-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 2);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end DualPortBootBRAM;

architecture arch of DualPortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"0b",
             2 => x"04",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"80",
            10 => x"0c",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"93",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"b4",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"b7",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"d2",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"cd",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"ff",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"8c",
           265 => x"0b",
           266 => x"04",
           267 => x"8c",
           268 => x"0b",
           269 => x"04",
           270 => x"8c",
           271 => x"0b",
           272 => x"04",
           273 => x"8c",
           274 => x"0b",
           275 => x"04",
           276 => x"8c",
           277 => x"0b",
           278 => x"04",
           279 => x"8d",
           280 => x"0b",
           281 => x"04",
           282 => x"8d",
           283 => x"0b",
           284 => x"04",
           285 => x"8d",
           286 => x"0b",
           287 => x"04",
           288 => x"8d",
           289 => x"0b",
           290 => x"04",
           291 => x"8e",
           292 => x"0b",
           293 => x"04",
           294 => x"8e",
           295 => x"0b",
           296 => x"04",
           297 => x"8e",
           298 => x"0b",
           299 => x"04",
           300 => x"8f",
           301 => x"0b",
           302 => x"04",
           303 => x"8f",
           304 => x"0b",
           305 => x"04",
           306 => x"8f",
           307 => x"0b",
           308 => x"04",
           309 => x"8f",
           310 => x"0b",
           311 => x"04",
           312 => x"90",
           313 => x"0b",
           314 => x"04",
           315 => x"90",
           316 => x"0b",
           317 => x"04",
           318 => x"90",
           319 => x"0b",
           320 => x"04",
           321 => x"90",
           322 => x"0b",
           323 => x"04",
           324 => x"91",
           325 => x"0b",
           326 => x"04",
           327 => x"91",
           328 => x"0b",
           329 => x"04",
           330 => x"91",
           331 => x"0b",
           332 => x"04",
           333 => x"91",
           334 => x"0b",
           335 => x"04",
           336 => x"92",
           337 => x"0b",
           338 => x"04",
           339 => x"92",
           340 => x"0b",
           341 => x"04",
           342 => x"92",
           343 => x"0b",
           344 => x"04",
           345 => x"93",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"81",
           385 => x"a4",
           386 => x"8b",
           387 => x"a4",
           388 => x"80",
           389 => x"e0",
           390 => x"e6",
           391 => x"a4",
           392 => x"80",
           393 => x"e0",
           394 => x"97",
           395 => x"a4",
           396 => x"80",
           397 => x"e0",
           398 => x"e1",
           399 => x"a4",
           400 => x"80",
           401 => x"e0",
           402 => x"e1",
           403 => x"a4",
           404 => x"80",
           405 => x"e0",
           406 => x"f6",
           407 => x"a4",
           408 => x"80",
           409 => x"e0",
           410 => x"da",
           411 => x"e0",
           412 => x"c0",
           413 => x"82",
           414 => x"80",
           415 => x"82",
           416 => x"80",
           417 => x"04",
           418 => x"0c",
           419 => x"82",
           420 => x"80",
           421 => x"04",
           422 => x"0c",
           423 => x"82",
           424 => x"80",
           425 => x"04",
           426 => x"0c",
           427 => x"82",
           428 => x"80",
           429 => x"04",
           430 => x"0c",
           431 => x"2d",
           432 => x"08",
           433 => x"90",
           434 => x"a4",
           435 => x"f6",
           436 => x"a4",
           437 => x"80",
           438 => x"e0",
           439 => x"80",
           440 => x"e0",
           441 => x"c0",
           442 => x"82",
           443 => x"80",
           444 => x"82",
           445 => x"80",
           446 => x"04",
           447 => x"0c",
           448 => x"2d",
           449 => x"08",
           450 => x"90",
           451 => x"a4",
           452 => x"a7",
           453 => x"a4",
           454 => x"80",
           455 => x"e0",
           456 => x"83",
           457 => x"e0",
           458 => x"c0",
           459 => x"82",
           460 => x"81",
           461 => x"82",
           462 => x"80",
           463 => x"04",
           464 => x"0c",
           465 => x"2d",
           466 => x"08",
           467 => x"90",
           468 => x"a4",
           469 => x"e5",
           470 => x"a4",
           471 => x"80",
           472 => x"e0",
           473 => x"91",
           474 => x"e0",
           475 => x"c0",
           476 => x"82",
           477 => x"82",
           478 => x"82",
           479 => x"80",
           480 => x"04",
           481 => x"0c",
           482 => x"2d",
           483 => x"08",
           484 => x"90",
           485 => x"a4",
           486 => x"a8",
           487 => x"a4",
           488 => x"80",
           489 => x"e0",
           490 => x"8d",
           491 => x"e0",
           492 => x"c0",
           493 => x"82",
           494 => x"82",
           495 => x"82",
           496 => x"80",
           497 => x"04",
           498 => x"0c",
           499 => x"2d",
           500 => x"08",
           501 => x"90",
           502 => x"a4",
           503 => x"97",
           504 => x"a4",
           505 => x"80",
           506 => x"e0",
           507 => x"8e",
           508 => x"e0",
           509 => x"c0",
           510 => x"82",
           511 => x"82",
           512 => x"82",
           513 => x"80",
           514 => x"04",
           515 => x"0c",
           516 => x"2d",
           517 => x"08",
           518 => x"90",
           519 => x"a4",
           520 => x"87",
           521 => x"a4",
           522 => x"80",
           523 => x"e0",
           524 => x"83",
           525 => x"e0",
           526 => x"c0",
           527 => x"82",
           528 => x"82",
           529 => x"82",
           530 => x"80",
           531 => x"04",
           532 => x"0c",
           533 => x"2d",
           534 => x"08",
           535 => x"90",
           536 => x"a4",
           537 => x"8e",
           538 => x"a4",
           539 => x"80",
           540 => x"e0",
           541 => x"9f",
           542 => x"e0",
           543 => x"c0",
           544 => x"82",
           545 => x"82",
           546 => x"82",
           547 => x"80",
           548 => x"04",
           549 => x"0c",
           550 => x"2d",
           551 => x"08",
           552 => x"90",
           553 => x"a4",
           554 => x"8c",
           555 => x"a4",
           556 => x"80",
           557 => x"e0",
           558 => x"b4",
           559 => x"e0",
           560 => x"c0",
           561 => x"82",
           562 => x"82",
           563 => x"82",
           564 => x"80",
           565 => x"04",
           566 => x"0c",
           567 => x"2d",
           568 => x"08",
           569 => x"90",
           570 => x"a4",
           571 => x"f5",
           572 => x"a4",
           573 => x"80",
           574 => x"e0",
           575 => x"b8",
           576 => x"e0",
           577 => x"c0",
           578 => x"82",
           579 => x"80",
           580 => x"82",
           581 => x"80",
           582 => x"04",
           583 => x"0c",
           584 => x"2d",
           585 => x"08",
           586 => x"90",
           587 => x"a4",
           588 => x"80",
           589 => x"a4",
           590 => x"80",
           591 => x"e0",
           592 => x"e0",
           593 => x"e0",
           594 => x"c0",
           595 => x"82",
           596 => x"81",
           597 => x"82",
           598 => x"80",
           599 => x"04",
           600 => x"0c",
           601 => x"2d",
           602 => x"08",
           603 => x"90",
           604 => x"a4",
           605 => x"bf",
           606 => x"a4",
           607 => x"80",
           608 => x"e0",
           609 => x"ac",
           610 => x"e0",
           611 => x"c0",
           612 => x"3c",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"10",
           621 => x"00",
           622 => x"ff",
           623 => x"06",
           624 => x"83",
           625 => x"10",
           626 => x"fc",
           627 => x"51",
           628 => x"80",
           629 => x"ff",
           630 => x"06",
           631 => x"52",
           632 => x"0a",
           633 => x"38",
           634 => x"51",
           635 => x"98",
           636 => x"84",
           637 => x"80",
           638 => x"05",
           639 => x"0b",
           640 => x"04",
           641 => x"80",
           642 => x"00",
           643 => x"08",
           644 => x"a4",
           645 => x"0d",
           646 => x"08",
           647 => x"82",
           648 => x"fc",
           649 => x"e0",
           650 => x"05",
           651 => x"e0",
           652 => x"05",
           653 => x"fb",
           654 => x"54",
           655 => x"82",
           656 => x"70",
           657 => x"08",
           658 => x"82",
           659 => x"f8",
           660 => x"82",
           661 => x"51",
           662 => x"0d",
           663 => x"0c",
           664 => x"a4",
           665 => x"e0",
           666 => x"3d",
           667 => x"a4",
           668 => x"08",
           669 => x"70",
           670 => x"81",
           671 => x"51",
           672 => x"38",
           673 => x"e0",
           674 => x"05",
           675 => x"38",
           676 => x"0b",
           677 => x"08",
           678 => x"81",
           679 => x"e0",
           680 => x"05",
           681 => x"82",
           682 => x"8c",
           683 => x"0b",
           684 => x"08",
           685 => x"82",
           686 => x"88",
           687 => x"e0",
           688 => x"05",
           689 => x"a4",
           690 => x"08",
           691 => x"f6",
           692 => x"82",
           693 => x"8c",
           694 => x"80",
           695 => x"e0",
           696 => x"05",
           697 => x"90",
           698 => x"98",
           699 => x"e0",
           700 => x"05",
           701 => x"e0",
           702 => x"05",
           703 => x"09",
           704 => x"38",
           705 => x"e0",
           706 => x"05",
           707 => x"39",
           708 => x"08",
           709 => x"82",
           710 => x"f8",
           711 => x"53",
           712 => x"82",
           713 => x"8c",
           714 => x"05",
           715 => x"08",
           716 => x"82",
           717 => x"fc",
           718 => x"05",
           719 => x"08",
           720 => x"ff",
           721 => x"e0",
           722 => x"05",
           723 => x"72",
           724 => x"a4",
           725 => x"08",
           726 => x"a4",
           727 => x"0c",
           728 => x"a4",
           729 => x"08",
           730 => x"0c",
           731 => x"82",
           732 => x"04",
           733 => x"08",
           734 => x"a4",
           735 => x"0d",
           736 => x"e0",
           737 => x"05",
           738 => x"a4",
           739 => x"08",
           740 => x"08",
           741 => x"fe",
           742 => x"e0",
           743 => x"05",
           744 => x"a4",
           745 => x"70",
           746 => x"08",
           747 => x"82",
           748 => x"fc",
           749 => x"82",
           750 => x"8c",
           751 => x"82",
           752 => x"e0",
           753 => x"51",
           754 => x"3f",
           755 => x"08",
           756 => x"a4",
           757 => x"0c",
           758 => x"08",
           759 => x"82",
           760 => x"88",
           761 => x"51",
           762 => x"34",
           763 => x"08",
           764 => x"70",
           765 => x"0c",
           766 => x"0d",
           767 => x"0c",
           768 => x"a4",
           769 => x"e0",
           770 => x"3d",
           771 => x"a4",
           772 => x"70",
           773 => x"08",
           774 => x"82",
           775 => x"fc",
           776 => x"82",
           777 => x"8c",
           778 => x"82",
           779 => x"88",
           780 => x"54",
           781 => x"e0",
           782 => x"82",
           783 => x"f8",
           784 => x"e0",
           785 => x"05",
           786 => x"e0",
           787 => x"54",
           788 => x"82",
           789 => x"04",
           790 => x"08",
           791 => x"a4",
           792 => x"0d",
           793 => x"e0",
           794 => x"05",
           795 => x"a4",
           796 => x"08",
           797 => x"8c",
           798 => x"e0",
           799 => x"05",
           800 => x"33",
           801 => x"70",
           802 => x"81",
           803 => x"51",
           804 => x"80",
           805 => x"ff",
           806 => x"a4",
           807 => x"0c",
           808 => x"82",
           809 => x"8c",
           810 => x"72",
           811 => x"82",
           812 => x"f8",
           813 => x"81",
           814 => x"72",
           815 => x"fa",
           816 => x"a4",
           817 => x"08",
           818 => x"e0",
           819 => x"05",
           820 => x"a4",
           821 => x"22",
           822 => x"51",
           823 => x"2e",
           824 => x"82",
           825 => x"f8",
           826 => x"af",
           827 => x"fc",
           828 => x"a4",
           829 => x"33",
           830 => x"26",
           831 => x"82",
           832 => x"f8",
           833 => x"72",
           834 => x"81",
           835 => x"38",
           836 => x"08",
           837 => x"70",
           838 => x"98",
           839 => x"53",
           840 => x"82",
           841 => x"e4",
           842 => x"83",
           843 => x"32",
           844 => x"51",
           845 => x"72",
           846 => x"38",
           847 => x"08",
           848 => x"70",
           849 => x"51",
           850 => x"e0",
           851 => x"05",
           852 => x"39",
           853 => x"08",
           854 => x"70",
           855 => x"98",
           856 => x"83",
           857 => x"73",
           858 => x"51",
           859 => x"53",
           860 => x"a4",
           861 => x"34",
           862 => x"08",
           863 => x"54",
           864 => x"08",
           865 => x"70",
           866 => x"51",
           867 => x"82",
           868 => x"e8",
           869 => x"e0",
           870 => x"05",
           871 => x"2b",
           872 => x"51",
           873 => x"80",
           874 => x"80",
           875 => x"e0",
           876 => x"05",
           877 => x"a4",
           878 => x"22",
           879 => x"70",
           880 => x"51",
           881 => x"db",
           882 => x"a4",
           883 => x"33",
           884 => x"70",
           885 => x"90",
           886 => x"2c",
           887 => x"51",
           888 => x"e0",
           889 => x"05",
           890 => x"39",
           891 => x"08",
           892 => x"70",
           893 => x"81",
           894 => x"53",
           895 => x"9d",
           896 => x"a4",
           897 => x"33",
           898 => x"70",
           899 => x"51",
           900 => x"38",
           901 => x"e0",
           902 => x"05",
           903 => x"a4",
           904 => x"33",
           905 => x"e0",
           906 => x"05",
           907 => x"e0",
           908 => x"05",
           909 => x"26",
           910 => x"82",
           911 => x"c4",
           912 => x"82",
           913 => x"dc",
           914 => x"51",
           915 => x"72",
           916 => x"a4",
           917 => x"22",
           918 => x"51",
           919 => x"e0",
           920 => x"05",
           921 => x"a4",
           922 => x"22",
           923 => x"51",
           924 => x"e0",
           925 => x"05",
           926 => x"39",
           927 => x"08",
           928 => x"70",
           929 => x"51",
           930 => x"e0",
           931 => x"05",
           932 => x"39",
           933 => x"08",
           934 => x"70",
           935 => x"51",
           936 => x"e0",
           937 => x"05",
           938 => x"39",
           939 => x"08",
           940 => x"70",
           941 => x"53",
           942 => x"a4",
           943 => x"23",
           944 => x"e0",
           945 => x"05",
           946 => x"39",
           947 => x"08",
           948 => x"70",
           949 => x"53",
           950 => x"a4",
           951 => x"23",
           952 => x"bf",
           953 => x"a4",
           954 => x"34",
           955 => x"08",
           956 => x"ff",
           957 => x"72",
           958 => x"08",
           959 => x"80",
           960 => x"e0",
           961 => x"05",
           962 => x"39",
           963 => x"08",
           964 => x"82",
           965 => x"90",
           966 => x"05",
           967 => x"08",
           968 => x"70",
           969 => x"72",
           970 => x"08",
           971 => x"82",
           972 => x"ec",
           973 => x"11",
           974 => x"82",
           975 => x"ec",
           976 => x"ef",
           977 => x"a4",
           978 => x"08",
           979 => x"08",
           980 => x"84",
           981 => x"a4",
           982 => x"0c",
           983 => x"e0",
           984 => x"05",
           985 => x"a4",
           986 => x"22",
           987 => x"70",
           988 => x"51",
           989 => x"80",
           990 => x"82",
           991 => x"e8",
           992 => x"98",
           993 => x"98",
           994 => x"e0",
           995 => x"05",
           996 => x"a4",
           997 => x"e0",
           998 => x"72",
           999 => x"08",
          1000 => x"99",
          1001 => x"a4",
          1002 => x"08",
          1003 => x"3f",
          1004 => x"08",
          1005 => x"e0",
          1006 => x"05",
          1007 => x"a4",
          1008 => x"22",
          1009 => x"a4",
          1010 => x"22",
          1011 => x"54",
          1012 => x"e0",
          1013 => x"05",
          1014 => x"39",
          1015 => x"08",
          1016 => x"82",
          1017 => x"90",
          1018 => x"05",
          1019 => x"08",
          1020 => x"70",
          1021 => x"a4",
          1022 => x"0c",
          1023 => x"08",
          1024 => x"70",
          1025 => x"81",
          1026 => x"51",
          1027 => x"2e",
          1028 => x"e0",
          1029 => x"05",
          1030 => x"2b",
          1031 => x"2c",
          1032 => x"a4",
          1033 => x"08",
          1034 => x"ec",
          1035 => x"98",
          1036 => x"82",
          1037 => x"f4",
          1038 => x"39",
          1039 => x"08",
          1040 => x"51",
          1041 => x"82",
          1042 => x"53",
          1043 => x"a4",
          1044 => x"23",
          1045 => x"08",
          1046 => x"53",
          1047 => x"08",
          1048 => x"73",
          1049 => x"54",
          1050 => x"a4",
          1051 => x"23",
          1052 => x"82",
          1053 => x"e4",
          1054 => x"82",
          1055 => x"06",
          1056 => x"72",
          1057 => x"38",
          1058 => x"08",
          1059 => x"82",
          1060 => x"90",
          1061 => x"05",
          1062 => x"08",
          1063 => x"70",
          1064 => x"a4",
          1065 => x"0c",
          1066 => x"82",
          1067 => x"90",
          1068 => x"e0",
          1069 => x"05",
          1070 => x"82",
          1071 => x"90",
          1072 => x"08",
          1073 => x"08",
          1074 => x"53",
          1075 => x"08",
          1076 => x"82",
          1077 => x"fc",
          1078 => x"e0",
          1079 => x"05",
          1080 => x"a4",
          1081 => x"a4",
          1082 => x"22",
          1083 => x"51",
          1084 => x"e0",
          1085 => x"05",
          1086 => x"a4",
          1087 => x"08",
          1088 => x"a4",
          1089 => x"0c",
          1090 => x"08",
          1091 => x"70",
          1092 => x"51",
          1093 => x"e0",
          1094 => x"05",
          1095 => x"39",
          1096 => x"e0",
          1097 => x"05",
          1098 => x"82",
          1099 => x"e4",
          1100 => x"80",
          1101 => x"53",
          1102 => x"a4",
          1103 => x"23",
          1104 => x"82",
          1105 => x"f8",
          1106 => x"0b",
          1107 => x"08",
          1108 => x"82",
          1109 => x"e4",
          1110 => x"82",
          1111 => x"06",
          1112 => x"72",
          1113 => x"38",
          1114 => x"08",
          1115 => x"82",
          1116 => x"90",
          1117 => x"05",
          1118 => x"08",
          1119 => x"70",
          1120 => x"a4",
          1121 => x"0c",
          1122 => x"82",
          1123 => x"90",
          1124 => x"e0",
          1125 => x"05",
          1126 => x"82",
          1127 => x"90",
          1128 => x"08",
          1129 => x"08",
          1130 => x"53",
          1131 => x"08",
          1132 => x"82",
          1133 => x"fc",
          1134 => x"e0",
          1135 => x"05",
          1136 => x"06",
          1137 => x"82",
          1138 => x"e4",
          1139 => x"e0",
          1140 => x"e0",
          1141 => x"05",
          1142 => x"a4",
          1143 => x"08",
          1144 => x"08",
          1145 => x"82",
          1146 => x"fc",
          1147 => x"55",
          1148 => x"54",
          1149 => x"3f",
          1150 => x"08",
          1151 => x"34",
          1152 => x"08",
          1153 => x"82",
          1154 => x"d4",
          1155 => x"e0",
          1156 => x"05",
          1157 => x"51",
          1158 => x"27",
          1159 => x"e0",
          1160 => x"05",
          1161 => x"33",
          1162 => x"a4",
          1163 => x"33",
          1164 => x"11",
          1165 => x"72",
          1166 => x"08",
          1167 => x"97",
          1168 => x"a4",
          1169 => x"08",
          1170 => x"b0",
          1171 => x"72",
          1172 => x"08",
          1173 => x"82",
          1174 => x"d4",
          1175 => x"82",
          1176 => x"d0",
          1177 => x"34",
          1178 => x"08",
          1179 => x"81",
          1180 => x"a4",
          1181 => x"0c",
          1182 => x"08",
          1183 => x"70",
          1184 => x"a4",
          1185 => x"08",
          1186 => x"c7",
          1187 => x"98",
          1188 => x"e0",
          1189 => x"05",
          1190 => x"e0",
          1191 => x"05",
          1192 => x"84",
          1193 => x"39",
          1194 => x"08",
          1195 => x"82",
          1196 => x"55",
          1197 => x"70",
          1198 => x"53",
          1199 => x"a4",
          1200 => x"34",
          1201 => x"08",
          1202 => x"70",
          1203 => x"53",
          1204 => x"94",
          1205 => x"a4",
          1206 => x"22",
          1207 => x"53",
          1208 => x"a4",
          1209 => x"23",
          1210 => x"08",
          1211 => x"70",
          1212 => x"81",
          1213 => x"53",
          1214 => x"80",
          1215 => x"e0",
          1216 => x"05",
          1217 => x"2b",
          1218 => x"08",
          1219 => x"82",
          1220 => x"cc",
          1221 => x"2c",
          1222 => x"08",
          1223 => x"82",
          1224 => x"f4",
          1225 => x"53",
          1226 => x"09",
          1227 => x"38",
          1228 => x"08",
          1229 => x"fe",
          1230 => x"82",
          1231 => x"c8",
          1232 => x"39",
          1233 => x"08",
          1234 => x"ff",
          1235 => x"82",
          1236 => x"c8",
          1237 => x"e0",
          1238 => x"05",
          1239 => x"a4",
          1240 => x"23",
          1241 => x"08",
          1242 => x"70",
          1243 => x"81",
          1244 => x"53",
          1245 => x"80",
          1246 => x"e0",
          1247 => x"05",
          1248 => x"2b",
          1249 => x"82",
          1250 => x"fc",
          1251 => x"51",
          1252 => x"74",
          1253 => x"82",
          1254 => x"e4",
          1255 => x"f7",
          1256 => x"72",
          1257 => x"08",
          1258 => x"9d",
          1259 => x"a4",
          1260 => x"33",
          1261 => x"a4",
          1262 => x"33",
          1263 => x"54",
          1264 => x"e0",
          1265 => x"05",
          1266 => x"a4",
          1267 => x"22",
          1268 => x"70",
          1269 => x"51",
          1270 => x"2e",
          1271 => x"e0",
          1272 => x"05",
          1273 => x"2b",
          1274 => x"70",
          1275 => x"88",
          1276 => x"51",
          1277 => x"54",
          1278 => x"08",
          1279 => x"70",
          1280 => x"53",
          1281 => x"a4",
          1282 => x"23",
          1283 => x"e0",
          1284 => x"05",
          1285 => x"2b",
          1286 => x"70",
          1287 => x"88",
          1288 => x"51",
          1289 => x"54",
          1290 => x"08",
          1291 => x"70",
          1292 => x"53",
          1293 => x"a4",
          1294 => x"23",
          1295 => x"08",
          1296 => x"70",
          1297 => x"51",
          1298 => x"38",
          1299 => x"08",
          1300 => x"ff",
          1301 => x"72",
          1302 => x"08",
          1303 => x"73",
          1304 => x"90",
          1305 => x"80",
          1306 => x"38",
          1307 => x"08",
          1308 => x"52",
          1309 => x"ee",
          1310 => x"82",
          1311 => x"e4",
          1312 => x"81",
          1313 => x"06",
          1314 => x"72",
          1315 => x"38",
          1316 => x"08",
          1317 => x"52",
          1318 => x"ca",
          1319 => x"39",
          1320 => x"08",
          1321 => x"70",
          1322 => x"81",
          1323 => x"53",
          1324 => x"90",
          1325 => x"a4",
          1326 => x"08",
          1327 => x"8a",
          1328 => x"39",
          1329 => x"08",
          1330 => x"70",
          1331 => x"81",
          1332 => x"53",
          1333 => x"8e",
          1334 => x"a4",
          1335 => x"08",
          1336 => x"8a",
          1337 => x"e0",
          1338 => x"05",
          1339 => x"2a",
          1340 => x"51",
          1341 => x"80",
          1342 => x"82",
          1343 => x"88",
          1344 => x"b0",
          1345 => x"3f",
          1346 => x"08",
          1347 => x"53",
          1348 => x"09",
          1349 => x"38",
          1350 => x"08",
          1351 => x"52",
          1352 => x"08",
          1353 => x"51",
          1354 => x"82",
          1355 => x"e4",
          1356 => x"88",
          1357 => x"06",
          1358 => x"72",
          1359 => x"38",
          1360 => x"08",
          1361 => x"ff",
          1362 => x"72",
          1363 => x"08",
          1364 => x"73",
          1365 => x"90",
          1366 => x"80",
          1367 => x"38",
          1368 => x"08",
          1369 => x"52",
          1370 => x"fa",
          1371 => x"82",
          1372 => x"e4",
          1373 => x"83",
          1374 => x"06",
          1375 => x"72",
          1376 => x"38",
          1377 => x"08",
          1378 => x"ff",
          1379 => x"72",
          1380 => x"08",
          1381 => x"73",
          1382 => x"98",
          1383 => x"80",
          1384 => x"38",
          1385 => x"08",
          1386 => x"52",
          1387 => x"b6",
          1388 => x"82",
          1389 => x"e4",
          1390 => x"87",
          1391 => x"06",
          1392 => x"72",
          1393 => x"e0",
          1394 => x"05",
          1395 => x"54",
          1396 => x"e0",
          1397 => x"05",
          1398 => x"2b",
          1399 => x"51",
          1400 => x"25",
          1401 => x"e0",
          1402 => x"05",
          1403 => x"51",
          1404 => x"d2",
          1405 => x"a4",
          1406 => x"33",
          1407 => x"e3",
          1408 => x"06",
          1409 => x"e0",
          1410 => x"05",
          1411 => x"e0",
          1412 => x"05",
          1413 => x"ce",
          1414 => x"39",
          1415 => x"08",
          1416 => x"53",
          1417 => x"2e",
          1418 => x"80",
          1419 => x"e0",
          1420 => x"05",
          1421 => x"51",
          1422 => x"e0",
          1423 => x"05",
          1424 => x"ff",
          1425 => x"72",
          1426 => x"2e",
          1427 => x"82",
          1428 => x"88",
          1429 => x"82",
          1430 => x"fc",
          1431 => x"33",
          1432 => x"a4",
          1433 => x"08",
          1434 => x"e0",
          1435 => x"05",
          1436 => x"f2",
          1437 => x"39",
          1438 => x"08",
          1439 => x"53",
          1440 => x"2e",
          1441 => x"80",
          1442 => x"e0",
          1443 => x"05",
          1444 => x"51",
          1445 => x"e0",
          1446 => x"05",
          1447 => x"ff",
          1448 => x"72",
          1449 => x"2e",
          1450 => x"82",
          1451 => x"88",
          1452 => x"82",
          1453 => x"fc",
          1454 => x"33",
          1455 => x"a6",
          1456 => x"a4",
          1457 => x"08",
          1458 => x"e0",
          1459 => x"05",
          1460 => x"39",
          1461 => x"08",
          1462 => x"82",
          1463 => x"a9",
          1464 => x"a4",
          1465 => x"08",
          1466 => x"a4",
          1467 => x"08",
          1468 => x"e0",
          1469 => x"05",
          1470 => x"a4",
          1471 => x"08",
          1472 => x"53",
          1473 => x"cc",
          1474 => x"a4",
          1475 => x"22",
          1476 => x"70",
          1477 => x"51",
          1478 => x"2e",
          1479 => x"82",
          1480 => x"ec",
          1481 => x"11",
          1482 => x"82",
          1483 => x"ec",
          1484 => x"90",
          1485 => x"2c",
          1486 => x"73",
          1487 => x"82",
          1488 => x"88",
          1489 => x"a0",
          1490 => x"3f",
          1491 => x"e0",
          1492 => x"05",
          1493 => x"e0",
          1494 => x"05",
          1495 => x"86",
          1496 => x"82",
          1497 => x"e4",
          1498 => x"b7",
          1499 => x"a4",
          1500 => x"33",
          1501 => x"2e",
          1502 => x"a8",
          1503 => x"82",
          1504 => x"e4",
          1505 => x"0b",
          1506 => x"08",
          1507 => x"80",
          1508 => x"a4",
          1509 => x"34",
          1510 => x"e0",
          1511 => x"05",
          1512 => x"39",
          1513 => x"08",
          1514 => x"52",
          1515 => x"08",
          1516 => x"51",
          1517 => x"e9",
          1518 => x"e0",
          1519 => x"05",
          1520 => x"08",
          1521 => x"a4",
          1522 => x"0c",
          1523 => x"e0",
          1524 => x"05",
          1525 => x"98",
          1526 => x"0d",
          1527 => x"0c",
          1528 => x"a4",
          1529 => x"e0",
          1530 => x"3d",
          1531 => x"f8",
          1532 => x"e0",
          1533 => x"05",
          1534 => x"e0",
          1535 => x"05",
          1536 => x"dd",
          1537 => x"98",
          1538 => x"e0",
          1539 => x"85",
          1540 => x"e0",
          1541 => x"82",
          1542 => x"02",
          1543 => x"0c",
          1544 => x"80",
          1545 => x"a4",
          1546 => x"0c",
          1547 => x"08",
          1548 => x"70",
          1549 => x"81",
          1550 => x"06",
          1551 => x"51",
          1552 => x"2e",
          1553 => x"0b",
          1554 => x"08",
          1555 => x"81",
          1556 => x"e0",
          1557 => x"05",
          1558 => x"33",
          1559 => x"08",
          1560 => x"81",
          1561 => x"a4",
          1562 => x"0c",
          1563 => x"e0",
          1564 => x"05",
          1565 => x"ff",
          1566 => x"80",
          1567 => x"82",
          1568 => x"82",
          1569 => x"53",
          1570 => x"08",
          1571 => x"52",
          1572 => x"51",
          1573 => x"82",
          1574 => x"53",
          1575 => x"ff",
          1576 => x"0b",
          1577 => x"08",
          1578 => x"ff",
          1579 => x"fb",
          1580 => x"fb",
          1581 => x"53",
          1582 => x"13",
          1583 => x"2d",
          1584 => x"08",
          1585 => x"2e",
          1586 => x"0b",
          1587 => x"08",
          1588 => x"82",
          1589 => x"f8",
          1590 => x"82",
          1591 => x"f4",
          1592 => x"82",
          1593 => x"f4",
          1594 => x"e0",
          1595 => x"3d",
          1596 => x"a4",
          1597 => x"e0",
          1598 => x"82",
          1599 => x"fb",
          1600 => x"0b",
          1601 => x"08",
          1602 => x"82",
          1603 => x"8c",
          1604 => x"11",
          1605 => x"2a",
          1606 => x"70",
          1607 => x"51",
          1608 => x"72",
          1609 => x"38",
          1610 => x"e0",
          1611 => x"05",
          1612 => x"39",
          1613 => x"08",
          1614 => x"53",
          1615 => x"e0",
          1616 => x"05",
          1617 => x"82",
          1618 => x"88",
          1619 => x"72",
          1620 => x"08",
          1621 => x"72",
          1622 => x"53",
          1623 => x"b6",
          1624 => x"a4",
          1625 => x"08",
          1626 => x"08",
          1627 => x"53",
          1628 => x"08",
          1629 => x"52",
          1630 => x"51",
          1631 => x"82",
          1632 => x"53",
          1633 => x"ff",
          1634 => x"0b",
          1635 => x"08",
          1636 => x"ff",
          1637 => x"e0",
          1638 => x"05",
          1639 => x"e0",
          1640 => x"05",
          1641 => x"e0",
          1642 => x"05",
          1643 => x"98",
          1644 => x"0d",
          1645 => x"0c",
          1646 => x"a4",
          1647 => x"e0",
          1648 => x"3d",
          1649 => x"fc",
          1650 => x"e0",
          1651 => x"05",
          1652 => x"3f",
          1653 => x"08",
          1654 => x"98",
          1655 => x"3d",
          1656 => x"a4",
          1657 => x"e0",
          1658 => x"82",
          1659 => x"fb",
          1660 => x"e0",
          1661 => x"05",
          1662 => x"33",
          1663 => x"70",
          1664 => x"81",
          1665 => x"51",
          1666 => x"80",
          1667 => x"ff",
          1668 => x"a4",
          1669 => x"0c",
          1670 => x"82",
          1671 => x"8c",
          1672 => x"11",
          1673 => x"2a",
          1674 => x"51",
          1675 => x"72",
          1676 => x"db",
          1677 => x"a4",
          1678 => x"08",
          1679 => x"08",
          1680 => x"54",
          1681 => x"08",
          1682 => x"25",
          1683 => x"e0",
          1684 => x"05",
          1685 => x"70",
          1686 => x"08",
          1687 => x"52",
          1688 => x"72",
          1689 => x"08",
          1690 => x"0c",
          1691 => x"08",
          1692 => x"8c",
          1693 => x"05",
          1694 => x"82",
          1695 => x"88",
          1696 => x"82",
          1697 => x"fc",
          1698 => x"53",
          1699 => x"82",
          1700 => x"8c",
          1701 => x"e0",
          1702 => x"05",
          1703 => x"e0",
          1704 => x"05",
          1705 => x"ff",
          1706 => x"12",
          1707 => x"54",
          1708 => x"e0",
          1709 => x"72",
          1710 => x"e0",
          1711 => x"05",
          1712 => x"08",
          1713 => x"12",
          1714 => x"a4",
          1715 => x"08",
          1716 => x"a4",
          1717 => x"0c",
          1718 => x"39",
          1719 => x"e0",
          1720 => x"05",
          1721 => x"a4",
          1722 => x"08",
          1723 => x"0c",
          1724 => x"82",
          1725 => x"04",
          1726 => x"08",
          1727 => x"a4",
          1728 => x"0d",
          1729 => x"08",
          1730 => x"85",
          1731 => x"81",
          1732 => x"06",
          1733 => x"52",
          1734 => x"8d",
          1735 => x"82",
          1736 => x"f8",
          1737 => x"94",
          1738 => x"a4",
          1739 => x"08",
          1740 => x"70",
          1741 => x"81",
          1742 => x"51",
          1743 => x"2e",
          1744 => x"82",
          1745 => x"88",
          1746 => x"e0",
          1747 => x"05",
          1748 => x"85",
          1749 => x"ff",
          1750 => x"52",
          1751 => x"34",
          1752 => x"08",
          1753 => x"8c",
          1754 => x"05",
          1755 => x"82",
          1756 => x"88",
          1757 => x"11",
          1758 => x"e0",
          1759 => x"05",
          1760 => x"52",
          1761 => x"82",
          1762 => x"88",
          1763 => x"11",
          1764 => x"2a",
          1765 => x"51",
          1766 => x"71",
          1767 => x"d7",
          1768 => x"a4",
          1769 => x"08",
          1770 => x"33",
          1771 => x"08",
          1772 => x"51",
          1773 => x"a4",
          1774 => x"08",
          1775 => x"e0",
          1776 => x"05",
          1777 => x"a4",
          1778 => x"08",
          1779 => x"12",
          1780 => x"07",
          1781 => x"85",
          1782 => x"0b",
          1783 => x"08",
          1784 => x"81",
          1785 => x"e0",
          1786 => x"05",
          1787 => x"81",
          1788 => x"52",
          1789 => x"82",
          1790 => x"88",
          1791 => x"e0",
          1792 => x"05",
          1793 => x"11",
          1794 => x"71",
          1795 => x"98",
          1796 => x"e0",
          1797 => x"05",
          1798 => x"e0",
          1799 => x"05",
          1800 => x"80",
          1801 => x"e0",
          1802 => x"05",
          1803 => x"a4",
          1804 => x"0c",
          1805 => x"08",
          1806 => x"85",
          1807 => x"e0",
          1808 => x"05",
          1809 => x"e0",
          1810 => x"05",
          1811 => x"09",
          1812 => x"38",
          1813 => x"08",
          1814 => x"90",
          1815 => x"82",
          1816 => x"ec",
          1817 => x"39",
          1818 => x"08",
          1819 => x"a0",
          1820 => x"82",
          1821 => x"ec",
          1822 => x"e0",
          1823 => x"05",
          1824 => x"e0",
          1825 => x"05",
          1826 => x"34",
          1827 => x"e0",
          1828 => x"05",
          1829 => x"82",
          1830 => x"88",
          1831 => x"11",
          1832 => x"8c",
          1833 => x"e0",
          1834 => x"05",
          1835 => x"ff",
          1836 => x"e0",
          1837 => x"05",
          1838 => x"52",
          1839 => x"08",
          1840 => x"82",
          1841 => x"89",
          1842 => x"e0",
          1843 => x"82",
          1844 => x"02",
          1845 => x"0c",
          1846 => x"82",
          1847 => x"88",
          1848 => x"e0",
          1849 => x"05",
          1850 => x"a4",
          1851 => x"08",
          1852 => x"08",
          1853 => x"82",
          1854 => x"90",
          1855 => x"2e",
          1856 => x"82",
          1857 => x"f8",
          1858 => x"e0",
          1859 => x"05",
          1860 => x"ac",
          1861 => x"a4",
          1862 => x"08",
          1863 => x"08",
          1864 => x"05",
          1865 => x"a4",
          1866 => x"08",
          1867 => x"90",
          1868 => x"a4",
          1869 => x"08",
          1870 => x"08",
          1871 => x"05",
          1872 => x"08",
          1873 => x"82",
          1874 => x"f8",
          1875 => x"e0",
          1876 => x"05",
          1877 => x"e0",
          1878 => x"05",
          1879 => x"a4",
          1880 => x"08",
          1881 => x"e0",
          1882 => x"05",
          1883 => x"a4",
          1884 => x"08",
          1885 => x"e0",
          1886 => x"05",
          1887 => x"a4",
          1888 => x"08",
          1889 => x"9c",
          1890 => x"a4",
          1891 => x"08",
          1892 => x"e0",
          1893 => x"05",
          1894 => x"a4",
          1895 => x"08",
          1896 => x"e0",
          1897 => x"05",
          1898 => x"a4",
          1899 => x"08",
          1900 => x"08",
          1901 => x"53",
          1902 => x"71",
          1903 => x"39",
          1904 => x"08",
          1905 => x"81",
          1906 => x"a4",
          1907 => x"0c",
          1908 => x"08",
          1909 => x"ff",
          1910 => x"a4",
          1911 => x"0c",
          1912 => x"08",
          1913 => x"80",
          1914 => x"82",
          1915 => x"f8",
          1916 => x"70",
          1917 => x"a4",
          1918 => x"08",
          1919 => x"e0",
          1920 => x"05",
          1921 => x"a4",
          1922 => x"08",
          1923 => x"71",
          1924 => x"a4",
          1925 => x"08",
          1926 => x"e0",
          1927 => x"05",
          1928 => x"39",
          1929 => x"08",
          1930 => x"70",
          1931 => x"0c",
          1932 => x"0d",
          1933 => x"0c",
          1934 => x"a4",
          1935 => x"e0",
          1936 => x"3d",
          1937 => x"a4",
          1938 => x"08",
          1939 => x"08",
          1940 => x"82",
          1941 => x"fc",
          1942 => x"71",
          1943 => x"a4",
          1944 => x"08",
          1945 => x"e0",
          1946 => x"05",
          1947 => x"ff",
          1948 => x"70",
          1949 => x"38",
          1950 => x"e0",
          1951 => x"05",
          1952 => x"82",
          1953 => x"fc",
          1954 => x"e0",
          1955 => x"05",
          1956 => x"a4",
          1957 => x"08",
          1958 => x"e0",
          1959 => x"84",
          1960 => x"e0",
          1961 => x"82",
          1962 => x"02",
          1963 => x"0c",
          1964 => x"82",
          1965 => x"88",
          1966 => x"e0",
          1967 => x"05",
          1968 => x"a4",
          1969 => x"08",
          1970 => x"82",
          1971 => x"8c",
          1972 => x"05",
          1973 => x"08",
          1974 => x"82",
          1975 => x"fc",
          1976 => x"51",
          1977 => x"82",
          1978 => x"fc",
          1979 => x"05",
          1980 => x"08",
          1981 => x"70",
          1982 => x"51",
          1983 => x"84",
          1984 => x"39",
          1985 => x"08",
          1986 => x"70",
          1987 => x"0c",
          1988 => x"0d",
          1989 => x"0c",
          1990 => x"a4",
          1991 => x"e0",
          1992 => x"3d",
          1993 => x"a4",
          1994 => x"08",
          1995 => x"08",
          1996 => x"82",
          1997 => x"8c",
          1998 => x"e0",
          1999 => x"05",
          2000 => x"a4",
          2001 => x"08",
          2002 => x"e5",
          2003 => x"a4",
          2004 => x"08",
          2005 => x"e0",
          2006 => x"05",
          2007 => x"a4",
          2008 => x"08",
          2009 => x"e0",
          2010 => x"05",
          2011 => x"a4",
          2012 => x"08",
          2013 => x"38",
          2014 => x"08",
          2015 => x"51",
          2016 => x"e0",
          2017 => x"05",
          2018 => x"82",
          2019 => x"f8",
          2020 => x"e0",
          2021 => x"05",
          2022 => x"71",
          2023 => x"e0",
          2024 => x"05",
          2025 => x"82",
          2026 => x"fc",
          2027 => x"ad",
          2028 => x"a4",
          2029 => x"08",
          2030 => x"98",
          2031 => x"3d",
          2032 => x"a4",
          2033 => x"e0",
          2034 => x"82",
          2035 => x"fd",
          2036 => x"e0",
          2037 => x"05",
          2038 => x"81",
          2039 => x"e0",
          2040 => x"05",
          2041 => x"33",
          2042 => x"08",
          2043 => x"81",
          2044 => x"a4",
          2045 => x"0c",
          2046 => x"08",
          2047 => x"70",
          2048 => x"ff",
          2049 => x"54",
          2050 => x"2e",
          2051 => x"ce",
          2052 => x"a4",
          2053 => x"08",
          2054 => x"82",
          2055 => x"88",
          2056 => x"05",
          2057 => x"08",
          2058 => x"70",
          2059 => x"51",
          2060 => x"38",
          2061 => x"e0",
          2062 => x"05",
          2063 => x"39",
          2064 => x"08",
          2065 => x"ff",
          2066 => x"a4",
          2067 => x"0c",
          2068 => x"08",
          2069 => x"80",
          2070 => x"ff",
          2071 => x"e0",
          2072 => x"05",
          2073 => x"80",
          2074 => x"e0",
          2075 => x"05",
          2076 => x"52",
          2077 => x"38",
          2078 => x"e0",
          2079 => x"05",
          2080 => x"39",
          2081 => x"08",
          2082 => x"ff",
          2083 => x"a4",
          2084 => x"0c",
          2085 => x"08",
          2086 => x"70",
          2087 => x"70",
          2088 => x"0b",
          2089 => x"08",
          2090 => x"ae",
          2091 => x"a4",
          2092 => x"08",
          2093 => x"e0",
          2094 => x"05",
          2095 => x"72",
          2096 => x"82",
          2097 => x"fc",
          2098 => x"55",
          2099 => x"8a",
          2100 => x"82",
          2101 => x"fc",
          2102 => x"e0",
          2103 => x"05",
          2104 => x"98",
          2105 => x"0d",
          2106 => x"0c",
          2107 => x"a4",
          2108 => x"e0",
          2109 => x"3d",
          2110 => x"a4",
          2111 => x"08",
          2112 => x"a4",
          2113 => x"08",
          2114 => x"3f",
          2115 => x"08",
          2116 => x"a4",
          2117 => x"0c",
          2118 => x"08",
          2119 => x"81",
          2120 => x"51",
          2121 => x"f7",
          2122 => x"98",
          2123 => x"e0",
          2124 => x"05",
          2125 => x"e0",
          2126 => x"05",
          2127 => x"80",
          2128 => x"a4",
          2129 => x"0c",
          2130 => x"e0",
          2131 => x"05",
          2132 => x"a4",
          2133 => x"08",
          2134 => x"74",
          2135 => x"a4",
          2136 => x"08",
          2137 => x"a4",
          2138 => x"08",
          2139 => x"a4",
          2140 => x"08",
          2141 => x"3f",
          2142 => x"08",
          2143 => x"a4",
          2144 => x"0c",
          2145 => x"a4",
          2146 => x"08",
          2147 => x"0c",
          2148 => x"82",
          2149 => x"04",
          2150 => x"08",
          2151 => x"a4",
          2152 => x"0d",
          2153 => x"08",
          2154 => x"82",
          2155 => x"f8",
          2156 => x"e0",
          2157 => x"05",
          2158 => x"80",
          2159 => x"a4",
          2160 => x"0c",
          2161 => x"82",
          2162 => x"f8",
          2163 => x"71",
          2164 => x"a4",
          2165 => x"08",
          2166 => x"e0",
          2167 => x"05",
          2168 => x"ff",
          2169 => x"70",
          2170 => x"38",
          2171 => x"08",
          2172 => x"ff",
          2173 => x"a4",
          2174 => x"0c",
          2175 => x"08",
          2176 => x"ff",
          2177 => x"ff",
          2178 => x"e0",
          2179 => x"05",
          2180 => x"82",
          2181 => x"f8",
          2182 => x"e0",
          2183 => x"05",
          2184 => x"a4",
          2185 => x"08",
          2186 => x"e0",
          2187 => x"05",
          2188 => x"e0",
          2189 => x"05",
          2190 => x"98",
          2191 => x"0d",
          2192 => x"0c",
          2193 => x"a4",
          2194 => x"e0",
          2195 => x"3d",
          2196 => x"a4",
          2197 => x"08",
          2198 => x"08",
          2199 => x"82",
          2200 => x"90",
          2201 => x"2e",
          2202 => x"82",
          2203 => x"90",
          2204 => x"05",
          2205 => x"08",
          2206 => x"82",
          2207 => x"90",
          2208 => x"05",
          2209 => x"08",
          2210 => x"82",
          2211 => x"90",
          2212 => x"2e",
          2213 => x"e0",
          2214 => x"05",
          2215 => x"82",
          2216 => x"fc",
          2217 => x"52",
          2218 => x"82",
          2219 => x"fc",
          2220 => x"05",
          2221 => x"08",
          2222 => x"ff",
          2223 => x"e0",
          2224 => x"05",
          2225 => x"e0",
          2226 => x"84",
          2227 => x"e0",
          2228 => x"82",
          2229 => x"02",
          2230 => x"0c",
          2231 => x"82",
          2232 => x"8c",
          2233 => x"82",
          2234 => x"88",
          2235 => x"93",
          2236 => x"98",
          2237 => x"e0",
          2238 => x"84",
          2239 => x"e0",
          2240 => x"82",
          2241 => x"02",
          2242 => x"0c",
          2243 => x"a0",
          2244 => x"a4",
          2245 => x"0c",
          2246 => x"08",
          2247 => x"80",
          2248 => x"82",
          2249 => x"8c",
          2250 => x"83",
          2251 => x"e0",
          2252 => x"82",
          2253 => x"e4",
          2254 => x"8f",
          2255 => x"a4",
          2256 => x"08",
          2257 => x"08",
          2258 => x"82",
          2259 => x"88",
          2260 => x"2e",
          2261 => x"e0",
          2262 => x"05",
          2263 => x"c9",
          2264 => x"98",
          2265 => x"a4",
          2266 => x"08",
          2267 => x"e0",
          2268 => x"05",
          2269 => x"39",
          2270 => x"08",
          2271 => x"82",
          2272 => x"fc",
          2273 => x"82",
          2274 => x"e0",
          2275 => x"e0",
          2276 => x"05",
          2277 => x"a4",
          2278 => x"0c",
          2279 => x"08",
          2280 => x"ff",
          2281 => x"82",
          2282 => x"f8",
          2283 => x"8d",
          2284 => x"82",
          2285 => x"e8",
          2286 => x"da",
          2287 => x"a4",
          2288 => x"08",
          2289 => x"71",
          2290 => x"08",
          2291 => x"2e",
          2292 => x"94",
          2293 => x"a4",
          2294 => x"08",
          2295 => x"a4",
          2296 => x"0c",
          2297 => x"39",
          2298 => x"08",
          2299 => x"81",
          2300 => x"a4",
          2301 => x"0c",
          2302 => x"08",
          2303 => x"82",
          2304 => x"f8",
          2305 => x"82",
          2306 => x"f4",
          2307 => x"e0",
          2308 => x"05",
          2309 => x"a4",
          2310 => x"08",
          2311 => x"a4",
          2312 => x"08",
          2313 => x"e0",
          2314 => x"05",
          2315 => x"0b",
          2316 => x"08",
          2317 => x"82",
          2318 => x"f8",
          2319 => x"2e",
          2320 => x"82",
          2321 => x"f4",
          2322 => x"82",
          2323 => x"fc",
          2324 => x"05",
          2325 => x"08",
          2326 => x"71",
          2327 => x"07",
          2328 => x"08",
          2329 => x"82",
          2330 => x"88",
          2331 => x"70",
          2332 => x"08",
          2333 => x"07",
          2334 => x"08",
          2335 => x"82",
          2336 => x"8c",
          2337 => x"e0",
          2338 => x"05",
          2339 => x"11",
          2340 => x"08",
          2341 => x"ff",
          2342 => x"2c",
          2343 => x"08",
          2344 => x"82",
          2345 => x"ec",
          2346 => x"06",
          2347 => x"08",
          2348 => x"82",
          2349 => x"8c",
          2350 => x"e0",
          2351 => x"05",
          2352 => x"e0",
          2353 => x"05",
          2354 => x"82",
          2355 => x"f4",
          2356 => x"e0",
          2357 => x"05",
          2358 => x"82",
          2359 => x"f8",
          2360 => x"52",
          2361 => x"51",
          2362 => x"cb",
          2363 => x"a4",
          2364 => x"08",
          2365 => x"e0",
          2366 => x"05",
          2367 => x"e0",
          2368 => x"05",
          2369 => x"a4",
          2370 => x"08",
          2371 => x"a4",
          2372 => x"0c",
          2373 => x"e0",
          2374 => x"05",
          2375 => x"98",
          2376 => x"0d",
          2377 => x"0c",
          2378 => x"a4",
          2379 => x"e0",
          2380 => x"3d",
          2381 => x"a4",
          2382 => x"08",
          2383 => x"08",
          2384 => x"82",
          2385 => x"fc",
          2386 => x"80",
          2387 => x"70",
          2388 => x"0b",
          2389 => x"08",
          2390 => x"8a",
          2391 => x"82",
          2392 => x"f0",
          2393 => x"e0",
          2394 => x"05",
          2395 => x"a4",
          2396 => x"0c",
          2397 => x"e0",
          2398 => x"05",
          2399 => x"e0",
          2400 => x"05",
          2401 => x"82",
          2402 => x"fc",
          2403 => x"e0",
          2404 => x"05",
          2405 => x"a4",
          2406 => x"0c",
          2407 => x"08",
          2408 => x"83",
          2409 => x"51",
          2410 => x"38",
          2411 => x"e0",
          2412 => x"05",
          2413 => x"80",
          2414 => x"a4",
          2415 => x"0c",
          2416 => x"08",
          2417 => x"82",
          2418 => x"f8",
          2419 => x"0b",
          2420 => x"08",
          2421 => x"31",
          2422 => x"08",
          2423 => x"71",
          2424 => x"a4",
          2425 => x"0c",
          2426 => x"08",
          2427 => x"82",
          2428 => x"f8",
          2429 => x"82",
          2430 => x"f4",
          2431 => x"e0",
          2432 => x"05",
          2433 => x"06",
          2434 => x"8c",
          2435 => x"82",
          2436 => x"e8",
          2437 => x"39",
          2438 => x"e0",
          2439 => x"05",
          2440 => x"a4",
          2441 => x"08",
          2442 => x"08",
          2443 => x"84",
          2444 => x"a4",
          2445 => x"08",
          2446 => x"a4",
          2447 => x"08",
          2448 => x"e0",
          2449 => x"05",
          2450 => x"a4",
          2451 => x"08",
          2452 => x"08",
          2453 => x"05",
          2454 => x"08",
          2455 => x"82",
          2456 => x"fc",
          2457 => x"06",
          2458 => x"8c",
          2459 => x"82",
          2460 => x"e4",
          2461 => x"39",
          2462 => x"e0",
          2463 => x"05",
          2464 => x"a4",
          2465 => x"08",
          2466 => x"08",
          2467 => x"82",
          2468 => x"a4",
          2469 => x"08",
          2470 => x"a4",
          2471 => x"08",
          2472 => x"e0",
          2473 => x"05",
          2474 => x"a4",
          2475 => x"08",
          2476 => x"08",
          2477 => x"05",
          2478 => x"08",
          2479 => x"82",
          2480 => x"a4",
          2481 => x"08",
          2482 => x"a4",
          2483 => x"08",
          2484 => x"81",
          2485 => x"06",
          2486 => x"75",
          2487 => x"a4",
          2488 => x"08",
          2489 => x"82",
          2490 => x"53",
          2491 => x"51",
          2492 => x"51",
          2493 => x"82",
          2494 => x"04",
          2495 => x"08",
          2496 => x"a4",
          2497 => x"0d",
          2498 => x"08",
          2499 => x"52",
          2500 => x"08",
          2501 => x"51",
          2502 => x"82",
          2503 => x"70",
          2504 => x"08",
          2505 => x"29",
          2506 => x"08",
          2507 => x"71",
          2508 => x"e0",
          2509 => x"51",
          2510 => x"0d",
          2511 => x"0c",
          2512 => x"a4",
          2513 => x"e0",
          2514 => x"3d",
          2515 => x"a4",
          2516 => x"08",
          2517 => x"a4",
          2518 => x"08",
          2519 => x"82",
          2520 => x"70",
          2521 => x"0c",
          2522 => x"0d",
          2523 => x"0c",
          2524 => x"a4",
          2525 => x"e0",
          2526 => x"3d",
          2527 => x"82",
          2528 => x"fc",
          2529 => x"e0",
          2530 => x"05",
          2531 => x"9b",
          2532 => x"a4",
          2533 => x"08",
          2534 => x"3f",
          2535 => x"08",
          2536 => x"a4",
          2537 => x"0c",
          2538 => x"82",
          2539 => x"fc",
          2540 => x"e0",
          2541 => x"05",
          2542 => x"a4",
          2543 => x"08",
          2544 => x"38",
          2545 => x"08",
          2546 => x"51",
          2547 => x"82",
          2548 => x"82",
          2549 => x"e4",
          2550 => x"31",
          2551 => x"08",
          2552 => x"52",
          2553 => x"e0",
          2554 => x"05",
          2555 => x"a4",
          2556 => x"08",
          2557 => x"a4",
          2558 => x"0c",
          2559 => x"08",
          2560 => x"82",
          2561 => x"f8",
          2562 => x"e0",
          2563 => x"05",
          2564 => x"52",
          2565 => x"a4",
          2566 => x"08",
          2567 => x"82",
          2568 => x"88",
          2569 => x"82",
          2570 => x"e8",
          2571 => x"82",
          2572 => x"e0",
          2573 => x"05",
          2574 => x"52",
          2575 => x"a4",
          2576 => x"08",
          2577 => x"06",
          2578 => x"0b",
          2579 => x"08",
          2580 => x"82",
          2581 => x"e0",
          2582 => x"05",
          2583 => x"82",
          2584 => x"f8",
          2585 => x"e0",
          2586 => x"05",
          2587 => x"a4",
          2588 => x"08",
          2589 => x"a4",
          2590 => x"0c",
          2591 => x"08",
          2592 => x"82",
          2593 => x"f8",
          2594 => x"82",
          2595 => x"88",
          2596 => x"2b",
          2597 => x"08",
          2598 => x"52",
          2599 => x"e0",
          2600 => x"05",
          2601 => x"a4",
          2602 => x"08",
          2603 => x"ab",
          2604 => x"a4",
          2605 => x"08",
          2606 => x"a4",
          2607 => x"08",
          2608 => x"e0",
          2609 => x"05",
          2610 => x"70",
          2611 => x"e0",
          2612 => x"05",
          2613 => x"a4",
          2614 => x"08",
          2615 => x"e0",
          2616 => x"05",
          2617 => x"e0",
          2618 => x"05",
          2619 => x"a4",
          2620 => x"08",
          2621 => x"08",
          2622 => x"31",
          2623 => x"e0",
          2624 => x"05",
          2625 => x"71",
          2626 => x"e0",
          2627 => x"05",
          2628 => x"a4",
          2629 => x"08",
          2630 => x"e0",
          2631 => x"05",
          2632 => x"a4",
          2633 => x"08",
          2634 => x"08",
          2635 => x"06",
          2636 => x"08",
          2637 => x"71",
          2638 => x"a4",
          2639 => x"0c",
          2640 => x"08",
          2641 => x"ff",
          2642 => x"a4",
          2643 => x"0c",
          2644 => x"51",
          2645 => x"53",
          2646 => x"82",
          2647 => x"f4",
          2648 => x"82",
          2649 => x"e8",
          2650 => x"82",
          2651 => x"e8",
          2652 => x"e0",
          2653 => x"3d",
          2654 => x"a4",
          2655 => x"e0",
          2656 => x"82",
          2657 => x"fb",
          2658 => x"0b",
          2659 => x"08",
          2660 => x"82",
          2661 => x"88",
          2662 => x"e0",
          2663 => x"05",
          2664 => x"e0",
          2665 => x"05",
          2666 => x"a4",
          2667 => x"08",
          2668 => x"08",
          2669 => x"2c",
          2670 => x"08",
          2671 => x"82",
          2672 => x"88",
          2673 => x"e0",
          2674 => x"05",
          2675 => x"82",
          2676 => x"f8",
          2677 => x"82",
          2678 => x"88",
          2679 => x"e0",
          2680 => x"05",
          2681 => x"a4",
          2682 => x"08",
          2683 => x"e0",
          2684 => x"05",
          2685 => x"e0",
          2686 => x"05",
          2687 => x"a4",
          2688 => x"08",
          2689 => x"08",
          2690 => x"32",
          2691 => x"08",
          2692 => x"82",
          2693 => x"8c",
          2694 => x"82",
          2695 => x"88",
          2696 => x"51",
          2697 => x"3f",
          2698 => x"08",
          2699 => x"a4",
          2700 => x"08",
          2701 => x"e0",
          2702 => x"05",
          2703 => x"82",
          2704 => x"51",
          2705 => x"3d",
          2706 => x"a4",
          2707 => x"e0",
          2708 => x"82",
          2709 => x"f7",
          2710 => x"0b",
          2711 => x"08",
          2712 => x"82",
          2713 => x"8c",
          2714 => x"80",
          2715 => x"e0",
          2716 => x"05",
          2717 => x"51",
          2718 => x"53",
          2719 => x"a4",
          2720 => x"34",
          2721 => x"06",
          2722 => x"2e",
          2723 => x"91",
          2724 => x"a4",
          2725 => x"08",
          2726 => x"05",
          2727 => x"ce",
          2728 => x"a4",
          2729 => x"33",
          2730 => x"2e",
          2731 => x"a4",
          2732 => x"82",
          2733 => x"f0",
          2734 => x"e0",
          2735 => x"05",
          2736 => x"81",
          2737 => x"70",
          2738 => x"72",
          2739 => x"a4",
          2740 => x"34",
          2741 => x"08",
          2742 => x"53",
          2743 => x"09",
          2744 => x"dc",
          2745 => x"a4",
          2746 => x"08",
          2747 => x"05",
          2748 => x"08",
          2749 => x"33",
          2750 => x"08",
          2751 => x"82",
          2752 => x"f8",
          2753 => x"e0",
          2754 => x"05",
          2755 => x"a4",
          2756 => x"08",
          2757 => x"b6",
          2758 => x"a4",
          2759 => x"08",
          2760 => x"84",
          2761 => x"39",
          2762 => x"e0",
          2763 => x"05",
          2764 => x"a4",
          2765 => x"08",
          2766 => x"05",
          2767 => x"08",
          2768 => x"33",
          2769 => x"08",
          2770 => x"81",
          2771 => x"0b",
          2772 => x"08",
          2773 => x"82",
          2774 => x"88",
          2775 => x"08",
          2776 => x"0c",
          2777 => x"53",
          2778 => x"e0",
          2779 => x"05",
          2780 => x"39",
          2781 => x"08",
          2782 => x"53",
          2783 => x"8d",
          2784 => x"82",
          2785 => x"ec",
          2786 => x"80",
          2787 => x"a4",
          2788 => x"33",
          2789 => x"27",
          2790 => x"e0",
          2791 => x"05",
          2792 => x"b9",
          2793 => x"8d",
          2794 => x"82",
          2795 => x"ec",
          2796 => x"d8",
          2797 => x"82",
          2798 => x"f4",
          2799 => x"39",
          2800 => x"08",
          2801 => x"53",
          2802 => x"90",
          2803 => x"a4",
          2804 => x"33",
          2805 => x"26",
          2806 => x"39",
          2807 => x"e0",
          2808 => x"05",
          2809 => x"39",
          2810 => x"e0",
          2811 => x"05",
          2812 => x"82",
          2813 => x"fc",
          2814 => x"e0",
          2815 => x"05",
          2816 => x"73",
          2817 => x"38",
          2818 => x"08",
          2819 => x"53",
          2820 => x"27",
          2821 => x"e0",
          2822 => x"05",
          2823 => x"51",
          2824 => x"e0",
          2825 => x"05",
          2826 => x"a4",
          2827 => x"33",
          2828 => x"53",
          2829 => x"a4",
          2830 => x"34",
          2831 => x"08",
          2832 => x"53",
          2833 => x"ad",
          2834 => x"a4",
          2835 => x"33",
          2836 => x"53",
          2837 => x"a4",
          2838 => x"34",
          2839 => x"08",
          2840 => x"53",
          2841 => x"8d",
          2842 => x"82",
          2843 => x"ec",
          2844 => x"98",
          2845 => x"a4",
          2846 => x"33",
          2847 => x"08",
          2848 => x"54",
          2849 => x"26",
          2850 => x"0b",
          2851 => x"08",
          2852 => x"80",
          2853 => x"e0",
          2854 => x"05",
          2855 => x"e0",
          2856 => x"05",
          2857 => x"e0",
          2858 => x"05",
          2859 => x"82",
          2860 => x"fc",
          2861 => x"e0",
          2862 => x"05",
          2863 => x"81",
          2864 => x"70",
          2865 => x"52",
          2866 => x"33",
          2867 => x"08",
          2868 => x"fe",
          2869 => x"e0",
          2870 => x"05",
          2871 => x"80",
          2872 => x"82",
          2873 => x"fc",
          2874 => x"82",
          2875 => x"fc",
          2876 => x"e0",
          2877 => x"05",
          2878 => x"a4",
          2879 => x"08",
          2880 => x"81",
          2881 => x"a4",
          2882 => x"0c",
          2883 => x"08",
          2884 => x"82",
          2885 => x"8b",
          2886 => x"e0",
          2887 => x"82",
          2888 => x"02",
          2889 => x"0c",
          2890 => x"80",
          2891 => x"a4",
          2892 => x"34",
          2893 => x"08",
          2894 => x"53",
          2895 => x"82",
          2896 => x"88",
          2897 => x"08",
          2898 => x"33",
          2899 => x"e0",
          2900 => x"05",
          2901 => x"ff",
          2902 => x"a0",
          2903 => x"06",
          2904 => x"e0",
          2905 => x"05",
          2906 => x"81",
          2907 => x"53",
          2908 => x"e0",
          2909 => x"05",
          2910 => x"ad",
          2911 => x"06",
          2912 => x"0b",
          2913 => x"08",
          2914 => x"82",
          2915 => x"88",
          2916 => x"08",
          2917 => x"0c",
          2918 => x"53",
          2919 => x"e0",
          2920 => x"05",
          2921 => x"a4",
          2922 => x"33",
          2923 => x"2e",
          2924 => x"81",
          2925 => x"e0",
          2926 => x"05",
          2927 => x"81",
          2928 => x"70",
          2929 => x"72",
          2930 => x"a4",
          2931 => x"34",
          2932 => x"08",
          2933 => x"82",
          2934 => x"e8",
          2935 => x"e0",
          2936 => x"05",
          2937 => x"2e",
          2938 => x"e0",
          2939 => x"05",
          2940 => x"2e",
          2941 => x"cd",
          2942 => x"82",
          2943 => x"f4",
          2944 => x"e0",
          2945 => x"05",
          2946 => x"81",
          2947 => x"70",
          2948 => x"72",
          2949 => x"a4",
          2950 => x"34",
          2951 => x"82",
          2952 => x"a4",
          2953 => x"34",
          2954 => x"08",
          2955 => x"70",
          2956 => x"71",
          2957 => x"51",
          2958 => x"82",
          2959 => x"f8",
          2960 => x"fe",
          2961 => x"a4",
          2962 => x"33",
          2963 => x"26",
          2964 => x"0b",
          2965 => x"08",
          2966 => x"83",
          2967 => x"e0",
          2968 => x"05",
          2969 => x"73",
          2970 => x"82",
          2971 => x"f8",
          2972 => x"72",
          2973 => x"38",
          2974 => x"0b",
          2975 => x"08",
          2976 => x"82",
          2977 => x"0b",
          2978 => x"08",
          2979 => x"b2",
          2980 => x"a4",
          2981 => x"33",
          2982 => x"27",
          2983 => x"e0",
          2984 => x"05",
          2985 => x"b9",
          2986 => x"8d",
          2987 => x"82",
          2988 => x"ec",
          2989 => x"a5",
          2990 => x"82",
          2991 => x"f4",
          2992 => x"0b",
          2993 => x"08",
          2994 => x"82",
          2995 => x"f8",
          2996 => x"a0",
          2997 => x"cf",
          2998 => x"a4",
          2999 => x"33",
          3000 => x"73",
          3001 => x"82",
          3002 => x"f8",
          3003 => x"11",
          3004 => x"82",
          3005 => x"f8",
          3006 => x"e0",
          3007 => x"05",
          3008 => x"51",
          3009 => x"e0",
          3010 => x"05",
          3011 => x"a4",
          3012 => x"33",
          3013 => x"27",
          3014 => x"e0",
          3015 => x"05",
          3016 => x"51",
          3017 => x"e0",
          3018 => x"05",
          3019 => x"a4",
          3020 => x"33",
          3021 => x"26",
          3022 => x"0b",
          3023 => x"08",
          3024 => x"81",
          3025 => x"e0",
          3026 => x"05",
          3027 => x"a4",
          3028 => x"33",
          3029 => x"74",
          3030 => x"80",
          3031 => x"a4",
          3032 => x"0c",
          3033 => x"82",
          3034 => x"f4",
          3035 => x"82",
          3036 => x"fc",
          3037 => x"82",
          3038 => x"f8",
          3039 => x"12",
          3040 => x"08",
          3041 => x"82",
          3042 => x"88",
          3043 => x"08",
          3044 => x"0c",
          3045 => x"51",
          3046 => x"72",
          3047 => x"a4",
          3048 => x"34",
          3049 => x"82",
          3050 => x"f0",
          3051 => x"72",
          3052 => x"38",
          3053 => x"08",
          3054 => x"30",
          3055 => x"08",
          3056 => x"82",
          3057 => x"8c",
          3058 => x"e0",
          3059 => x"05",
          3060 => x"53",
          3061 => x"e0",
          3062 => x"05",
          3063 => x"a4",
          3064 => x"08",
          3065 => x"0c",
          3066 => x"82",
          3067 => x"04",
          3068 => x"7a",
          3069 => x"56",
          3070 => x"80",
          3071 => x"38",
          3072 => x"15",
          3073 => x"16",
          3074 => x"d2",
          3075 => x"54",
          3076 => x"09",
          3077 => x"38",
          3078 => x"f1",
          3079 => x"76",
          3080 => x"db",
          3081 => x"08",
          3082 => x"8d",
          3083 => x"98",
          3084 => x"98",
          3085 => x"53",
          3086 => x"58",
          3087 => x"82",
          3088 => x"8b",
          3089 => x"33",
          3090 => x"2e",
          3091 => x"81",
          3092 => x"ff",
          3093 => x"98",
          3094 => x"38",
          3095 => x"82",
          3096 => x"8a",
          3097 => x"81",
          3098 => x"e0",
          3099 => x"ff",
          3100 => x"52",
          3101 => x"81",
          3102 => x"84",
          3103 => x"fc",
          3104 => x"08",
          3105 => x"e4",
          3106 => x"39",
          3107 => x"51",
          3108 => x"82",
          3109 => x"80",
          3110 => x"be",
          3111 => x"eb",
          3112 => x"a0",
          3113 => x"39",
          3114 => x"51",
          3115 => x"82",
          3116 => x"80",
          3117 => x"be",
          3118 => x"cf",
          3119 => x"ec",
          3120 => x"39",
          3121 => x"51",
          3122 => x"82",
          3123 => x"bb",
          3124 => x"b8",
          3125 => x"82",
          3126 => x"af",
          3127 => x"f4",
          3128 => x"82",
          3129 => x"a3",
          3130 => x"a4",
          3131 => x"82",
          3132 => x"97",
          3133 => x"cc",
          3134 => x"82",
          3135 => x"8b",
          3136 => x"fc",
          3137 => x"82",
          3138 => x"ce",
          3139 => x"3d",
          3140 => x"3d",
          3141 => x"56",
          3142 => x"e7",
          3143 => x"74",
          3144 => x"e8",
          3145 => x"39",
          3146 => x"74",
          3147 => x"3f",
          3148 => x"08",
          3149 => x"e3",
          3150 => x"e0",
          3151 => x"79",
          3152 => x"82",
          3153 => x"ff",
          3154 => x"87",
          3155 => x"ec",
          3156 => x"02",
          3157 => x"e3",
          3158 => x"57",
          3159 => x"30",
          3160 => x"73",
          3161 => x"59",
          3162 => x"77",
          3163 => x"83",
          3164 => x"74",
          3165 => x"81",
          3166 => x"55",
          3167 => x"81",
          3168 => x"53",
          3169 => x"3d",
          3170 => x"81",
          3171 => x"82",
          3172 => x"57",
          3173 => x"08",
          3174 => x"e0",
          3175 => x"c0",
          3176 => x"82",
          3177 => x"59",
          3178 => x"05",
          3179 => x"53",
          3180 => x"51",
          3181 => x"3f",
          3182 => x"08",
          3183 => x"98",
          3184 => x"7a",
          3185 => x"2e",
          3186 => x"19",
          3187 => x"59",
          3188 => x"3d",
          3189 => x"81",
          3190 => x"76",
          3191 => x"07",
          3192 => x"30",
          3193 => x"72",
          3194 => x"51",
          3195 => x"2e",
          3196 => x"c1",
          3197 => x"c0",
          3198 => x"52",
          3199 => x"92",
          3200 => x"75",
          3201 => x"0c",
          3202 => x"04",
          3203 => x"7c",
          3204 => x"b7",
          3205 => x"59",
          3206 => x"53",
          3207 => x"51",
          3208 => x"82",
          3209 => x"a8",
          3210 => x"2e",
          3211 => x"81",
          3212 => x"9c",
          3213 => x"f8",
          3214 => x"60",
          3215 => x"98",
          3216 => x"7e",
          3217 => x"82",
          3218 => x"58",
          3219 => x"04",
          3220 => x"98",
          3221 => x"0d",
          3222 => x"0d",
          3223 => x"02",
          3224 => x"cf",
          3225 => x"73",
          3226 => x"5f",
          3227 => x"5e",
          3228 => x"38",
          3229 => x"82",
          3230 => x"81",
          3231 => x"88",
          3232 => x"2e",
          3233 => x"58",
          3234 => x"2e",
          3235 => x"39",
          3236 => x"d2",
          3237 => x"7a",
          3238 => x"c4",
          3239 => x"ec",
          3240 => x"cc",
          3241 => x"e4",
          3242 => x"74",
          3243 => x"80",
          3244 => x"2e",
          3245 => x"a0",
          3246 => x"80",
          3247 => x"19",
          3248 => x"27",
          3249 => x"22",
          3250 => x"d0",
          3251 => x"bc",
          3252 => x"82",
          3253 => x"ff",
          3254 => x"82",
          3255 => x"c3",
          3256 => x"53",
          3257 => x"8e",
          3258 => x"52",
          3259 => x"51",
          3260 => x"3f",
          3261 => x"c1",
          3262 => x"ae",
          3263 => x"15",
          3264 => x"74",
          3265 => x"7a",
          3266 => x"72",
          3267 => x"c1",
          3268 => x"ad",
          3269 => x"39",
          3270 => x"51",
          3271 => x"3f",
          3272 => x"82",
          3273 => x"52",
          3274 => x"ba",
          3275 => x"39",
          3276 => x"51",
          3277 => x"3f",
          3278 => x"78",
          3279 => x"38",
          3280 => x"33",
          3281 => x"56",
          3282 => x"83",
          3283 => x"80",
          3284 => x"27",
          3285 => x"53",
          3286 => x"70",
          3287 => x"51",
          3288 => x"2e",
          3289 => x"80",
          3290 => x"38",
          3291 => x"08",
          3292 => x"88",
          3293 => x"fc",
          3294 => x"51",
          3295 => x"81",
          3296 => x"b6",
          3297 => x"f4",
          3298 => x"3f",
          3299 => x"1c",
          3300 => x"51",
          3301 => x"82",
          3302 => x"98",
          3303 => x"2c",
          3304 => x"a0",
          3305 => x"06",
          3306 => x"51",
          3307 => x"82",
          3308 => x"98",
          3309 => x"2c",
          3310 => x"70",
          3311 => x"32",
          3312 => x"72",
          3313 => x"07",
          3314 => x"58",
          3315 => x"57",
          3316 => x"d6",
          3317 => x"2e",
          3318 => x"7c",
          3319 => x"79",
          3320 => x"38",
          3321 => x"82",
          3322 => x"8f",
          3323 => x"fc",
          3324 => x"9b",
          3325 => x"8a",
          3326 => x"3f",
          3327 => x"52",
          3328 => x"51",
          3329 => x"3f",
          3330 => x"22",
          3331 => x"3f",
          3332 => x"54",
          3333 => x"53",
          3334 => x"33",
          3335 => x"98",
          3336 => x"e8",
          3337 => x"2e",
          3338 => x"89",
          3339 => x"0d",
          3340 => x"0d",
          3341 => x"80",
          3342 => x"f4",
          3343 => x"99",
          3344 => x"c2",
          3345 => x"d4",
          3346 => x"99",
          3347 => x"81",
          3348 => x"06",
          3349 => x"80",
          3350 => x"81",
          3351 => x"3f",
          3352 => x"51",
          3353 => x"80",
          3354 => x"3f",
          3355 => x"70",
          3356 => x"52",
          3357 => x"92",
          3358 => x"99",
          3359 => x"c2",
          3360 => x"98",
          3361 => x"98",
          3362 => x"83",
          3363 => x"06",
          3364 => x"80",
          3365 => x"81",
          3366 => x"3f",
          3367 => x"51",
          3368 => x"80",
          3369 => x"3f",
          3370 => x"70",
          3371 => x"52",
          3372 => x"92",
          3373 => x"98",
          3374 => x"c3",
          3375 => x"dc",
          3376 => x"98",
          3377 => x"85",
          3378 => x"06",
          3379 => x"80",
          3380 => x"81",
          3381 => x"3f",
          3382 => x"51",
          3383 => x"80",
          3384 => x"3f",
          3385 => x"70",
          3386 => x"52",
          3387 => x"92",
          3388 => x"98",
          3389 => x"c3",
          3390 => x"a0",
          3391 => x"97",
          3392 => x"87",
          3393 => x"06",
          3394 => x"80",
          3395 => x"81",
          3396 => x"3f",
          3397 => x"51",
          3398 => x"80",
          3399 => x"3f",
          3400 => x"70",
          3401 => x"52",
          3402 => x"92",
          3403 => x"97",
          3404 => x"c3",
          3405 => x"e4",
          3406 => x"97",
          3407 => x"f8",
          3408 => x"0d",
          3409 => x"0d",
          3410 => x"05",
          3411 => x"70",
          3412 => x"80",
          3413 => x"d9",
          3414 => x"0b",
          3415 => x"33",
          3416 => x"38",
          3417 => x"c4",
          3418 => x"f7",
          3419 => x"8b",
          3420 => x"e0",
          3421 => x"70",
          3422 => x"08",
          3423 => x"82",
          3424 => x"51",
          3425 => x"0b",
          3426 => x"34",
          3427 => x"db",
          3428 => x"73",
          3429 => x"81",
          3430 => x"82",
          3431 => x"74",
          3432 => x"81",
          3433 => x"82",
          3434 => x"80",
          3435 => x"82",
          3436 => x"51",
          3437 => x"91",
          3438 => x"a8",
          3439 => x"e7",
          3440 => x"0b",
          3441 => x"9c",
          3442 => x"82",
          3443 => x"54",
          3444 => x"09",
          3445 => x"38",
          3446 => x"53",
          3447 => x"51",
          3448 => x"80",
          3449 => x"98",
          3450 => x"0d",
          3451 => x"0d",
          3452 => x"5e",
          3453 => x"f7",
          3454 => x"81",
          3455 => x"80",
          3456 => x"82",
          3457 => x"81",
          3458 => x"78",
          3459 => x"81",
          3460 => x"97",
          3461 => x"53",
          3462 => x"52",
          3463 => x"f9",
          3464 => x"78",
          3465 => x"c4",
          3466 => x"9a",
          3467 => x"98",
          3468 => x"88",
          3469 => x"ac",
          3470 => x"39",
          3471 => x"5e",
          3472 => x"51",
          3473 => x"3f",
          3474 => x"47",
          3475 => x"52",
          3476 => x"f1",
          3477 => x"ff",
          3478 => x"f3",
          3479 => x"e0",
          3480 => x"2b",
          3481 => x"51",
          3482 => x"c2",
          3483 => x"38",
          3484 => x"24",
          3485 => x"bd",
          3486 => x"38",
          3487 => x"90",
          3488 => x"2e",
          3489 => x"78",
          3490 => x"da",
          3491 => x"39",
          3492 => x"2e",
          3493 => x"78",
          3494 => x"85",
          3495 => x"bf",
          3496 => x"38",
          3497 => x"78",
          3498 => x"89",
          3499 => x"80",
          3500 => x"38",
          3501 => x"2e",
          3502 => x"78",
          3503 => x"89",
          3504 => x"a7",
          3505 => x"83",
          3506 => x"38",
          3507 => x"24",
          3508 => x"81",
          3509 => x"f1",
          3510 => x"39",
          3511 => x"2e",
          3512 => x"8a",
          3513 => x"3d",
          3514 => x"53",
          3515 => x"51",
          3516 => x"82",
          3517 => x"80",
          3518 => x"38",
          3519 => x"fc",
          3520 => x"84",
          3521 => x"97",
          3522 => x"98",
          3523 => x"fe",
          3524 => x"3d",
          3525 => x"53",
          3526 => x"51",
          3527 => x"82",
          3528 => x"86",
          3529 => x"98",
          3530 => x"c4",
          3531 => x"a5",
          3532 => x"64",
          3533 => x"7b",
          3534 => x"38",
          3535 => x"7a",
          3536 => x"5c",
          3537 => x"26",
          3538 => x"db",
          3539 => x"ff",
          3540 => x"ff",
          3541 => x"eb",
          3542 => x"e0",
          3543 => x"2e",
          3544 => x"b5",
          3545 => x"11",
          3546 => x"05",
          3547 => x"3f",
          3548 => x"08",
          3549 => x"c8",
          3550 => x"fe",
          3551 => x"ff",
          3552 => x"eb",
          3553 => x"e0",
          3554 => x"2e",
          3555 => x"82",
          3556 => x"ff",
          3557 => x"64",
          3558 => x"27",
          3559 => x"62",
          3560 => x"81",
          3561 => x"79",
          3562 => x"05",
          3563 => x"b5",
          3564 => x"11",
          3565 => x"05",
          3566 => x"3f",
          3567 => x"08",
          3568 => x"fc",
          3569 => x"fe",
          3570 => x"ff",
          3571 => x"ea",
          3572 => x"e0",
          3573 => x"2e",
          3574 => x"b5",
          3575 => x"11",
          3576 => x"05",
          3577 => x"3f",
          3578 => x"08",
          3579 => x"d0",
          3580 => x"84",
          3581 => x"94",
          3582 => x"79",
          3583 => x"38",
          3584 => x"7b",
          3585 => x"5b",
          3586 => x"92",
          3587 => x"7a",
          3588 => x"53",
          3589 => x"c5",
          3590 => x"a3",
          3591 => x"1a",
          3592 => x"44",
          3593 => x"8a",
          3594 => x"3f",
          3595 => x"b5",
          3596 => x"11",
          3597 => x"05",
          3598 => x"3f",
          3599 => x"08",
          3600 => x"82",
          3601 => x"59",
          3602 => x"89",
          3603 => x"b4",
          3604 => x"cd",
          3605 => x"fd",
          3606 => x"80",
          3607 => x"82",
          3608 => x"45",
          3609 => x"de",
          3610 => x"78",
          3611 => x"38",
          3612 => x"08",
          3613 => x"82",
          3614 => x"59",
          3615 => x"88",
          3616 => x"cc",
          3617 => x"39",
          3618 => x"33",
          3619 => x"2e",
          3620 => x"de",
          3621 => x"89",
          3622 => x"e4",
          3623 => x"05",
          3624 => x"fe",
          3625 => x"ff",
          3626 => x"e8",
          3627 => x"e0",
          3628 => x"de",
          3629 => x"fc",
          3630 => x"80",
          3631 => x"82",
          3632 => x"44",
          3633 => x"82",
          3634 => x"59",
          3635 => x"88",
          3636 => x"c0",
          3637 => x"39",
          3638 => x"33",
          3639 => x"2e",
          3640 => x"de",
          3641 => x"aa",
          3642 => x"ff",
          3643 => x"80",
          3644 => x"82",
          3645 => x"44",
          3646 => x"de",
          3647 => x"78",
          3648 => x"38",
          3649 => x"08",
          3650 => x"82",
          3651 => x"88",
          3652 => x"3d",
          3653 => x"53",
          3654 => x"51",
          3655 => x"82",
          3656 => x"80",
          3657 => x"80",
          3658 => x"7a",
          3659 => x"38",
          3660 => x"90",
          3661 => x"70",
          3662 => x"2a",
          3663 => x"51",
          3664 => x"78",
          3665 => x"38",
          3666 => x"83",
          3667 => x"82",
          3668 => x"ff",
          3669 => x"80",
          3670 => x"62",
          3671 => x"64",
          3672 => x"3f",
          3673 => x"51",
          3674 => x"b5",
          3675 => x"11",
          3676 => x"05",
          3677 => x"3f",
          3678 => x"08",
          3679 => x"c0",
          3680 => x"fe",
          3681 => x"ff",
          3682 => x"e7",
          3683 => x"e0",
          3684 => x"2e",
          3685 => x"59",
          3686 => x"05",
          3687 => x"64",
          3688 => x"b5",
          3689 => x"11",
          3690 => x"05",
          3691 => x"3f",
          3692 => x"08",
          3693 => x"88",
          3694 => x"33",
          3695 => x"c5",
          3696 => x"a0",
          3697 => x"fb",
          3698 => x"80",
          3699 => x"51",
          3700 => x"3f",
          3701 => x"33",
          3702 => x"2e",
          3703 => x"9f",
          3704 => x"38",
          3705 => x"fc",
          3706 => x"84",
          3707 => x"af",
          3708 => x"98",
          3709 => x"91",
          3710 => x"02",
          3711 => x"33",
          3712 => x"81",
          3713 => x"b1",
          3714 => x"d4",
          3715 => x"87",
          3716 => x"39",
          3717 => x"f4",
          3718 => x"84",
          3719 => x"ae",
          3720 => x"98",
          3721 => x"f8",
          3722 => x"3d",
          3723 => x"53",
          3724 => x"51",
          3725 => x"82",
          3726 => x"80",
          3727 => x"61",
          3728 => x"c2",
          3729 => x"70",
          3730 => x"23",
          3731 => x"3d",
          3732 => x"53",
          3733 => x"51",
          3734 => x"82",
          3735 => x"df",
          3736 => x"39",
          3737 => x"54",
          3738 => x"d8",
          3739 => x"9c",
          3740 => x"f8",
          3741 => x"f8",
          3742 => x"ff",
          3743 => x"79",
          3744 => x"59",
          3745 => x"f7",
          3746 => x"9f",
          3747 => x"61",
          3748 => x"d0",
          3749 => x"fe",
          3750 => x"ff",
          3751 => x"df",
          3752 => x"e0",
          3753 => x"2e",
          3754 => x"59",
          3755 => x"05",
          3756 => x"82",
          3757 => x"78",
          3758 => x"39",
          3759 => x"51",
          3760 => x"3f",
          3761 => x"b5",
          3762 => x"11",
          3763 => x"05",
          3764 => x"3f",
          3765 => x"08",
          3766 => x"e4",
          3767 => x"fe",
          3768 => x"ff",
          3769 => x"de",
          3770 => x"e0",
          3771 => x"2e",
          3772 => x"61",
          3773 => x"61",
          3774 => x"b5",
          3775 => x"11",
          3776 => x"05",
          3777 => x"3f",
          3778 => x"08",
          3779 => x"b0",
          3780 => x"08",
          3781 => x"c5",
          3782 => x"9d",
          3783 => x"fb",
          3784 => x"80",
          3785 => x"51",
          3786 => x"3f",
          3787 => x"33",
          3788 => x"2e",
          3789 => x"9f",
          3790 => x"38",
          3791 => x"f0",
          3792 => x"84",
          3793 => x"86",
          3794 => x"98",
          3795 => x"8d",
          3796 => x"71",
          3797 => x"84",
          3798 => x"b5",
          3799 => x"d4",
          3800 => x"b3",
          3801 => x"39",
          3802 => x"80",
          3803 => x"84",
          3804 => x"ab",
          3805 => x"98",
          3806 => x"f5",
          3807 => x"52",
          3808 => x"51",
          3809 => x"3f",
          3810 => x"04",
          3811 => x"80",
          3812 => x"84",
          3813 => x"87",
          3814 => x"98",
          3815 => x"f5",
          3816 => x"52",
          3817 => x"51",
          3818 => x"3f",
          3819 => x"2d",
          3820 => x"08",
          3821 => x"88",
          3822 => x"98",
          3823 => x"c6",
          3824 => x"9c",
          3825 => x"f8",
          3826 => x"c8",
          3827 => x"c7",
          3828 => x"99",
          3829 => x"39",
          3830 => x"51",
          3831 => x"3f",
          3832 => x"a6",
          3833 => x"3f",
          3834 => x"97",
          3835 => x"78",
          3836 => x"cc",
          3837 => x"52",
          3838 => x"f1",
          3839 => x"98",
          3840 => x"e0",
          3841 => x"2e",
          3842 => x"82",
          3843 => x"46",
          3844 => x"84",
          3845 => x"cc",
          3846 => x"98",
          3847 => x"06",
          3848 => x"80",
          3849 => x"38",
          3850 => x"08",
          3851 => x"3f",
          3852 => x"08",
          3853 => x"c1",
          3854 => x"7a",
          3855 => x"38",
          3856 => x"89",
          3857 => x"2e",
          3858 => x"ca",
          3859 => x"2e",
          3860 => x"c2",
          3861 => x"f8",
          3862 => x"82",
          3863 => x"80",
          3864 => x"80",
          3865 => x"ff",
          3866 => x"ff",
          3867 => x"b8",
          3868 => x"b5",
          3869 => x"05",
          3870 => x"3f",
          3871 => x"55",
          3872 => x"54",
          3873 => x"c7",
          3874 => x"3d",
          3875 => x"51",
          3876 => x"3f",
          3877 => x"54",
          3878 => x"c7",
          3879 => x"3d",
          3880 => x"51",
          3881 => x"3f",
          3882 => x"58",
          3883 => x"57",
          3884 => x"55",
          3885 => x"80",
          3886 => x"80",
          3887 => x"3d",
          3888 => x"51",
          3889 => x"82",
          3890 => x"82",
          3891 => x"09",
          3892 => x"72",
          3893 => x"51",
          3894 => x"80",
          3895 => x"26",
          3896 => x"5a",
          3897 => x"59",
          3898 => x"8d",
          3899 => x"70",
          3900 => x"5c",
          3901 => x"c3",
          3902 => x"32",
          3903 => x"07",
          3904 => x"38",
          3905 => x"09",
          3906 => x"38",
          3907 => x"51",
          3908 => x"3f",
          3909 => x"f1",
          3910 => x"39",
          3911 => x"51",
          3912 => x"3f",
          3913 => x"f5",
          3914 => x"0b",
          3915 => x"34",
          3916 => x"8c",
          3917 => x"55",
          3918 => x"52",
          3919 => x"93",
          3920 => x"98",
          3921 => x"75",
          3922 => x"87",
          3923 => x"73",
          3924 => x"3f",
          3925 => x"98",
          3926 => x"0c",
          3927 => x"9c",
          3928 => x"55",
          3929 => x"52",
          3930 => x"e7",
          3931 => x"98",
          3932 => x"75",
          3933 => x"87",
          3934 => x"73",
          3935 => x"3f",
          3936 => x"98",
          3937 => x"0c",
          3938 => x"0b",
          3939 => x"84",
          3940 => x"83",
          3941 => x"94",
          3942 => x"82",
          3943 => x"85",
          3944 => x"02",
          3945 => x"05",
          3946 => x"82",
          3947 => x"87",
          3948 => x"13",
          3949 => x"0c",
          3950 => x"0c",
          3951 => x"3f",
          3952 => x"82",
          3953 => x"ff",
          3954 => x"82",
          3955 => x"ff",
          3956 => x"80",
          3957 => x"93",
          3958 => x"51",
          3959 => x"f0",
          3960 => x"04",
          3961 => x"76",
          3962 => x"55",
          3963 => x"54",
          3964 => x"81",
          3965 => x"33",
          3966 => x"2e",
          3967 => x"86",
          3968 => x"53",
          3969 => x"33",
          3970 => x"2e",
          3971 => x"86",
          3972 => x"53",
          3973 => x"52",
          3974 => x"09",
          3975 => x"38",
          3976 => x"12",
          3977 => x"33",
          3978 => x"a2",
          3979 => x"81",
          3980 => x"2e",
          3981 => x"ea",
          3982 => x"81",
          3983 => x"72",
          3984 => x"70",
          3985 => x"38",
          3986 => x"80",
          3987 => x"73",
          3988 => x"72",
          3989 => x"70",
          3990 => x"81",
          3991 => x"81",
          3992 => x"32",
          3993 => x"80",
          3994 => x"51",
          3995 => x"80",
          3996 => x"80",
          3997 => x"05",
          3998 => x"75",
          3999 => x"70",
          4000 => x"0c",
          4001 => x"04",
          4002 => x"76",
          4003 => x"80",
          4004 => x"86",
          4005 => x"52",
          4006 => x"b2",
          4007 => x"98",
          4008 => x"80",
          4009 => x"74",
          4010 => x"e0",
          4011 => x"3d",
          4012 => x"3d",
          4013 => x"11",
          4014 => x"52",
          4015 => x"70",
          4016 => x"98",
          4017 => x"33",
          4018 => x"82",
          4019 => x"26",
          4020 => x"84",
          4021 => x"83",
          4022 => x"26",
          4023 => x"85",
          4024 => x"84",
          4025 => x"26",
          4026 => x"86",
          4027 => x"85",
          4028 => x"26",
          4029 => x"88",
          4030 => x"86",
          4031 => x"e7",
          4032 => x"38",
          4033 => x"54",
          4034 => x"87",
          4035 => x"cc",
          4036 => x"87",
          4037 => x"0c",
          4038 => x"c0",
          4039 => x"82",
          4040 => x"c0",
          4041 => x"83",
          4042 => x"c0",
          4043 => x"84",
          4044 => x"c0",
          4045 => x"85",
          4046 => x"c0",
          4047 => x"86",
          4048 => x"c0",
          4049 => x"74",
          4050 => x"a4",
          4051 => x"c0",
          4052 => x"80",
          4053 => x"98",
          4054 => x"52",
          4055 => x"98",
          4056 => x"0d",
          4057 => x"0d",
          4058 => x"c0",
          4059 => x"81",
          4060 => x"c0",
          4061 => x"5e",
          4062 => x"87",
          4063 => x"08",
          4064 => x"1c",
          4065 => x"98",
          4066 => x"79",
          4067 => x"87",
          4068 => x"08",
          4069 => x"1c",
          4070 => x"98",
          4071 => x"79",
          4072 => x"87",
          4073 => x"08",
          4074 => x"1c",
          4075 => x"98",
          4076 => x"7b",
          4077 => x"87",
          4078 => x"08",
          4079 => x"1c",
          4080 => x"0c",
          4081 => x"ff",
          4082 => x"83",
          4083 => x"58",
          4084 => x"57",
          4085 => x"56",
          4086 => x"55",
          4087 => x"54",
          4088 => x"53",
          4089 => x"ff",
          4090 => x"c8",
          4091 => x"94",
          4092 => x"3d",
          4093 => x"3d",
          4094 => x"05",
          4095 => x"52",
          4096 => x"09",
          4097 => x"38",
          4098 => x"83",
          4099 => x"70",
          4100 => x"07",
          4101 => x"70",
          4102 => x"38",
          4103 => x"84",
          4104 => x"3f",
          4105 => x"08",
          4106 => x"98",
          4107 => x"71",
          4108 => x"81",
          4109 => x"80",
          4110 => x"2e",
          4111 => x"83",
          4112 => x"72",
          4113 => x"30",
          4114 => x"76",
          4115 => x"51",
          4116 => x"38",
          4117 => x"98",
          4118 => x"0d",
          4119 => x"0d",
          4120 => x"54",
          4121 => x"53",
          4122 => x"8a",
          4123 => x"98",
          4124 => x"70",
          4125 => x"07",
          4126 => x"54",
          4127 => x"25",
          4128 => x"82",
          4129 => x"85",
          4130 => x"fb",
          4131 => x"9f",
          4132 => x"de",
          4133 => x"81",
          4134 => x"55",
          4135 => x"94",
          4136 => x"80",
          4137 => x"87",
          4138 => x"51",
          4139 => x"96",
          4140 => x"06",
          4141 => x"70",
          4142 => x"38",
          4143 => x"70",
          4144 => x"51",
          4145 => x"72",
          4146 => x"81",
          4147 => x"70",
          4148 => x"38",
          4149 => x"70",
          4150 => x"51",
          4151 => x"38",
          4152 => x"06",
          4153 => x"94",
          4154 => x"80",
          4155 => x"87",
          4156 => x"52",
          4157 => x"74",
          4158 => x"0c",
          4159 => x"04",
          4160 => x"02",
          4161 => x"70",
          4162 => x"2a",
          4163 => x"70",
          4164 => x"34",
          4165 => x"04",
          4166 => x"02",
          4167 => x"58",
          4168 => x"09",
          4169 => x"38",
          4170 => x"51",
          4171 => x"de",
          4172 => x"81",
          4173 => x"56",
          4174 => x"84",
          4175 => x"2e",
          4176 => x"c0",
          4177 => x"72",
          4178 => x"2a",
          4179 => x"55",
          4180 => x"80",
          4181 => x"73",
          4182 => x"81",
          4183 => x"72",
          4184 => x"81",
          4185 => x"06",
          4186 => x"80",
          4187 => x"73",
          4188 => x"81",
          4189 => x"72",
          4190 => x"75",
          4191 => x"53",
          4192 => x"80",
          4193 => x"2e",
          4194 => x"c0",
          4195 => x"77",
          4196 => x"0b",
          4197 => x"0c",
          4198 => x"04",
          4199 => x"79",
          4200 => x"33",
          4201 => x"06",
          4202 => x"70",
          4203 => x"fc",
          4204 => x"ff",
          4205 => x"82",
          4206 => x"70",
          4207 => x"59",
          4208 => x"87",
          4209 => x"51",
          4210 => x"86",
          4211 => x"94",
          4212 => x"08",
          4213 => x"70",
          4214 => x"54",
          4215 => x"2e",
          4216 => x"91",
          4217 => x"06",
          4218 => x"d7",
          4219 => x"32",
          4220 => x"51",
          4221 => x"2e",
          4222 => x"93",
          4223 => x"06",
          4224 => x"ff",
          4225 => x"81",
          4226 => x"87",
          4227 => x"52",
          4228 => x"86",
          4229 => x"94",
          4230 => x"72",
          4231 => x"74",
          4232 => x"ff",
          4233 => x"57",
          4234 => x"38",
          4235 => x"98",
          4236 => x"0d",
          4237 => x"0d",
          4238 => x"33",
          4239 => x"06",
          4240 => x"c0",
          4241 => x"72",
          4242 => x"38",
          4243 => x"94",
          4244 => x"70",
          4245 => x"81",
          4246 => x"51",
          4247 => x"e2",
          4248 => x"ff",
          4249 => x"c0",
          4250 => x"70",
          4251 => x"38",
          4252 => x"90",
          4253 => x"70",
          4254 => x"82",
          4255 => x"51",
          4256 => x"04",
          4257 => x"82",
          4258 => x"81",
          4259 => x"e0",
          4260 => x"fe",
          4261 => x"de",
          4262 => x"81",
          4263 => x"53",
          4264 => x"84",
          4265 => x"2e",
          4266 => x"c0",
          4267 => x"71",
          4268 => x"2a",
          4269 => x"51",
          4270 => x"52",
          4271 => x"a0",
          4272 => x"ff",
          4273 => x"c0",
          4274 => x"70",
          4275 => x"38",
          4276 => x"90",
          4277 => x"70",
          4278 => x"98",
          4279 => x"51",
          4280 => x"98",
          4281 => x"0d",
          4282 => x"0d",
          4283 => x"80",
          4284 => x"2a",
          4285 => x"51",
          4286 => x"84",
          4287 => x"c0",
          4288 => x"82",
          4289 => x"87",
          4290 => x"08",
          4291 => x"0c",
          4292 => x"94",
          4293 => x"bc",
          4294 => x"9e",
          4295 => x"de",
          4296 => x"c0",
          4297 => x"82",
          4298 => x"87",
          4299 => x"08",
          4300 => x"0c",
          4301 => x"ac",
          4302 => x"cc",
          4303 => x"9e",
          4304 => x"de",
          4305 => x"c0",
          4306 => x"82",
          4307 => x"87",
          4308 => x"08",
          4309 => x"0c",
          4310 => x"bc",
          4311 => x"dc",
          4312 => x"9e",
          4313 => x"de",
          4314 => x"c0",
          4315 => x"82",
          4316 => x"87",
          4317 => x"08",
          4318 => x"de",
          4319 => x"c0",
          4320 => x"82",
          4321 => x"87",
          4322 => x"08",
          4323 => x"0c",
          4324 => x"8c",
          4325 => x"f4",
          4326 => x"82",
          4327 => x"80",
          4328 => x"9e",
          4329 => x"84",
          4330 => x"51",
          4331 => x"80",
          4332 => x"81",
          4333 => x"de",
          4334 => x"0b",
          4335 => x"90",
          4336 => x"80",
          4337 => x"52",
          4338 => x"2e",
          4339 => x"52",
          4340 => x"fa",
          4341 => x"87",
          4342 => x"08",
          4343 => x"0a",
          4344 => x"52",
          4345 => x"83",
          4346 => x"71",
          4347 => x"34",
          4348 => x"c0",
          4349 => x"70",
          4350 => x"06",
          4351 => x"70",
          4352 => x"38",
          4353 => x"82",
          4354 => x"80",
          4355 => x"9e",
          4356 => x"a0",
          4357 => x"51",
          4358 => x"80",
          4359 => x"81",
          4360 => x"de",
          4361 => x"0b",
          4362 => x"90",
          4363 => x"80",
          4364 => x"52",
          4365 => x"2e",
          4366 => x"52",
          4367 => x"fe",
          4368 => x"87",
          4369 => x"08",
          4370 => x"80",
          4371 => x"52",
          4372 => x"83",
          4373 => x"71",
          4374 => x"34",
          4375 => x"c0",
          4376 => x"70",
          4377 => x"06",
          4378 => x"70",
          4379 => x"38",
          4380 => x"82",
          4381 => x"80",
          4382 => x"9e",
          4383 => x"81",
          4384 => x"51",
          4385 => x"80",
          4386 => x"81",
          4387 => x"df",
          4388 => x"0b",
          4389 => x"90",
          4390 => x"c0",
          4391 => x"52",
          4392 => x"2e",
          4393 => x"52",
          4394 => x"82",
          4395 => x"87",
          4396 => x"08",
          4397 => x"06",
          4398 => x"70",
          4399 => x"38",
          4400 => x"82",
          4401 => x"87",
          4402 => x"08",
          4403 => x"06",
          4404 => x"51",
          4405 => x"82",
          4406 => x"80",
          4407 => x"9e",
          4408 => x"84",
          4409 => x"52",
          4410 => x"2e",
          4411 => x"52",
          4412 => x"85",
          4413 => x"9e",
          4414 => x"83",
          4415 => x"84",
          4416 => x"51",
          4417 => x"86",
          4418 => x"87",
          4419 => x"08",
          4420 => x"51",
          4421 => x"80",
          4422 => x"81",
          4423 => x"df",
          4424 => x"c0",
          4425 => x"70",
          4426 => x"51",
          4427 => x"88",
          4428 => x"0d",
          4429 => x"0d",
          4430 => x"51",
          4431 => x"3f",
          4432 => x"33",
          4433 => x"2e",
          4434 => x"c8",
          4435 => x"89",
          4436 => x"c8",
          4437 => x"a5",
          4438 => x"de",
          4439 => x"73",
          4440 => x"38",
          4441 => x"08",
          4442 => x"08",
          4443 => x"82",
          4444 => x"ff",
          4445 => x"82",
          4446 => x"54",
          4447 => x"94",
          4448 => x"cc",
          4449 => x"d0",
          4450 => x"52",
          4451 => x"51",
          4452 => x"3f",
          4453 => x"33",
          4454 => x"2e",
          4455 => x"de",
          4456 => x"de",
          4457 => x"54",
          4458 => x"94",
          4459 => x"dc",
          4460 => x"fd",
          4461 => x"80",
          4462 => x"82",
          4463 => x"82",
          4464 => x"11",
          4465 => x"c9",
          4466 => x"88",
          4467 => x"de",
          4468 => x"73",
          4469 => x"38",
          4470 => x"08",
          4471 => x"08",
          4472 => x"82",
          4473 => x"ff",
          4474 => x"82",
          4475 => x"54",
          4476 => x"8e",
          4477 => x"84",
          4478 => x"c9",
          4479 => x"88",
          4480 => x"df",
          4481 => x"73",
          4482 => x"38",
          4483 => x"33",
          4484 => x"88",
          4485 => x"f4",
          4486 => x"85",
          4487 => x"80",
          4488 => x"82",
          4489 => x"52",
          4490 => x"51",
          4491 => x"3f",
          4492 => x"33",
          4493 => x"2e",
          4494 => x"ca",
          4495 => x"a3",
          4496 => x"de",
          4497 => x"73",
          4498 => x"38",
          4499 => x"51",
          4500 => x"3f",
          4501 => x"33",
          4502 => x"2e",
          4503 => x"ca",
          4504 => x"a3",
          4505 => x"df",
          4506 => x"73",
          4507 => x"38",
          4508 => x"51",
          4509 => x"3f",
          4510 => x"33",
          4511 => x"2e",
          4512 => x"ca",
          4513 => x"a3",
          4514 => x"cb",
          4515 => x"a3",
          4516 => x"de",
          4517 => x"82",
          4518 => x"ff",
          4519 => x"82",
          4520 => x"52",
          4521 => x"51",
          4522 => x"3f",
          4523 => x"08",
          4524 => x"e0",
          4525 => x"d4",
          4526 => x"88",
          4527 => x"d7",
          4528 => x"e8",
          4529 => x"cc",
          4530 => x"86",
          4531 => x"de",
          4532 => x"bd",
          4533 => x"75",
          4534 => x"f7",
          4535 => x"98",
          4536 => x"c0",
          4537 => x"31",
          4538 => x"e0",
          4539 => x"82",
          4540 => x"ff",
          4541 => x"82",
          4542 => x"54",
          4543 => x"aa",
          4544 => x"f0",
          4545 => x"84",
          4546 => x"51",
          4547 => x"3f",
          4548 => x"08",
          4549 => x"29",
          4550 => x"54",
          4551 => x"98",
          4552 => x"cc",
          4553 => x"85",
          4554 => x"de",
          4555 => x"73",
          4556 => x"38",
          4557 => x"08",
          4558 => x"c0",
          4559 => x"ff",
          4560 => x"82",
          4561 => x"bd",
          4562 => x"76",
          4563 => x"54",
          4564 => x"08",
          4565 => x"90",
          4566 => x"b0",
          4567 => x"ff",
          4568 => x"87",
          4569 => x"fe",
          4570 => x"92",
          4571 => x"05",
          4572 => x"26",
          4573 => x"84",
          4574 => x"cc",
          4575 => x"08",
          4576 => x"bc",
          4577 => x"82",
          4578 => x"97",
          4579 => x"cc",
          4580 => x"82",
          4581 => x"8b",
          4582 => x"d8",
          4583 => x"82",
          4584 => x"ff",
          4585 => x"84",
          4586 => x"71",
          4587 => x"04",
          4588 => x"c0",
          4589 => x"04",
          4590 => x"08",
          4591 => x"84",
          4592 => x"3d",
          4593 => x"2b",
          4594 => x"79",
          4595 => x"98",
          4596 => x"13",
          4597 => x"51",
          4598 => x"51",
          4599 => x"82",
          4600 => x"33",
          4601 => x"74",
          4602 => x"82",
          4603 => x"08",
          4604 => x"05",
          4605 => x"71",
          4606 => x"52",
          4607 => x"09",
          4608 => x"38",
          4609 => x"82",
          4610 => x"85",
          4611 => x"fb",
          4612 => x"02",
          4613 => x"05",
          4614 => x"55",
          4615 => x"80",
          4616 => x"82",
          4617 => x"52",
          4618 => x"a3",
          4619 => x"fb",
          4620 => x"a0",
          4621 => x"ae",
          4622 => x"fc",
          4623 => x"51",
          4624 => x"3f",
          4625 => x"05",
          4626 => x"34",
          4627 => x"06",
          4628 => x"77",
          4629 => x"b4",
          4630 => x"34",
          4631 => x"04",
          4632 => x"7c",
          4633 => x"b7",
          4634 => x"88",
          4635 => x"33",
          4636 => x"33",
          4637 => x"82",
          4638 => x"70",
          4639 => x"59",
          4640 => x"74",
          4641 => x"38",
          4642 => x"fd",
          4643 => x"e8",
          4644 => x"29",
          4645 => x"05",
          4646 => x"54",
          4647 => x"9d",
          4648 => x"e0",
          4649 => x"0c",
          4650 => x"33",
          4651 => x"82",
          4652 => x"70",
          4653 => x"5a",
          4654 => x"a7",
          4655 => x"78",
          4656 => x"ff",
          4657 => x"82",
          4658 => x"81",
          4659 => x"82",
          4660 => x"74",
          4661 => x"55",
          4662 => x"87",
          4663 => x"82",
          4664 => x"77",
          4665 => x"38",
          4666 => x"08",
          4667 => x"2e",
          4668 => x"df",
          4669 => x"74",
          4670 => x"3d",
          4671 => x"76",
          4672 => x"75",
          4673 => x"84",
          4674 => x"e4",
          4675 => x"51",
          4676 => x"3f",
          4677 => x"08",
          4678 => x"e8",
          4679 => x"0d",
          4680 => x"0d",
          4681 => x"53",
          4682 => x"08",
          4683 => x"2e",
          4684 => x"51",
          4685 => x"80",
          4686 => x"14",
          4687 => x"54",
          4688 => x"e6",
          4689 => x"82",
          4690 => x"82",
          4691 => x"52",
          4692 => x"95",
          4693 => x"80",
          4694 => x"82",
          4695 => x"51",
          4696 => x"80",
          4697 => x"e4",
          4698 => x"0d",
          4699 => x"0d",
          4700 => x"52",
          4701 => x"08",
          4702 => x"e9",
          4703 => x"98",
          4704 => x"38",
          4705 => x"08",
          4706 => x"52",
          4707 => x"52",
          4708 => x"c1",
          4709 => x"98",
          4710 => x"ba",
          4711 => x"ff",
          4712 => x"82",
          4713 => x"55",
          4714 => x"e0",
          4715 => x"9d",
          4716 => x"98",
          4717 => x"70",
          4718 => x"80",
          4719 => x"53",
          4720 => x"17",
          4721 => x"52",
          4722 => x"c0",
          4723 => x"2e",
          4724 => x"ff",
          4725 => x"3d",
          4726 => x"3d",
          4727 => x"08",
          4728 => x"5a",
          4729 => x"58",
          4730 => x"82",
          4731 => x"51",
          4732 => x"3f",
          4733 => x"08",
          4734 => x"ff",
          4735 => x"e4",
          4736 => x"80",
          4737 => x"3d",
          4738 => x"81",
          4739 => x"82",
          4740 => x"80",
          4741 => x"75",
          4742 => x"9d",
          4743 => x"98",
          4744 => x"58",
          4745 => x"82",
          4746 => x"25",
          4747 => x"e0",
          4748 => x"05",
          4749 => x"55",
          4750 => x"74",
          4751 => x"70",
          4752 => x"2a",
          4753 => x"78",
          4754 => x"38",
          4755 => x"38",
          4756 => x"08",
          4757 => x"53",
          4758 => x"89",
          4759 => x"98",
          4760 => x"89",
          4761 => x"e8",
          4762 => x"a0",
          4763 => x"2e",
          4764 => x"9b",
          4765 => x"79",
          4766 => x"ab",
          4767 => x"ff",
          4768 => x"ab",
          4769 => x"82",
          4770 => x"74",
          4771 => x"77",
          4772 => x"0c",
          4773 => x"04",
          4774 => x"7c",
          4775 => x"71",
          4776 => x"59",
          4777 => x"a0",
          4778 => x"06",
          4779 => x"33",
          4780 => x"77",
          4781 => x"38",
          4782 => x"5b",
          4783 => x"56",
          4784 => x"a0",
          4785 => x"06",
          4786 => x"75",
          4787 => x"80",
          4788 => x"29",
          4789 => x"05",
          4790 => x"55",
          4791 => x"3f",
          4792 => x"08",
          4793 => x"74",
          4794 => x"a9",
          4795 => x"e0",
          4796 => x"c5",
          4797 => x"33",
          4798 => x"2e",
          4799 => x"82",
          4800 => x"b5",
          4801 => x"3f",
          4802 => x"1a",
          4803 => x"fc",
          4804 => x"05",
          4805 => x"3f",
          4806 => x"08",
          4807 => x"38",
          4808 => x"78",
          4809 => x"fd",
          4810 => x"e0",
          4811 => x"ff",
          4812 => x"85",
          4813 => x"91",
          4814 => x"70",
          4815 => x"51",
          4816 => x"27",
          4817 => x"80",
          4818 => x"e0",
          4819 => x"3d",
          4820 => x"3d",
          4821 => x"08",
          4822 => x"b4",
          4823 => x"5f",
          4824 => x"af",
          4825 => x"df",
          4826 => x"df",
          4827 => x"5b",
          4828 => x"38",
          4829 => x"e0",
          4830 => x"73",
          4831 => x"55",
          4832 => x"81",
          4833 => x"70",
          4834 => x"56",
          4835 => x"81",
          4836 => x"51",
          4837 => x"82",
          4838 => x"82",
          4839 => x"82",
          4840 => x"80",
          4841 => x"38",
          4842 => x"52",
          4843 => x"08",
          4844 => x"f3",
          4845 => x"98",
          4846 => x"8c",
          4847 => x"94",
          4848 => x"d3",
          4849 => x"39",
          4850 => x"08",
          4851 => x"e4",
          4852 => x"f8",
          4853 => x"70",
          4854 => x"9a",
          4855 => x"e0",
          4856 => x"82",
          4857 => x"74",
          4858 => x"06",
          4859 => x"82",
          4860 => x"51",
          4861 => x"3f",
          4862 => x"08",
          4863 => x"82",
          4864 => x"25",
          4865 => x"e0",
          4866 => x"05",
          4867 => x"55",
          4868 => x"80",
          4869 => x"ff",
          4870 => x"51",
          4871 => x"81",
          4872 => x"ff",
          4873 => x"93",
          4874 => x"38",
          4875 => x"ff",
          4876 => x"06",
          4877 => x"86",
          4878 => x"df",
          4879 => x"8c",
          4880 => x"e4",
          4881 => x"84",
          4882 => x"3f",
          4883 => x"80",
          4884 => x"3f",
          4885 => x"08",
          4886 => x"98",
          4887 => x"78",
          4888 => x"38",
          4889 => x"06",
          4890 => x"33",
          4891 => x"70",
          4892 => x"f7",
          4893 => x"98",
          4894 => x"2c",
          4895 => x"05",
          4896 => x"82",
          4897 => x"70",
          4898 => x"33",
          4899 => x"51",
          4900 => x"59",
          4901 => x"56",
          4902 => x"80",
          4903 => x"74",
          4904 => x"74",
          4905 => x"29",
          4906 => x"05",
          4907 => x"51",
          4908 => x"24",
          4909 => x"76",
          4910 => x"77",
          4911 => x"3f",
          4912 => x"08",
          4913 => x"54",
          4914 => x"d7",
          4915 => x"f7",
          4916 => x"56",
          4917 => x"81",
          4918 => x"81",
          4919 => x"70",
          4920 => x"81",
          4921 => x"51",
          4922 => x"26",
          4923 => x"53",
          4924 => x"51",
          4925 => x"82",
          4926 => x"81",
          4927 => x"73",
          4928 => x"39",
          4929 => x"80",
          4930 => x"38",
          4931 => x"74",
          4932 => x"34",
          4933 => x"70",
          4934 => x"f7",
          4935 => x"98",
          4936 => x"2c",
          4937 => x"70",
          4938 => x"cd",
          4939 => x"5e",
          4940 => x"57",
          4941 => x"74",
          4942 => x"81",
          4943 => x"38",
          4944 => x"14",
          4945 => x"80",
          4946 => x"d4",
          4947 => x"82",
          4948 => x"92",
          4949 => x"f7",
          4950 => x"82",
          4951 => x"78",
          4952 => x"75",
          4953 => x"54",
          4954 => x"fd",
          4955 => x"84",
          4956 => x"e0",
          4957 => x"08",
          4958 => x"dc",
          4959 => x"7e",
          4960 => x"38",
          4961 => x"33",
          4962 => x"27",
          4963 => x"98",
          4964 => x"2c",
          4965 => x"75",
          4966 => x"74",
          4967 => x"33",
          4968 => x"74",
          4969 => x"29",
          4970 => x"05",
          4971 => x"82",
          4972 => x"56",
          4973 => x"39",
          4974 => x"33",
          4975 => x"54",
          4976 => x"dc",
          4977 => x"54",
          4978 => x"74",
          4979 => x"d8",
          4980 => x"7e",
          4981 => x"81",
          4982 => x"82",
          4983 => x"82",
          4984 => x"70",
          4985 => x"29",
          4986 => x"05",
          4987 => x"82",
          4988 => x"5a",
          4989 => x"74",
          4990 => x"38",
          4991 => x"08",
          4992 => x"70",
          4993 => x"ff",
          4994 => x"74",
          4995 => x"29",
          4996 => x"05",
          4997 => x"82",
          4998 => x"56",
          4999 => x"75",
          5000 => x"82",
          5001 => x"70",
          5002 => x"98",
          5003 => x"d8",
          5004 => x"56",
          5005 => x"25",
          5006 => x"82",
          5007 => x"52",
          5008 => x"97",
          5009 => x"81",
          5010 => x"81",
          5011 => x"70",
          5012 => x"f7",
          5013 => x"51",
          5014 => x"24",
          5015 => x"ec",
          5016 => x"34",
          5017 => x"1b",
          5018 => x"dc",
          5019 => x"82",
          5020 => x"f3",
          5021 => x"fd",
          5022 => x"dc",
          5023 => x"ff",
          5024 => x"73",
          5025 => x"c4",
          5026 => x"d8",
          5027 => x"54",
          5028 => x"d8",
          5029 => x"54",
          5030 => x"dc",
          5031 => x"fc",
          5032 => x"51",
          5033 => x"3f",
          5034 => x"33",
          5035 => x"70",
          5036 => x"f7",
          5037 => x"51",
          5038 => x"74",
          5039 => x"74",
          5040 => x"14",
          5041 => x"82",
          5042 => x"52",
          5043 => x"ff",
          5044 => x"74",
          5045 => x"29",
          5046 => x"05",
          5047 => x"82",
          5048 => x"58",
          5049 => x"75",
          5050 => x"82",
          5051 => x"52",
          5052 => x"95",
          5053 => x"f7",
          5054 => x"98",
          5055 => x"2c",
          5056 => x"33",
          5057 => x"57",
          5058 => x"fa",
          5059 => x"fb",
          5060 => x"88",
          5061 => x"ce",
          5062 => x"80",
          5063 => x"80",
          5064 => x"98",
          5065 => x"d8",
          5066 => x"55",
          5067 => x"de",
          5068 => x"39",
          5069 => x"33",
          5070 => x"80",
          5071 => x"fb",
          5072 => x"8a",
          5073 => x"9e",
          5074 => x"d8",
          5075 => x"f6",
          5076 => x"e0",
          5077 => x"ff",
          5078 => x"96",
          5079 => x"d8",
          5080 => x"80",
          5081 => x"81",
          5082 => x"79",
          5083 => x"3f",
          5084 => x"7a",
          5085 => x"82",
          5086 => x"80",
          5087 => x"d8",
          5088 => x"e0",
          5089 => x"3d",
          5090 => x"f7",
          5091 => x"73",
          5092 => x"b8",
          5093 => x"fc",
          5094 => x"51",
          5095 => x"3f",
          5096 => x"33",
          5097 => x"73",
          5098 => x"34",
          5099 => x"06",
          5100 => x"82",
          5101 => x"82",
          5102 => x"55",
          5103 => x"2e",
          5104 => x"ff",
          5105 => x"82",
          5106 => x"74",
          5107 => x"98",
          5108 => x"ff",
          5109 => x"55",
          5110 => x"ad",
          5111 => x"54",
          5112 => x"74",
          5113 => x"fc",
          5114 => x"33",
          5115 => x"f6",
          5116 => x"80",
          5117 => x"80",
          5118 => x"98",
          5119 => x"d8",
          5120 => x"55",
          5121 => x"d5",
          5122 => x"fc",
          5123 => x"51",
          5124 => x"3f",
          5125 => x"33",
          5126 => x"70",
          5127 => x"f7",
          5128 => x"51",
          5129 => x"74",
          5130 => x"38",
          5131 => x"08",
          5132 => x"ff",
          5133 => x"74",
          5134 => x"29",
          5135 => x"05",
          5136 => x"82",
          5137 => x"58",
          5138 => x"75",
          5139 => x"f7",
          5140 => x"f7",
          5141 => x"81",
          5142 => x"f7",
          5143 => x"56",
          5144 => x"27",
          5145 => x"82",
          5146 => x"52",
          5147 => x"73",
          5148 => x"34",
          5149 => x"33",
          5150 => x"92",
          5151 => x"f7",
          5152 => x"81",
          5153 => x"f7",
          5154 => x"56",
          5155 => x"26",
          5156 => x"b8",
          5157 => x"dc",
          5158 => x"82",
          5159 => x"ee",
          5160 => x"0b",
          5161 => x"34",
          5162 => x"f7",
          5163 => x"9c",
          5164 => x"38",
          5165 => x"08",
          5166 => x"2e",
          5167 => x"51",
          5168 => x"3f",
          5169 => x"08",
          5170 => x"34",
          5171 => x"08",
          5172 => x"81",
          5173 => x"52",
          5174 => x"9c",
          5175 => x"5b",
          5176 => x"7a",
          5177 => x"df",
          5178 => x"11",
          5179 => x"74",
          5180 => x"38",
          5181 => x"9a",
          5182 => x"e0",
          5183 => x"f7",
          5184 => x"e0",
          5185 => x"ff",
          5186 => x"53",
          5187 => x"51",
          5188 => x"3f",
          5189 => x"80",
          5190 => x"08",
          5191 => x"2e",
          5192 => x"74",
          5193 => x"91",
          5194 => x"7a",
          5195 => x"81",
          5196 => x"82",
          5197 => x"55",
          5198 => x"a4",
          5199 => x"ff",
          5200 => x"82",
          5201 => x"82",
          5202 => x"82",
          5203 => x"81",
          5204 => x"05",
          5205 => x"79",
          5206 => x"bd",
          5207 => x"39",
          5208 => x"82",
          5209 => x"70",
          5210 => x"74",
          5211 => x"38",
          5212 => x"99",
          5213 => x"e0",
          5214 => x"f7",
          5215 => x"e0",
          5216 => x"ff",
          5217 => x"53",
          5218 => x"51",
          5219 => x"3f",
          5220 => x"73",
          5221 => x"5b",
          5222 => x"82",
          5223 => x"74",
          5224 => x"f7",
          5225 => x"f7",
          5226 => x"79",
          5227 => x"3f",
          5228 => x"82",
          5229 => x"70",
          5230 => x"82",
          5231 => x"59",
          5232 => x"77",
          5233 => x"38",
          5234 => x"08",
          5235 => x"54",
          5236 => x"dc",
          5237 => x"70",
          5238 => x"ff",
          5239 => x"f4",
          5240 => x"f7",
          5241 => x"73",
          5242 => x"e0",
          5243 => x"fc",
          5244 => x"51",
          5245 => x"3f",
          5246 => x"33",
          5247 => x"73",
          5248 => x"34",
          5249 => x"f9",
          5250 => x"fa",
          5251 => x"e0",
          5252 => x"80",
          5253 => x"84",
          5254 => x"80",
          5255 => x"84",
          5256 => x"ff",
          5257 => x"82",
          5258 => x"54",
          5259 => x"74",
          5260 => x"76",
          5261 => x"82",
          5262 => x"54",
          5263 => x"34",
          5264 => x"34",
          5265 => x"08",
          5266 => x"15",
          5267 => x"15",
          5268 => x"88",
          5269 => x"84",
          5270 => x"fe",
          5271 => x"70",
          5272 => x"06",
          5273 => x"58",
          5274 => x"74",
          5275 => x"73",
          5276 => x"82",
          5277 => x"70",
          5278 => x"e0",
          5279 => x"f8",
          5280 => x"55",
          5281 => x"34",
          5282 => x"34",
          5283 => x"04",
          5284 => x"73",
          5285 => x"84",
          5286 => x"38",
          5287 => x"2a",
          5288 => x"83",
          5289 => x"51",
          5290 => x"82",
          5291 => x"83",
          5292 => x"f9",
          5293 => x"a6",
          5294 => x"84",
          5295 => x"22",
          5296 => x"e0",
          5297 => x"83",
          5298 => x"74",
          5299 => x"11",
          5300 => x"12",
          5301 => x"2b",
          5302 => x"05",
          5303 => x"71",
          5304 => x"06",
          5305 => x"2a",
          5306 => x"59",
          5307 => x"57",
          5308 => x"71",
          5309 => x"81",
          5310 => x"e0",
          5311 => x"75",
          5312 => x"54",
          5313 => x"34",
          5314 => x"34",
          5315 => x"08",
          5316 => x"33",
          5317 => x"71",
          5318 => x"70",
          5319 => x"ff",
          5320 => x"52",
          5321 => x"05",
          5322 => x"ff",
          5323 => x"2a",
          5324 => x"71",
          5325 => x"72",
          5326 => x"53",
          5327 => x"34",
          5328 => x"08",
          5329 => x"76",
          5330 => x"17",
          5331 => x"0d",
          5332 => x"0d",
          5333 => x"08",
          5334 => x"9e",
          5335 => x"83",
          5336 => x"86",
          5337 => x"12",
          5338 => x"2b",
          5339 => x"07",
          5340 => x"52",
          5341 => x"05",
          5342 => x"85",
          5343 => x"88",
          5344 => x"88",
          5345 => x"56",
          5346 => x"13",
          5347 => x"13",
          5348 => x"88",
          5349 => x"84",
          5350 => x"12",
          5351 => x"2b",
          5352 => x"07",
          5353 => x"52",
          5354 => x"12",
          5355 => x"33",
          5356 => x"07",
          5357 => x"54",
          5358 => x"70",
          5359 => x"73",
          5360 => x"82",
          5361 => x"13",
          5362 => x"12",
          5363 => x"2b",
          5364 => x"ff",
          5365 => x"88",
          5366 => x"53",
          5367 => x"73",
          5368 => x"14",
          5369 => x"0d",
          5370 => x"0d",
          5371 => x"22",
          5372 => x"08",
          5373 => x"71",
          5374 => x"81",
          5375 => x"88",
          5376 => x"88",
          5377 => x"33",
          5378 => x"71",
          5379 => x"90",
          5380 => x"5f",
          5381 => x"5a",
          5382 => x"54",
          5383 => x"80",
          5384 => x"51",
          5385 => x"82",
          5386 => x"70",
          5387 => x"81",
          5388 => x"8b",
          5389 => x"2b",
          5390 => x"70",
          5391 => x"33",
          5392 => x"07",
          5393 => x"8f",
          5394 => x"51",
          5395 => x"53",
          5396 => x"72",
          5397 => x"2a",
          5398 => x"82",
          5399 => x"83",
          5400 => x"e0",
          5401 => x"16",
          5402 => x"12",
          5403 => x"2b",
          5404 => x"07",
          5405 => x"55",
          5406 => x"33",
          5407 => x"71",
          5408 => x"70",
          5409 => x"06",
          5410 => x"57",
          5411 => x"52",
          5412 => x"71",
          5413 => x"88",
          5414 => x"fb",
          5415 => x"e0",
          5416 => x"84",
          5417 => x"22",
          5418 => x"72",
          5419 => x"33",
          5420 => x"71",
          5421 => x"83",
          5422 => x"5b",
          5423 => x"52",
          5424 => x"33",
          5425 => x"71",
          5426 => x"02",
          5427 => x"05",
          5428 => x"70",
          5429 => x"51",
          5430 => x"71",
          5431 => x"81",
          5432 => x"e0",
          5433 => x"15",
          5434 => x"12",
          5435 => x"2b",
          5436 => x"07",
          5437 => x"52",
          5438 => x"12",
          5439 => x"33",
          5440 => x"07",
          5441 => x"54",
          5442 => x"70",
          5443 => x"72",
          5444 => x"82",
          5445 => x"14",
          5446 => x"83",
          5447 => x"88",
          5448 => x"e0",
          5449 => x"54",
          5450 => x"04",
          5451 => x"7b",
          5452 => x"08",
          5453 => x"70",
          5454 => x"06",
          5455 => x"53",
          5456 => x"82",
          5457 => x"76",
          5458 => x"11",
          5459 => x"83",
          5460 => x"8b",
          5461 => x"2b",
          5462 => x"70",
          5463 => x"33",
          5464 => x"71",
          5465 => x"53",
          5466 => x"53",
          5467 => x"59",
          5468 => x"25",
          5469 => x"80",
          5470 => x"51",
          5471 => x"81",
          5472 => x"14",
          5473 => x"33",
          5474 => x"71",
          5475 => x"76",
          5476 => x"2a",
          5477 => x"58",
          5478 => x"14",
          5479 => x"ff",
          5480 => x"87",
          5481 => x"e0",
          5482 => x"19",
          5483 => x"85",
          5484 => x"88",
          5485 => x"88",
          5486 => x"5b",
          5487 => x"84",
          5488 => x"85",
          5489 => x"e0",
          5490 => x"53",
          5491 => x"14",
          5492 => x"87",
          5493 => x"e0",
          5494 => x"76",
          5495 => x"75",
          5496 => x"82",
          5497 => x"18",
          5498 => x"12",
          5499 => x"2b",
          5500 => x"80",
          5501 => x"88",
          5502 => x"55",
          5503 => x"74",
          5504 => x"15",
          5505 => x"0d",
          5506 => x"0d",
          5507 => x"e0",
          5508 => x"38",
          5509 => x"71",
          5510 => x"38",
          5511 => x"8c",
          5512 => x"0d",
          5513 => x"0d",
          5514 => x"58",
          5515 => x"82",
          5516 => x"83",
          5517 => x"82",
          5518 => x"84",
          5519 => x"12",
          5520 => x"2b",
          5521 => x"59",
          5522 => x"81",
          5523 => x"75",
          5524 => x"cb",
          5525 => x"29",
          5526 => x"81",
          5527 => x"88",
          5528 => x"81",
          5529 => x"79",
          5530 => x"ff",
          5531 => x"7f",
          5532 => x"51",
          5533 => x"77",
          5534 => x"38",
          5535 => x"85",
          5536 => x"5a",
          5537 => x"33",
          5538 => x"71",
          5539 => x"57",
          5540 => x"38",
          5541 => x"ff",
          5542 => x"7a",
          5543 => x"80",
          5544 => x"82",
          5545 => x"11",
          5546 => x"12",
          5547 => x"2b",
          5548 => x"ff",
          5549 => x"52",
          5550 => x"55",
          5551 => x"83",
          5552 => x"80",
          5553 => x"26",
          5554 => x"74",
          5555 => x"2e",
          5556 => x"77",
          5557 => x"81",
          5558 => x"75",
          5559 => x"3f",
          5560 => x"82",
          5561 => x"79",
          5562 => x"f7",
          5563 => x"e0",
          5564 => x"1c",
          5565 => x"87",
          5566 => x"8b",
          5567 => x"2b",
          5568 => x"5e",
          5569 => x"7a",
          5570 => x"ff",
          5571 => x"88",
          5572 => x"56",
          5573 => x"15",
          5574 => x"ff",
          5575 => x"85",
          5576 => x"e0",
          5577 => x"83",
          5578 => x"72",
          5579 => x"33",
          5580 => x"71",
          5581 => x"70",
          5582 => x"5b",
          5583 => x"56",
          5584 => x"19",
          5585 => x"19",
          5586 => x"88",
          5587 => x"84",
          5588 => x"12",
          5589 => x"2b",
          5590 => x"07",
          5591 => x"55",
          5592 => x"78",
          5593 => x"76",
          5594 => x"82",
          5595 => x"70",
          5596 => x"84",
          5597 => x"12",
          5598 => x"2b",
          5599 => x"2a",
          5600 => x"52",
          5601 => x"84",
          5602 => x"85",
          5603 => x"e0",
          5604 => x"84",
          5605 => x"82",
          5606 => x"8d",
          5607 => x"fe",
          5608 => x"52",
          5609 => x"08",
          5610 => x"db",
          5611 => x"71",
          5612 => x"38",
          5613 => x"ed",
          5614 => x"98",
          5615 => x"82",
          5616 => x"84",
          5617 => x"ee",
          5618 => x"66",
          5619 => x"70",
          5620 => x"e0",
          5621 => x"2e",
          5622 => x"84",
          5623 => x"3f",
          5624 => x"7e",
          5625 => x"3f",
          5626 => x"08",
          5627 => x"39",
          5628 => x"7b",
          5629 => x"3f",
          5630 => x"ba",
          5631 => x"f5",
          5632 => x"e0",
          5633 => x"ff",
          5634 => x"e0",
          5635 => x"71",
          5636 => x"70",
          5637 => x"06",
          5638 => x"73",
          5639 => x"81",
          5640 => x"88",
          5641 => x"75",
          5642 => x"ff",
          5643 => x"88",
          5644 => x"73",
          5645 => x"70",
          5646 => x"33",
          5647 => x"07",
          5648 => x"53",
          5649 => x"48",
          5650 => x"54",
          5651 => x"56",
          5652 => x"80",
          5653 => x"76",
          5654 => x"06",
          5655 => x"83",
          5656 => x"42",
          5657 => x"33",
          5658 => x"71",
          5659 => x"70",
          5660 => x"70",
          5661 => x"33",
          5662 => x"71",
          5663 => x"53",
          5664 => x"56",
          5665 => x"25",
          5666 => x"75",
          5667 => x"ff",
          5668 => x"54",
          5669 => x"81",
          5670 => x"18",
          5671 => x"2e",
          5672 => x"8f",
          5673 => x"f6",
          5674 => x"83",
          5675 => x"58",
          5676 => x"7f",
          5677 => x"74",
          5678 => x"78",
          5679 => x"3f",
          5680 => x"7f",
          5681 => x"75",
          5682 => x"38",
          5683 => x"11",
          5684 => x"33",
          5685 => x"07",
          5686 => x"f4",
          5687 => x"52",
          5688 => x"b7",
          5689 => x"98",
          5690 => x"ff",
          5691 => x"7c",
          5692 => x"2b",
          5693 => x"08",
          5694 => x"53",
          5695 => x"87",
          5696 => x"e0",
          5697 => x"84",
          5698 => x"ff",
          5699 => x"5c",
          5700 => x"60",
          5701 => x"74",
          5702 => x"38",
          5703 => x"c9",
          5704 => x"88",
          5705 => x"11",
          5706 => x"33",
          5707 => x"07",
          5708 => x"f4",
          5709 => x"52",
          5710 => x"df",
          5711 => x"98",
          5712 => x"ff",
          5713 => x"7c",
          5714 => x"2b",
          5715 => x"08",
          5716 => x"53",
          5717 => x"86",
          5718 => x"e0",
          5719 => x"84",
          5720 => x"05",
          5721 => x"73",
          5722 => x"06",
          5723 => x"7b",
          5724 => x"f9",
          5725 => x"e0",
          5726 => x"82",
          5727 => x"80",
          5728 => x"7d",
          5729 => x"82",
          5730 => x"51",
          5731 => x"3f",
          5732 => x"98",
          5733 => x"7a",
          5734 => x"38",
          5735 => x"52",
          5736 => x"8f",
          5737 => x"83",
          5738 => x"88",
          5739 => x"05",
          5740 => x"3f",
          5741 => x"82",
          5742 => x"94",
          5743 => x"fc",
          5744 => x"77",
          5745 => x"54",
          5746 => x"82",
          5747 => x"55",
          5748 => x"08",
          5749 => x"38",
          5750 => x"52",
          5751 => x"08",
          5752 => x"e1",
          5753 => x"e0",
          5754 => x"3d",
          5755 => x"3d",
          5756 => x"05",
          5757 => x"52",
          5758 => x"87",
          5759 => x"94",
          5760 => x"71",
          5761 => x"0c",
          5762 => x"04",
          5763 => x"02",
          5764 => x"02",
          5765 => x"05",
          5766 => x"83",
          5767 => x"26",
          5768 => x"72",
          5769 => x"c0",
          5770 => x"53",
          5771 => x"74",
          5772 => x"38",
          5773 => x"73",
          5774 => x"c0",
          5775 => x"51",
          5776 => x"85",
          5777 => x"98",
          5778 => x"52",
          5779 => x"82",
          5780 => x"70",
          5781 => x"38",
          5782 => x"8c",
          5783 => x"ec",
          5784 => x"fc",
          5785 => x"52",
          5786 => x"87",
          5787 => x"08",
          5788 => x"2e",
          5789 => x"82",
          5790 => x"34",
          5791 => x"13",
          5792 => x"82",
          5793 => x"86",
          5794 => x"f3",
          5795 => x"62",
          5796 => x"05",
          5797 => x"57",
          5798 => x"83",
          5799 => x"fe",
          5800 => x"e0",
          5801 => x"06",
          5802 => x"71",
          5803 => x"71",
          5804 => x"2b",
          5805 => x"80",
          5806 => x"92",
          5807 => x"c0",
          5808 => x"41",
          5809 => x"5a",
          5810 => x"87",
          5811 => x"0c",
          5812 => x"84",
          5813 => x"08",
          5814 => x"70",
          5815 => x"53",
          5816 => x"2e",
          5817 => x"08",
          5818 => x"70",
          5819 => x"34",
          5820 => x"80",
          5821 => x"53",
          5822 => x"2e",
          5823 => x"53",
          5824 => x"26",
          5825 => x"80",
          5826 => x"87",
          5827 => x"08",
          5828 => x"38",
          5829 => x"8c",
          5830 => x"80",
          5831 => x"78",
          5832 => x"99",
          5833 => x"0c",
          5834 => x"8c",
          5835 => x"08",
          5836 => x"51",
          5837 => x"38",
          5838 => x"8d",
          5839 => x"17",
          5840 => x"81",
          5841 => x"53",
          5842 => x"2e",
          5843 => x"fc",
          5844 => x"52",
          5845 => x"7d",
          5846 => x"ed",
          5847 => x"80",
          5848 => x"71",
          5849 => x"38",
          5850 => x"53",
          5851 => x"98",
          5852 => x"0d",
          5853 => x"0d",
          5854 => x"02",
          5855 => x"05",
          5856 => x"58",
          5857 => x"80",
          5858 => x"fc",
          5859 => x"e0",
          5860 => x"06",
          5861 => x"71",
          5862 => x"81",
          5863 => x"38",
          5864 => x"2b",
          5865 => x"80",
          5866 => x"92",
          5867 => x"c0",
          5868 => x"40",
          5869 => x"5a",
          5870 => x"c0",
          5871 => x"76",
          5872 => x"76",
          5873 => x"75",
          5874 => x"2a",
          5875 => x"51",
          5876 => x"80",
          5877 => x"7a",
          5878 => x"5c",
          5879 => x"81",
          5880 => x"81",
          5881 => x"06",
          5882 => x"80",
          5883 => x"87",
          5884 => x"08",
          5885 => x"38",
          5886 => x"8c",
          5887 => x"80",
          5888 => x"77",
          5889 => x"99",
          5890 => x"0c",
          5891 => x"8c",
          5892 => x"08",
          5893 => x"51",
          5894 => x"38",
          5895 => x"8d",
          5896 => x"70",
          5897 => x"84",
          5898 => x"5b",
          5899 => x"2e",
          5900 => x"fc",
          5901 => x"52",
          5902 => x"7d",
          5903 => x"f8",
          5904 => x"80",
          5905 => x"71",
          5906 => x"38",
          5907 => x"53",
          5908 => x"98",
          5909 => x"0d",
          5910 => x"0d",
          5911 => x"05",
          5912 => x"02",
          5913 => x"05",
          5914 => x"54",
          5915 => x"fe",
          5916 => x"98",
          5917 => x"53",
          5918 => x"80",
          5919 => x"0b",
          5920 => x"8c",
          5921 => x"71",
          5922 => x"dc",
          5923 => x"24",
          5924 => x"84",
          5925 => x"92",
          5926 => x"54",
          5927 => x"8d",
          5928 => x"39",
          5929 => x"80",
          5930 => x"cb",
          5931 => x"70",
          5932 => x"81",
          5933 => x"52",
          5934 => x"8a",
          5935 => x"98",
          5936 => x"71",
          5937 => x"c0",
          5938 => x"52",
          5939 => x"81",
          5940 => x"c0",
          5941 => x"53",
          5942 => x"82",
          5943 => x"71",
          5944 => x"39",
          5945 => x"39",
          5946 => x"77",
          5947 => x"81",
          5948 => x"72",
          5949 => x"84",
          5950 => x"73",
          5951 => x"0c",
          5952 => x"04",
          5953 => x"74",
          5954 => x"71",
          5955 => x"2b",
          5956 => x"98",
          5957 => x"84",
          5958 => x"fd",
          5959 => x"83",
          5960 => x"12",
          5961 => x"2b",
          5962 => x"07",
          5963 => x"70",
          5964 => x"2b",
          5965 => x"07",
          5966 => x"0c",
          5967 => x"56",
          5968 => x"3d",
          5969 => x"3d",
          5970 => x"84",
          5971 => x"22",
          5972 => x"72",
          5973 => x"54",
          5974 => x"2a",
          5975 => x"34",
          5976 => x"04",
          5977 => x"73",
          5978 => x"70",
          5979 => x"05",
          5980 => x"88",
          5981 => x"72",
          5982 => x"54",
          5983 => x"2a",
          5984 => x"70",
          5985 => x"34",
          5986 => x"51",
          5987 => x"83",
          5988 => x"fe",
          5989 => x"75",
          5990 => x"51",
          5991 => x"92",
          5992 => x"81",
          5993 => x"73",
          5994 => x"55",
          5995 => x"51",
          5996 => x"3d",
          5997 => x"3d",
          5998 => x"76",
          5999 => x"72",
          6000 => x"05",
          6001 => x"11",
          6002 => x"38",
          6003 => x"04",
          6004 => x"78",
          6005 => x"56",
          6006 => x"81",
          6007 => x"74",
          6008 => x"56",
          6009 => x"31",
          6010 => x"52",
          6011 => x"80",
          6012 => x"71",
          6013 => x"38",
          6014 => x"98",
          6015 => x"0d",
          6016 => x"0d",
          6017 => x"51",
          6018 => x"73",
          6019 => x"81",
          6020 => x"33",
          6021 => x"38",
          6022 => x"e0",
          6023 => x"3d",
          6024 => x"0b",
          6025 => x"0c",
          6026 => x"0d",
          6027 => x"70",
          6028 => x"52",
          6029 => x"55",
          6030 => x"3f",
          6031 => x"e0",
          6032 => x"38",
          6033 => x"98",
          6034 => x"52",
          6035 => x"f9",
          6036 => x"e0",
          6037 => x"ff",
          6038 => x"72",
          6039 => x"38",
          6040 => x"72",
          6041 => x"e0",
          6042 => x"3d",
          6043 => x"3d",
          6044 => x"80",
          6045 => x"33",
          6046 => x"7a",
          6047 => x"38",
          6048 => x"16",
          6049 => x"16",
          6050 => x"17",
          6051 => x"f9",
          6052 => x"e0",
          6053 => x"2e",
          6054 => x"b7",
          6055 => x"98",
          6056 => x"34",
          6057 => x"70",
          6058 => x"31",
          6059 => x"59",
          6060 => x"77",
          6061 => x"82",
          6062 => x"74",
          6063 => x"81",
          6064 => x"81",
          6065 => x"53",
          6066 => x"16",
          6067 => x"a5",
          6068 => x"81",
          6069 => x"e0",
          6070 => x"3d",
          6071 => x"3d",
          6072 => x"56",
          6073 => x"74",
          6074 => x"2e",
          6075 => x"51",
          6076 => x"82",
          6077 => x"57",
          6078 => x"08",
          6079 => x"54",
          6080 => x"16",
          6081 => x"33",
          6082 => x"3f",
          6083 => x"08",
          6084 => x"38",
          6085 => x"57",
          6086 => x"0c",
          6087 => x"98",
          6088 => x"0d",
          6089 => x"0d",
          6090 => x"57",
          6091 => x"82",
          6092 => x"58",
          6093 => x"08",
          6094 => x"76",
          6095 => x"83",
          6096 => x"06",
          6097 => x"84",
          6098 => x"78",
          6099 => x"81",
          6100 => x"38",
          6101 => x"82",
          6102 => x"52",
          6103 => x"52",
          6104 => x"3f",
          6105 => x"52",
          6106 => x"51",
          6107 => x"84",
          6108 => x"d2",
          6109 => x"fb",
          6110 => x"8a",
          6111 => x"52",
          6112 => x"51",
          6113 => x"94",
          6114 => x"84",
          6115 => x"fb",
          6116 => x"17",
          6117 => x"a4",
          6118 => x"c8",
          6119 => x"08",
          6120 => x"b4",
          6121 => x"55",
          6122 => x"81",
          6123 => x"f7",
          6124 => x"84",
          6125 => x"53",
          6126 => x"17",
          6127 => x"99",
          6128 => x"98",
          6129 => x"83",
          6130 => x"77",
          6131 => x"0c",
          6132 => x"04",
          6133 => x"77",
          6134 => x"12",
          6135 => x"55",
          6136 => x"56",
          6137 => x"8d",
          6138 => x"22",
          6139 => x"b0",
          6140 => x"57",
          6141 => x"e0",
          6142 => x"3d",
          6143 => x"3d",
          6144 => x"70",
          6145 => x"57",
          6146 => x"81",
          6147 => x"9c",
          6148 => x"81",
          6149 => x"74",
          6150 => x"72",
          6151 => x"f5",
          6152 => x"24",
          6153 => x"81",
          6154 => x"81",
          6155 => x"83",
          6156 => x"38",
          6157 => x"76",
          6158 => x"70",
          6159 => x"16",
          6160 => x"74",
          6161 => x"96",
          6162 => x"98",
          6163 => x"38",
          6164 => x"06",
          6165 => x"33",
          6166 => x"89",
          6167 => x"08",
          6168 => x"54",
          6169 => x"fc",
          6170 => x"e0",
          6171 => x"fe",
          6172 => x"ff",
          6173 => x"11",
          6174 => x"2b",
          6175 => x"81",
          6176 => x"2a",
          6177 => x"51",
          6178 => x"e2",
          6179 => x"ff",
          6180 => x"da",
          6181 => x"2a",
          6182 => x"05",
          6183 => x"fc",
          6184 => x"e0",
          6185 => x"c6",
          6186 => x"83",
          6187 => x"05",
          6188 => x"f8",
          6189 => x"e0",
          6190 => x"ff",
          6191 => x"ae",
          6192 => x"2a",
          6193 => x"05",
          6194 => x"fc",
          6195 => x"e0",
          6196 => x"38",
          6197 => x"83",
          6198 => x"05",
          6199 => x"f8",
          6200 => x"e0",
          6201 => x"0a",
          6202 => x"39",
          6203 => x"82",
          6204 => x"89",
          6205 => x"f8",
          6206 => x"7c",
          6207 => x"56",
          6208 => x"77",
          6209 => x"38",
          6210 => x"08",
          6211 => x"38",
          6212 => x"72",
          6213 => x"9d",
          6214 => x"24",
          6215 => x"81",
          6216 => x"82",
          6217 => x"83",
          6218 => x"38",
          6219 => x"76",
          6220 => x"70",
          6221 => x"18",
          6222 => x"76",
          6223 => x"9e",
          6224 => x"98",
          6225 => x"e0",
          6226 => x"d9",
          6227 => x"ff",
          6228 => x"05",
          6229 => x"81",
          6230 => x"54",
          6231 => x"80",
          6232 => x"77",
          6233 => x"f0",
          6234 => x"8f",
          6235 => x"51",
          6236 => x"34",
          6237 => x"17",
          6238 => x"2a",
          6239 => x"05",
          6240 => x"fa",
          6241 => x"e0",
          6242 => x"82",
          6243 => x"81",
          6244 => x"83",
          6245 => x"b8",
          6246 => x"2a",
          6247 => x"8f",
          6248 => x"2a",
          6249 => x"f0",
          6250 => x"06",
          6251 => x"72",
          6252 => x"ec",
          6253 => x"2a",
          6254 => x"05",
          6255 => x"fa",
          6256 => x"e0",
          6257 => x"82",
          6258 => x"80",
          6259 => x"83",
          6260 => x"52",
          6261 => x"fe",
          6262 => x"b8",
          6263 => x"e6",
          6264 => x"76",
          6265 => x"17",
          6266 => x"75",
          6267 => x"3f",
          6268 => x"08",
          6269 => x"98",
          6270 => x"77",
          6271 => x"77",
          6272 => x"fc",
          6273 => x"b8",
          6274 => x"51",
          6275 => x"8b",
          6276 => x"98",
          6277 => x"06",
          6278 => x"72",
          6279 => x"3f",
          6280 => x"17",
          6281 => x"e0",
          6282 => x"3d",
          6283 => x"3d",
          6284 => x"7e",
          6285 => x"56",
          6286 => x"75",
          6287 => x"74",
          6288 => x"27",
          6289 => x"80",
          6290 => x"ff",
          6291 => x"75",
          6292 => x"3f",
          6293 => x"08",
          6294 => x"98",
          6295 => x"38",
          6296 => x"54",
          6297 => x"81",
          6298 => x"39",
          6299 => x"08",
          6300 => x"39",
          6301 => x"51",
          6302 => x"82",
          6303 => x"58",
          6304 => x"08",
          6305 => x"c7",
          6306 => x"98",
          6307 => x"d2",
          6308 => x"98",
          6309 => x"cf",
          6310 => x"74",
          6311 => x"fc",
          6312 => x"e0",
          6313 => x"38",
          6314 => x"fe",
          6315 => x"08",
          6316 => x"74",
          6317 => x"38",
          6318 => x"17",
          6319 => x"33",
          6320 => x"73",
          6321 => x"77",
          6322 => x"26",
          6323 => x"80",
          6324 => x"e0",
          6325 => x"3d",
          6326 => x"3d",
          6327 => x"71",
          6328 => x"5b",
          6329 => x"90",
          6330 => x"77",
          6331 => x"38",
          6332 => x"78",
          6333 => x"81",
          6334 => x"79",
          6335 => x"f9",
          6336 => x"55",
          6337 => x"98",
          6338 => x"e0",
          6339 => x"98",
          6340 => x"e0",
          6341 => x"2e",
          6342 => x"9c",
          6343 => x"e0",
          6344 => x"82",
          6345 => x"58",
          6346 => x"70",
          6347 => x"80",
          6348 => x"38",
          6349 => x"09",
          6350 => x"e2",
          6351 => x"56",
          6352 => x"76",
          6353 => x"82",
          6354 => x"7a",
          6355 => x"3f",
          6356 => x"e0",
          6357 => x"2e",
          6358 => x"86",
          6359 => x"98",
          6360 => x"e0",
          6361 => x"70",
          6362 => x"07",
          6363 => x"7c",
          6364 => x"98",
          6365 => x"51",
          6366 => x"81",
          6367 => x"e0",
          6368 => x"2e",
          6369 => x"17",
          6370 => x"74",
          6371 => x"73",
          6372 => x"27",
          6373 => x"58",
          6374 => x"80",
          6375 => x"56",
          6376 => x"9c",
          6377 => x"26",
          6378 => x"56",
          6379 => x"81",
          6380 => x"52",
          6381 => x"c6",
          6382 => x"98",
          6383 => x"b8",
          6384 => x"82",
          6385 => x"81",
          6386 => x"06",
          6387 => x"e0",
          6388 => x"82",
          6389 => x"09",
          6390 => x"72",
          6391 => x"70",
          6392 => x"51",
          6393 => x"80",
          6394 => x"78",
          6395 => x"06",
          6396 => x"73",
          6397 => x"39",
          6398 => x"52",
          6399 => x"f7",
          6400 => x"98",
          6401 => x"98",
          6402 => x"82",
          6403 => x"07",
          6404 => x"55",
          6405 => x"2e",
          6406 => x"80",
          6407 => x"75",
          6408 => x"76",
          6409 => x"3f",
          6410 => x"08",
          6411 => x"38",
          6412 => x"0c",
          6413 => x"fe",
          6414 => x"08",
          6415 => x"74",
          6416 => x"ff",
          6417 => x"0c",
          6418 => x"81",
          6419 => x"84",
          6420 => x"39",
          6421 => x"81",
          6422 => x"8c",
          6423 => x"8c",
          6424 => x"98",
          6425 => x"39",
          6426 => x"55",
          6427 => x"98",
          6428 => x"0d",
          6429 => x"0d",
          6430 => x"55",
          6431 => x"82",
          6432 => x"58",
          6433 => x"e0",
          6434 => x"d8",
          6435 => x"74",
          6436 => x"3f",
          6437 => x"08",
          6438 => x"08",
          6439 => x"59",
          6440 => x"77",
          6441 => x"70",
          6442 => x"8a",
          6443 => x"84",
          6444 => x"56",
          6445 => x"58",
          6446 => x"97",
          6447 => x"75",
          6448 => x"52",
          6449 => x"51",
          6450 => x"82",
          6451 => x"80",
          6452 => x"8a",
          6453 => x"32",
          6454 => x"72",
          6455 => x"2a",
          6456 => x"56",
          6457 => x"98",
          6458 => x"0d",
          6459 => x"0d",
          6460 => x"08",
          6461 => x"74",
          6462 => x"26",
          6463 => x"74",
          6464 => x"72",
          6465 => x"74",
          6466 => x"88",
          6467 => x"73",
          6468 => x"33",
          6469 => x"27",
          6470 => x"16",
          6471 => x"9b",
          6472 => x"2a",
          6473 => x"88",
          6474 => x"58",
          6475 => x"80",
          6476 => x"16",
          6477 => x"0c",
          6478 => x"8a",
          6479 => x"89",
          6480 => x"72",
          6481 => x"38",
          6482 => x"51",
          6483 => x"82",
          6484 => x"54",
          6485 => x"08",
          6486 => x"38",
          6487 => x"e0",
          6488 => x"8b",
          6489 => x"08",
          6490 => x"08",
          6491 => x"82",
          6492 => x"74",
          6493 => x"cb",
          6494 => x"75",
          6495 => x"3f",
          6496 => x"08",
          6497 => x"73",
          6498 => x"98",
          6499 => x"82",
          6500 => x"2e",
          6501 => x"39",
          6502 => x"39",
          6503 => x"13",
          6504 => x"74",
          6505 => x"16",
          6506 => x"18",
          6507 => x"77",
          6508 => x"0c",
          6509 => x"04",
          6510 => x"7a",
          6511 => x"12",
          6512 => x"59",
          6513 => x"80",
          6514 => x"86",
          6515 => x"98",
          6516 => x"14",
          6517 => x"55",
          6518 => x"81",
          6519 => x"83",
          6520 => x"77",
          6521 => x"81",
          6522 => x"0c",
          6523 => x"55",
          6524 => x"76",
          6525 => x"17",
          6526 => x"74",
          6527 => x"9b",
          6528 => x"39",
          6529 => x"ff",
          6530 => x"2a",
          6531 => x"81",
          6532 => x"52",
          6533 => x"e6",
          6534 => x"98",
          6535 => x"55",
          6536 => x"e0",
          6537 => x"80",
          6538 => x"55",
          6539 => x"08",
          6540 => x"f4",
          6541 => x"08",
          6542 => x"08",
          6543 => x"38",
          6544 => x"77",
          6545 => x"84",
          6546 => x"39",
          6547 => x"52",
          6548 => x"86",
          6549 => x"98",
          6550 => x"55",
          6551 => x"08",
          6552 => x"c4",
          6553 => x"82",
          6554 => x"81",
          6555 => x"81",
          6556 => x"98",
          6557 => x"b0",
          6558 => x"98",
          6559 => x"51",
          6560 => x"82",
          6561 => x"a0",
          6562 => x"15",
          6563 => x"75",
          6564 => x"3f",
          6565 => x"08",
          6566 => x"76",
          6567 => x"77",
          6568 => x"9c",
          6569 => x"55",
          6570 => x"98",
          6571 => x"0d",
          6572 => x"0d",
          6573 => x"08",
          6574 => x"80",
          6575 => x"fc",
          6576 => x"e0",
          6577 => x"82",
          6578 => x"80",
          6579 => x"e0",
          6580 => x"98",
          6581 => x"78",
          6582 => x"3f",
          6583 => x"08",
          6584 => x"98",
          6585 => x"38",
          6586 => x"08",
          6587 => x"70",
          6588 => x"58",
          6589 => x"2e",
          6590 => x"83",
          6591 => x"82",
          6592 => x"55",
          6593 => x"81",
          6594 => x"07",
          6595 => x"2e",
          6596 => x"16",
          6597 => x"2e",
          6598 => x"88",
          6599 => x"82",
          6600 => x"56",
          6601 => x"51",
          6602 => x"82",
          6603 => x"54",
          6604 => x"08",
          6605 => x"9b",
          6606 => x"2e",
          6607 => x"83",
          6608 => x"73",
          6609 => x"0c",
          6610 => x"04",
          6611 => x"76",
          6612 => x"54",
          6613 => x"82",
          6614 => x"83",
          6615 => x"76",
          6616 => x"53",
          6617 => x"2e",
          6618 => x"90",
          6619 => x"51",
          6620 => x"82",
          6621 => x"90",
          6622 => x"53",
          6623 => x"98",
          6624 => x"0d",
          6625 => x"0d",
          6626 => x"83",
          6627 => x"54",
          6628 => x"55",
          6629 => x"3f",
          6630 => x"51",
          6631 => x"2e",
          6632 => x"8b",
          6633 => x"2a",
          6634 => x"51",
          6635 => x"86",
          6636 => x"fd",
          6637 => x"54",
          6638 => x"53",
          6639 => x"71",
          6640 => x"05",
          6641 => x"05",
          6642 => x"05",
          6643 => x"06",
          6644 => x"51",
          6645 => x"e4",
          6646 => x"e0",
          6647 => x"3d",
          6648 => x"3d",
          6649 => x"40",
          6650 => x"08",
          6651 => x"ff",
          6652 => x"98",
          6653 => x"2e",
          6654 => x"98",
          6655 => x"7d",
          6656 => x"3f",
          6657 => x"08",
          6658 => x"98",
          6659 => x"38",
          6660 => x"70",
          6661 => x"73",
          6662 => x"5b",
          6663 => x"8b",
          6664 => x"06",
          6665 => x"06",
          6666 => x"86",
          6667 => x"e0",
          6668 => x"73",
          6669 => x"09",
          6670 => x"38",
          6671 => x"e0",
          6672 => x"73",
          6673 => x"81",
          6674 => x"81",
          6675 => x"07",
          6676 => x"38",
          6677 => x"08",
          6678 => x"54",
          6679 => x"2e",
          6680 => x"83",
          6681 => x"75",
          6682 => x"38",
          6683 => x"81",
          6684 => x"8f",
          6685 => x"06",
          6686 => x"73",
          6687 => x"81",
          6688 => x"72",
          6689 => x"38",
          6690 => x"74",
          6691 => x"70",
          6692 => x"ac",
          6693 => x"5d",
          6694 => x"2e",
          6695 => x"81",
          6696 => x"15",
          6697 => x"73",
          6698 => x"06",
          6699 => x"8c",
          6700 => x"16",
          6701 => x"cc",
          6702 => x"98",
          6703 => x"ff",
          6704 => x"80",
          6705 => x"33",
          6706 => x"06",
          6707 => x"05",
          6708 => x"7b",
          6709 => x"d2",
          6710 => x"75",
          6711 => x"a4",
          6712 => x"98",
          6713 => x"ff",
          6714 => x"80",
          6715 => x"73",
          6716 => x"80",
          6717 => x"10",
          6718 => x"53",
          6719 => x"81",
          6720 => x"39",
          6721 => x"ff",
          6722 => x"06",
          6723 => x"17",
          6724 => x"27",
          6725 => x"33",
          6726 => x"70",
          6727 => x"54",
          6728 => x"2e",
          6729 => x"81",
          6730 => x"38",
          6731 => x"53",
          6732 => x"ff",
          6733 => x"ff",
          6734 => x"84",
          6735 => x"53",
          6736 => x"39",
          6737 => x"74",
          6738 => x"3f",
          6739 => x"08",
          6740 => x"53",
          6741 => x"a7",
          6742 => x"ac",
          6743 => x"39",
          6744 => x"51",
          6745 => x"82",
          6746 => x"5b",
          6747 => x"08",
          6748 => x"19",
          6749 => x"38",
          6750 => x"0b",
          6751 => x"7a",
          6752 => x"0c",
          6753 => x"04",
          6754 => x"60",
          6755 => x"59",
          6756 => x"51",
          6757 => x"82",
          6758 => x"58",
          6759 => x"08",
          6760 => x"81",
          6761 => x"5c",
          6762 => x"1a",
          6763 => x"08",
          6764 => x"ea",
          6765 => x"e0",
          6766 => x"82",
          6767 => x"83",
          6768 => x"19",
          6769 => x"57",
          6770 => x"38",
          6771 => x"f6",
          6772 => x"33",
          6773 => x"81",
          6774 => x"54",
          6775 => x"34",
          6776 => x"2e",
          6777 => x"74",
          6778 => x"81",
          6779 => x"74",
          6780 => x"38",
          6781 => x"38",
          6782 => x"09",
          6783 => x"f7",
          6784 => x"33",
          6785 => x"70",
          6786 => x"55",
          6787 => x"a1",
          6788 => x"2a",
          6789 => x"51",
          6790 => x"2e",
          6791 => x"17",
          6792 => x"bf",
          6793 => x"1c",
          6794 => x"0c",
          6795 => x"75",
          6796 => x"81",
          6797 => x"38",
          6798 => x"56",
          6799 => x"09",
          6800 => x"ac",
          6801 => x"08",
          6802 => x"5d",
          6803 => x"82",
          6804 => x"83",
          6805 => x"55",
          6806 => x"38",
          6807 => x"bf",
          6808 => x"f3",
          6809 => x"81",
          6810 => x"82",
          6811 => x"33",
          6812 => x"e5",
          6813 => x"e0",
          6814 => x"ff",
          6815 => x"79",
          6816 => x"38",
          6817 => x"26",
          6818 => x"75",
          6819 => x"a0",
          6820 => x"98",
          6821 => x"1e",
          6822 => x"55",
          6823 => x"55",
          6824 => x"3f",
          6825 => x"98",
          6826 => x"81",
          6827 => x"38",
          6828 => x"39",
          6829 => x"ff",
          6830 => x"06",
          6831 => x"1b",
          6832 => x"27",
          6833 => x"76",
          6834 => x"2a",
          6835 => x"51",
          6836 => x"80",
          6837 => x"73",
          6838 => x"38",
          6839 => x"70",
          6840 => x"73",
          6841 => x"1c",
          6842 => x"06",
          6843 => x"39",
          6844 => x"73",
          6845 => x"7b",
          6846 => x"51",
          6847 => x"82",
          6848 => x"81",
          6849 => x"73",
          6850 => x"38",
          6851 => x"81",
          6852 => x"95",
          6853 => x"a0",
          6854 => x"19",
          6855 => x"b0",
          6856 => x"98",
          6857 => x"9e",
          6858 => x"5c",
          6859 => x"1a",
          6860 => x"78",
          6861 => x"3f",
          6862 => x"08",
          6863 => x"98",
          6864 => x"fc",
          6865 => x"82",
          6866 => x"90",
          6867 => x"ee",
          6868 => x"70",
          6869 => x"33",
          6870 => x"56",
          6871 => x"55",
          6872 => x"38",
          6873 => x"08",
          6874 => x"56",
          6875 => x"2e",
          6876 => x"1d",
          6877 => x"70",
          6878 => x"5d",
          6879 => x"53",
          6880 => x"53",
          6881 => x"53",
          6882 => x"87",
          6883 => x"cb",
          6884 => x"06",
          6885 => x"2e",
          6886 => x"80",
          6887 => x"1b",
          6888 => x"8c",
          6889 => x"56",
          6890 => x"7d",
          6891 => x"e3",
          6892 => x"7b",
          6893 => x"38",
          6894 => x"22",
          6895 => x"ff",
          6896 => x"73",
          6897 => x"38",
          6898 => x"ff",
          6899 => x"59",
          6900 => x"74",
          6901 => x"10",
          6902 => x"2a",
          6903 => x"70",
          6904 => x"56",
          6905 => x"80",
          6906 => x"75",
          6907 => x"32",
          6908 => x"57",
          6909 => x"db",
          6910 => x"75",
          6911 => x"84",
          6912 => x"57",
          6913 => x"07",
          6914 => x"b9",
          6915 => x"38",
          6916 => x"73",
          6917 => x"16",
          6918 => x"84",
          6919 => x"56",
          6920 => x"94",
          6921 => x"17",
          6922 => x"74",
          6923 => x"27",
          6924 => x"33",
          6925 => x"2e",
          6926 => x"19",
          6927 => x"54",
          6928 => x"82",
          6929 => x"80",
          6930 => x"ff",
          6931 => x"74",
          6932 => x"81",
          6933 => x"15",
          6934 => x"27",
          6935 => x"19",
          6936 => x"54",
          6937 => x"3d",
          6938 => x"05",
          6939 => x"81",
          6940 => x"a0",
          6941 => x"26",
          6942 => x"17",
          6943 => x"33",
          6944 => x"75",
          6945 => x"75",
          6946 => x"79",
          6947 => x"3f",
          6948 => x"08",
          6949 => x"1b",
          6950 => x"7b",
          6951 => x"38",
          6952 => x"80",
          6953 => x"f0",
          6954 => x"98",
          6955 => x"e0",
          6956 => x"2e",
          6957 => x"82",
          6958 => x"80",
          6959 => x"ab",
          6960 => x"80",
          6961 => x"70",
          6962 => x"81",
          6963 => x"5e",
          6964 => x"80",
          6965 => x"8d",
          6966 => x"51",
          6967 => x"3f",
          6968 => x"08",
          6969 => x"52",
          6970 => x"c5",
          6971 => x"98",
          6972 => x"e0",
          6973 => x"9e",
          6974 => x"59",
          6975 => x"81",
          6976 => x"85",
          6977 => x"08",
          6978 => x"54",
          6979 => x"dd",
          6980 => x"98",
          6981 => x"e0",
          6982 => x"fa",
          6983 => x"51",
          6984 => x"82",
          6985 => x"81",
          6986 => x"98",
          6987 => x"7b",
          6988 => x"3f",
          6989 => x"08",
          6990 => x"98",
          6991 => x"38",
          6992 => x"9c",
          6993 => x"81",
          6994 => x"57",
          6995 => x"17",
          6996 => x"8b",
          6997 => x"e0",
          6998 => x"17",
          6999 => x"98",
          7000 => x"16",
          7001 => x"3f",
          7002 => x"f3",
          7003 => x"55",
          7004 => x"ff",
          7005 => x"74",
          7006 => x"22",
          7007 => x"51",
          7008 => x"82",
          7009 => x"33",
          7010 => x"df",
          7011 => x"85",
          7012 => x"ff",
          7013 => x"57",
          7014 => x"d4",
          7015 => x"ff",
          7016 => x"38",
          7017 => x"70",
          7018 => x"73",
          7019 => x"80",
          7020 => x"77",
          7021 => x"0b",
          7022 => x"80",
          7023 => x"ef",
          7024 => x"e0",
          7025 => x"82",
          7026 => x"80",
          7027 => x"19",
          7028 => x"d7",
          7029 => x"08",
          7030 => x"e2",
          7031 => x"e0",
          7032 => x"82",
          7033 => x"ae",
          7034 => x"82",
          7035 => x"52",
          7036 => x"51",
          7037 => x"8b",
          7038 => x"52",
          7039 => x"51",
          7040 => x"9c",
          7041 => x"1b",
          7042 => x"55",
          7043 => x"16",
          7044 => x"83",
          7045 => x"55",
          7046 => x"98",
          7047 => x"0d",
          7048 => x"0d",
          7049 => x"90",
          7050 => x"13",
          7051 => x"57",
          7052 => x"2e",
          7053 => x"52",
          7054 => x"b1",
          7055 => x"98",
          7056 => x"e0",
          7057 => x"c9",
          7058 => x"08",
          7059 => x"e1",
          7060 => x"e0",
          7061 => x"82",
          7062 => x"ab",
          7063 => x"08",
          7064 => x"34",
          7065 => x"17",
          7066 => x"08",
          7067 => x"38",
          7068 => x"08",
          7069 => x"ee",
          7070 => x"e0",
          7071 => x"82",
          7072 => x"80",
          7073 => x"73",
          7074 => x"81",
          7075 => x"82",
          7076 => x"e0",
          7077 => x"3d",
          7078 => x"3d",
          7079 => x"71",
          7080 => x"5c",
          7081 => x"19",
          7082 => x"08",
          7083 => x"e2",
          7084 => x"08",
          7085 => x"bb",
          7086 => x"71",
          7087 => x"08",
          7088 => x"57",
          7089 => x"72",
          7090 => x"9d",
          7091 => x"14",
          7092 => x"1b",
          7093 => x"7a",
          7094 => x"d0",
          7095 => x"83",
          7096 => x"51",
          7097 => x"ff",
          7098 => x"74",
          7099 => x"39",
          7100 => x"11",
          7101 => x"31",
          7102 => x"83",
          7103 => x"90",
          7104 => x"51",
          7105 => x"3f",
          7106 => x"08",
          7107 => x"06",
          7108 => x"75",
          7109 => x"81",
          7110 => x"38",
          7111 => x"53",
          7112 => x"74",
          7113 => x"82",
          7114 => x"74",
          7115 => x"70",
          7116 => x"25",
          7117 => x"07",
          7118 => x"73",
          7119 => x"38",
          7120 => x"39",
          7121 => x"81",
          7122 => x"57",
          7123 => x"1d",
          7124 => x"11",
          7125 => x"54",
          7126 => x"f1",
          7127 => x"70",
          7128 => x"30",
          7129 => x"51",
          7130 => x"94",
          7131 => x"0b",
          7132 => x"80",
          7133 => x"58",
          7134 => x"1c",
          7135 => x"33",
          7136 => x"56",
          7137 => x"2e",
          7138 => x"85",
          7139 => x"06",
          7140 => x"e5",
          7141 => x"32",
          7142 => x"72",
          7143 => x"51",
          7144 => x"8b",
          7145 => x"72",
          7146 => x"38",
          7147 => x"81",
          7148 => x"81",
          7149 => x"76",
          7150 => x"58",
          7151 => x"57",
          7152 => x"ff",
          7153 => x"17",
          7154 => x"80",
          7155 => x"34",
          7156 => x"53",
          7157 => x"38",
          7158 => x"bf",
          7159 => x"34",
          7160 => x"e1",
          7161 => x"89",
          7162 => x"5a",
          7163 => x"2e",
          7164 => x"96",
          7165 => x"55",
          7166 => x"ff",
          7167 => x"55",
          7168 => x"aa",
          7169 => x"08",
          7170 => x"51",
          7171 => x"27",
          7172 => x"84",
          7173 => x"39",
          7174 => x"53",
          7175 => x"53",
          7176 => x"8a",
          7177 => x"70",
          7178 => x"06",
          7179 => x"76",
          7180 => x"58",
          7181 => x"81",
          7182 => x"71",
          7183 => x"55",
          7184 => x"b5",
          7185 => x"94",
          7186 => x"0b",
          7187 => x"9c",
          7188 => x"11",
          7189 => x"72",
          7190 => x"89",
          7191 => x"1c",
          7192 => x"13",
          7193 => x"34",
          7194 => x"9c",
          7195 => x"d9",
          7196 => x"e0",
          7197 => x"0c",
          7198 => x"d9",
          7199 => x"e0",
          7200 => x"19",
          7201 => x"51",
          7202 => x"82",
          7203 => x"84",
          7204 => x"3d",
          7205 => x"3d",
          7206 => x"08",
          7207 => x"64",
          7208 => x"55",
          7209 => x"2e",
          7210 => x"55",
          7211 => x"2e",
          7212 => x"80",
          7213 => x"7f",
          7214 => x"88",
          7215 => x"39",
          7216 => x"80",
          7217 => x"56",
          7218 => x"af",
          7219 => x"06",
          7220 => x"56",
          7221 => x"32",
          7222 => x"80",
          7223 => x"51",
          7224 => x"dc",
          7225 => x"1f",
          7226 => x"33",
          7227 => x"9f",
          7228 => x"ff",
          7229 => x"1f",
          7230 => x"7d",
          7231 => x"3f",
          7232 => x"08",
          7233 => x"39",
          7234 => x"08",
          7235 => x"5b",
          7236 => x"92",
          7237 => x"51",
          7238 => x"82",
          7239 => x"ff",
          7240 => x"38",
          7241 => x"0b",
          7242 => x"08",
          7243 => x"78",
          7244 => x"e0",
          7245 => x"2a",
          7246 => x"75",
          7247 => x"59",
          7248 => x"08",
          7249 => x"06",
          7250 => x"70",
          7251 => x"27",
          7252 => x"07",
          7253 => x"56",
          7254 => x"75",
          7255 => x"ae",
          7256 => x"ff",
          7257 => x"75",
          7258 => x"c4",
          7259 => x"3f",
          7260 => x"08",
          7261 => x"78",
          7262 => x"81",
          7263 => x"10",
          7264 => x"74",
          7265 => x"59",
          7266 => x"81",
          7267 => x"61",
          7268 => x"56",
          7269 => x"2e",
          7270 => x"83",
          7271 => x"73",
          7272 => x"70",
          7273 => x"25",
          7274 => x"51",
          7275 => x"38",
          7276 => x"76",
          7277 => x"57",
          7278 => x"09",
          7279 => x"38",
          7280 => x"73",
          7281 => x"38",
          7282 => x"78",
          7283 => x"81",
          7284 => x"38",
          7285 => x"54",
          7286 => x"09",
          7287 => x"c1",
          7288 => x"54",
          7289 => x"09",
          7290 => x"38",
          7291 => x"54",
          7292 => x"80",
          7293 => x"56",
          7294 => x"78",
          7295 => x"38",
          7296 => x"75",
          7297 => x"57",
          7298 => x"58",
          7299 => x"e9",
          7300 => x"07",
          7301 => x"1f",
          7302 => x"39",
          7303 => x"a8",
          7304 => x"1a",
          7305 => x"74",
          7306 => x"71",
          7307 => x"70",
          7308 => x"2a",
          7309 => x"58",
          7310 => x"ae",
          7311 => x"73",
          7312 => x"19",
          7313 => x"38",
          7314 => x"11",
          7315 => x"74",
          7316 => x"38",
          7317 => x"90",
          7318 => x"07",
          7319 => x"39",
          7320 => x"70",
          7321 => x"06",
          7322 => x"73",
          7323 => x"81",
          7324 => x"81",
          7325 => x"1b",
          7326 => x"55",
          7327 => x"2e",
          7328 => x"8f",
          7329 => x"ff",
          7330 => x"73",
          7331 => x"81",
          7332 => x"76",
          7333 => x"78",
          7334 => x"38",
          7335 => x"05",
          7336 => x"54",
          7337 => x"9d",
          7338 => x"1a",
          7339 => x"ff",
          7340 => x"80",
          7341 => x"fe",
          7342 => x"55",
          7343 => x"2e",
          7344 => x"eb",
          7345 => x"a0",
          7346 => x"51",
          7347 => x"80",
          7348 => x"88",
          7349 => x"1a",
          7350 => x"1f",
          7351 => x"75",
          7352 => x"94",
          7353 => x"2e",
          7354 => x"ae",
          7355 => x"70",
          7356 => x"51",
          7357 => x"2e",
          7358 => x"80",
          7359 => x"76",
          7360 => x"d1",
          7361 => x"73",
          7362 => x"26",
          7363 => x"5b",
          7364 => x"70",
          7365 => x"07",
          7366 => x"7e",
          7367 => x"55",
          7368 => x"2e",
          7369 => x"8b",
          7370 => x"38",
          7371 => x"8b",
          7372 => x"07",
          7373 => x"26",
          7374 => x"78",
          7375 => x"8b",
          7376 => x"81",
          7377 => x"5f",
          7378 => x"80",
          7379 => x"af",
          7380 => x"07",
          7381 => x"52",
          7382 => x"ce",
          7383 => x"e0",
          7384 => x"ff",
          7385 => x"87",
          7386 => x"06",
          7387 => x"73",
          7388 => x"38",
          7389 => x"06",
          7390 => x"11",
          7391 => x"81",
          7392 => x"a4",
          7393 => x"54",
          7394 => x"8a",
          7395 => x"07",
          7396 => x"fe",
          7397 => x"18",
          7398 => x"88",
          7399 => x"73",
          7400 => x"18",
          7401 => x"39",
          7402 => x"92",
          7403 => x"82",
          7404 => x"d4",
          7405 => x"e0",
          7406 => x"2e",
          7407 => x"df",
          7408 => x"58",
          7409 => x"ff",
          7410 => x"73",
          7411 => x"38",
          7412 => x"5c",
          7413 => x"54",
          7414 => x"8e",
          7415 => x"07",
          7416 => x"83",
          7417 => x"58",
          7418 => x"18",
          7419 => x"75",
          7420 => x"18",
          7421 => x"39",
          7422 => x"54",
          7423 => x"2e",
          7424 => x"86",
          7425 => x"a0",
          7426 => x"88",
          7427 => x"06",
          7428 => x"82",
          7429 => x"06",
          7430 => x"06",
          7431 => x"2e",
          7432 => x"83",
          7433 => x"83",
          7434 => x"06",
          7435 => x"82",
          7436 => x"81",
          7437 => x"06",
          7438 => x"9f",
          7439 => x"06",
          7440 => x"2e",
          7441 => x"90",
          7442 => x"82",
          7443 => x"06",
          7444 => x"80",
          7445 => x"76",
          7446 => x"76",
          7447 => x"7d",
          7448 => x"3f",
          7449 => x"08",
          7450 => x"56",
          7451 => x"98",
          7452 => x"be",
          7453 => x"98",
          7454 => x"09",
          7455 => x"e8",
          7456 => x"2a",
          7457 => x"76",
          7458 => x"51",
          7459 => x"2e",
          7460 => x"81",
          7461 => x"80",
          7462 => x"38",
          7463 => x"ab",
          7464 => x"56",
          7465 => x"74",
          7466 => x"73",
          7467 => x"56",
          7468 => x"82",
          7469 => x"06",
          7470 => x"ac",
          7471 => x"33",
          7472 => x"70",
          7473 => x"55",
          7474 => x"2e",
          7475 => x"1e",
          7476 => x"06",
          7477 => x"05",
          7478 => x"e4",
          7479 => x"e0",
          7480 => x"1f",
          7481 => x"39",
          7482 => x"98",
          7483 => x"0d",
          7484 => x"0d",
          7485 => x"7b",
          7486 => x"73",
          7487 => x"55",
          7488 => x"2e",
          7489 => x"75",
          7490 => x"57",
          7491 => x"26",
          7492 => x"ba",
          7493 => x"70",
          7494 => x"ba",
          7495 => x"06",
          7496 => x"73",
          7497 => x"70",
          7498 => x"51",
          7499 => x"89",
          7500 => x"82",
          7501 => x"ff",
          7502 => x"56",
          7503 => x"2e",
          7504 => x"80",
          7505 => x"98",
          7506 => x"08",
          7507 => x"76",
          7508 => x"58",
          7509 => x"81",
          7510 => x"ff",
          7511 => x"53",
          7512 => x"26",
          7513 => x"13",
          7514 => x"06",
          7515 => x"9f",
          7516 => x"99",
          7517 => x"e0",
          7518 => x"ff",
          7519 => x"72",
          7520 => x"2a",
          7521 => x"72",
          7522 => x"06",
          7523 => x"ff",
          7524 => x"30",
          7525 => x"70",
          7526 => x"07",
          7527 => x"9f",
          7528 => x"54",
          7529 => x"80",
          7530 => x"81",
          7531 => x"59",
          7532 => x"25",
          7533 => x"8b",
          7534 => x"24",
          7535 => x"76",
          7536 => x"78",
          7537 => x"82",
          7538 => x"51",
          7539 => x"98",
          7540 => x"0d",
          7541 => x"0d",
          7542 => x"0b",
          7543 => x"ff",
          7544 => x"0c",
          7545 => x"51",
          7546 => x"84",
          7547 => x"98",
          7548 => x"38",
          7549 => x"51",
          7550 => x"82",
          7551 => x"83",
          7552 => x"54",
          7553 => x"82",
          7554 => x"09",
          7555 => x"e3",
          7556 => x"b8",
          7557 => x"57",
          7558 => x"2e",
          7559 => x"83",
          7560 => x"74",
          7561 => x"70",
          7562 => x"25",
          7563 => x"51",
          7564 => x"38",
          7565 => x"2e",
          7566 => x"b5",
          7567 => x"82",
          7568 => x"80",
          7569 => x"cf",
          7570 => x"e0",
          7571 => x"82",
          7572 => x"80",
          7573 => x"85",
          7574 => x"dc",
          7575 => x"16",
          7576 => x"3f",
          7577 => x"08",
          7578 => x"98",
          7579 => x"83",
          7580 => x"74",
          7581 => x"0c",
          7582 => x"04",
          7583 => x"61",
          7584 => x"80",
          7585 => x"58",
          7586 => x"0c",
          7587 => x"e1",
          7588 => x"98",
          7589 => x"56",
          7590 => x"e0",
          7591 => x"87",
          7592 => x"e0",
          7593 => x"29",
          7594 => x"05",
          7595 => x"53",
          7596 => x"80",
          7597 => x"38",
          7598 => x"76",
          7599 => x"74",
          7600 => x"72",
          7601 => x"38",
          7602 => x"51",
          7603 => x"82",
          7604 => x"81",
          7605 => x"81",
          7606 => x"72",
          7607 => x"80",
          7608 => x"38",
          7609 => x"70",
          7610 => x"53",
          7611 => x"86",
          7612 => x"f2",
          7613 => x"34",
          7614 => x"82",
          7615 => x"33",
          7616 => x"81",
          7617 => x"33",
          7618 => x"3f",
          7619 => x"08",
          7620 => x"70",
          7621 => x"55",
          7622 => x"86",
          7623 => x"80",
          7624 => x"74",
          7625 => x"81",
          7626 => x"8a",
          7627 => x"b8",
          7628 => x"53",
          7629 => x"fd",
          7630 => x"e0",
          7631 => x"ff",
          7632 => x"82",
          7633 => x"76",
          7634 => x"9c",
          7635 => x"8d",
          7636 => x"72",
          7637 => x"90",
          7638 => x"74",
          7639 => x"56",
          7640 => x"33",
          7641 => x"72",
          7642 => x"38",
          7643 => x"51",
          7644 => x"82",
          7645 => x"57",
          7646 => x"84",
          7647 => x"ff",
          7648 => x"56",
          7649 => x"25",
          7650 => x"18",
          7651 => x"11",
          7652 => x"70",
          7653 => x"71",
          7654 => x"71",
          7655 => x"f0",
          7656 => x"51",
          7657 => x"74",
          7658 => x"57",
          7659 => x"90",
          7660 => x"73",
          7661 => x"3f",
          7662 => x"08",
          7663 => x"57",
          7664 => x"e0",
          7665 => x"54",
          7666 => x"2e",
          7667 => x"83",
          7668 => x"81",
          7669 => x"38",
          7670 => x"8c",
          7671 => x"84",
          7672 => x"83",
          7673 => x"38",
          7674 => x"84",
          7675 => x"38",
          7676 => x"81",
          7677 => x"38",
          7678 => x"51",
          7679 => x"82",
          7680 => x"83",
          7681 => x"53",
          7682 => x"2e",
          7683 => x"84",
          7684 => x"ce",
          7685 => x"ec",
          7686 => x"98",
          7687 => x"ff",
          7688 => x"8d",
          7689 => x"14",
          7690 => x"3f",
          7691 => x"08",
          7692 => x"15",
          7693 => x"14",
          7694 => x"34",
          7695 => x"33",
          7696 => x"81",
          7697 => x"54",
          7698 => x"72",
          7699 => x"98",
          7700 => x"ff",
          7701 => x"29",
          7702 => x"33",
          7703 => x"72",
          7704 => x"72",
          7705 => x"38",
          7706 => x"06",
          7707 => x"2e",
          7708 => x"56",
          7709 => x"80",
          7710 => x"c9",
          7711 => x"e0",
          7712 => x"82",
          7713 => x"88",
          7714 => x"8f",
          7715 => x"56",
          7716 => x"38",
          7717 => x"51",
          7718 => x"82",
          7719 => x"83",
          7720 => x"55",
          7721 => x"80",
          7722 => x"c8",
          7723 => x"e0",
          7724 => x"80",
          7725 => x"c8",
          7726 => x"e0",
          7727 => x"ff",
          7728 => x"8d",
          7729 => x"2e",
          7730 => x"88",
          7731 => x"14",
          7732 => x"05",
          7733 => x"75",
          7734 => x"38",
          7735 => x"52",
          7736 => x"51",
          7737 => x"3f",
          7738 => x"08",
          7739 => x"98",
          7740 => x"82",
          7741 => x"e0",
          7742 => x"ff",
          7743 => x"26",
          7744 => x"57",
          7745 => x"f5",
          7746 => x"82",
          7747 => x"f5",
          7748 => x"81",
          7749 => x"8d",
          7750 => x"2e",
          7751 => x"82",
          7752 => x"16",
          7753 => x"16",
          7754 => x"70",
          7755 => x"7a",
          7756 => x"0c",
          7757 => x"83",
          7758 => x"06",
          7759 => x"e2",
          7760 => x"c0",
          7761 => x"98",
          7762 => x"ff",
          7763 => x"56",
          7764 => x"38",
          7765 => x"38",
          7766 => x"51",
          7767 => x"82",
          7768 => x"ac",
          7769 => x"82",
          7770 => x"39",
          7771 => x"80",
          7772 => x"38",
          7773 => x"15",
          7774 => x"53",
          7775 => x"8d",
          7776 => x"15",
          7777 => x"76",
          7778 => x"51",
          7779 => x"13",
          7780 => x"8d",
          7781 => x"15",
          7782 => x"cc",
          7783 => x"94",
          7784 => x"0b",
          7785 => x"ff",
          7786 => x"15",
          7787 => x"2e",
          7788 => x"81",
          7789 => x"e8",
          7790 => x"c8",
          7791 => x"98",
          7792 => x"ff",
          7793 => x"81",
          7794 => x"06",
          7795 => x"81",
          7796 => x"51",
          7797 => x"82",
          7798 => x"80",
          7799 => x"e0",
          7800 => x"15",
          7801 => x"14",
          7802 => x"3f",
          7803 => x"08",
          7804 => x"06",
          7805 => x"d4",
          7806 => x"81",
          7807 => x"38",
          7808 => x"c6",
          7809 => x"e0",
          7810 => x"8b",
          7811 => x"2e",
          7812 => x"b3",
          7813 => x"14",
          7814 => x"3f",
          7815 => x"08",
          7816 => x"e4",
          7817 => x"81",
          7818 => x"84",
          7819 => x"c5",
          7820 => x"e0",
          7821 => x"15",
          7822 => x"14",
          7823 => x"3f",
          7824 => x"08",
          7825 => x"76",
          7826 => x"f7",
          7827 => x"05",
          7828 => x"f7",
          7829 => x"86",
          7830 => x"f7",
          7831 => x"15",
          7832 => x"98",
          7833 => x"56",
          7834 => x"98",
          7835 => x"0d",
          7836 => x"0d",
          7837 => x"55",
          7838 => x"ba",
          7839 => x"53",
          7840 => x"b2",
          7841 => x"52",
          7842 => x"aa",
          7843 => x"22",
          7844 => x"57",
          7845 => x"2e",
          7846 => x"9a",
          7847 => x"33",
          7848 => x"ca",
          7849 => x"98",
          7850 => x"52",
          7851 => x"71",
          7852 => x"55",
          7853 => x"53",
          7854 => x"0c",
          7855 => x"e0",
          7856 => x"3d",
          7857 => x"3d",
          7858 => x"05",
          7859 => x"89",
          7860 => x"52",
          7861 => x"3f",
          7862 => x"0b",
          7863 => x"08",
          7864 => x"82",
          7865 => x"84",
          7866 => x"e0",
          7867 => x"55",
          7868 => x"2e",
          7869 => x"74",
          7870 => x"73",
          7871 => x"38",
          7872 => x"78",
          7873 => x"54",
          7874 => x"92",
          7875 => x"89",
          7876 => x"84",
          7877 => x"e4",
          7878 => x"98",
          7879 => x"82",
          7880 => x"88",
          7881 => x"ea",
          7882 => x"02",
          7883 => x"eb",
          7884 => x"59",
          7885 => x"80",
          7886 => x"38",
          7887 => x"70",
          7888 => x"cc",
          7889 => x"3d",
          7890 => x"58",
          7891 => x"82",
          7892 => x"55",
          7893 => x"08",
          7894 => x"7a",
          7895 => x"8c",
          7896 => x"56",
          7897 => x"82",
          7898 => x"55",
          7899 => x"08",
          7900 => x"80",
          7901 => x"70",
          7902 => x"57",
          7903 => x"83",
          7904 => x"77",
          7905 => x"73",
          7906 => x"ab",
          7907 => x"2e",
          7908 => x"84",
          7909 => x"06",
          7910 => x"51",
          7911 => x"82",
          7912 => x"55",
          7913 => x"b2",
          7914 => x"06",
          7915 => x"b8",
          7916 => x"2a",
          7917 => x"51",
          7918 => x"2e",
          7919 => x"55",
          7920 => x"77",
          7921 => x"74",
          7922 => x"77",
          7923 => x"81",
          7924 => x"73",
          7925 => x"af",
          7926 => x"7a",
          7927 => x"3f",
          7928 => x"08",
          7929 => x"b2",
          7930 => x"8e",
          7931 => x"f4",
          7932 => x"a0",
          7933 => x"34",
          7934 => x"52",
          7935 => x"85",
          7936 => x"62",
          7937 => x"c2",
          7938 => x"54",
          7939 => x"15",
          7940 => x"2e",
          7941 => x"7a",
          7942 => x"51",
          7943 => x"75",
          7944 => x"d0",
          7945 => x"86",
          7946 => x"98",
          7947 => x"e0",
          7948 => x"ca",
          7949 => x"74",
          7950 => x"02",
          7951 => x"70",
          7952 => x"81",
          7953 => x"56",
          7954 => x"86",
          7955 => x"82",
          7956 => x"81",
          7957 => x"06",
          7958 => x"80",
          7959 => x"75",
          7960 => x"73",
          7961 => x"38",
          7962 => x"92",
          7963 => x"7a",
          7964 => x"3f",
          7965 => x"08",
          7966 => x"90",
          7967 => x"55",
          7968 => x"08",
          7969 => x"77",
          7970 => x"81",
          7971 => x"73",
          7972 => x"38",
          7973 => x"07",
          7974 => x"11",
          7975 => x"0c",
          7976 => x"0c",
          7977 => x"52",
          7978 => x"3f",
          7979 => x"08",
          7980 => x"08",
          7981 => x"63",
          7982 => x"5a",
          7983 => x"82",
          7984 => x"82",
          7985 => x"8c",
          7986 => x"7a",
          7987 => x"17",
          7988 => x"23",
          7989 => x"34",
          7990 => x"1a",
          7991 => x"9c",
          7992 => x"0b",
          7993 => x"77",
          7994 => x"81",
          7995 => x"73",
          7996 => x"8d",
          7997 => x"98",
          7998 => x"81",
          7999 => x"e0",
          8000 => x"1a",
          8001 => x"22",
          8002 => x"7b",
          8003 => x"a8",
          8004 => x"78",
          8005 => x"3f",
          8006 => x"08",
          8007 => x"98",
          8008 => x"83",
          8009 => x"82",
          8010 => x"ff",
          8011 => x"06",
          8012 => x"55",
          8013 => x"56",
          8014 => x"76",
          8015 => x"51",
          8016 => x"27",
          8017 => x"70",
          8018 => x"5a",
          8019 => x"76",
          8020 => x"74",
          8021 => x"83",
          8022 => x"73",
          8023 => x"38",
          8024 => x"51",
          8025 => x"82",
          8026 => x"85",
          8027 => x"8e",
          8028 => x"2a",
          8029 => x"08",
          8030 => x"0c",
          8031 => x"79",
          8032 => x"73",
          8033 => x"0c",
          8034 => x"04",
          8035 => x"60",
          8036 => x"40",
          8037 => x"80",
          8038 => x"3d",
          8039 => x"78",
          8040 => x"3f",
          8041 => x"08",
          8042 => x"98",
          8043 => x"91",
          8044 => x"74",
          8045 => x"38",
          8046 => x"c7",
          8047 => x"33",
          8048 => x"87",
          8049 => x"2e",
          8050 => x"95",
          8051 => x"91",
          8052 => x"56",
          8053 => x"81",
          8054 => x"34",
          8055 => x"a3",
          8056 => x"08",
          8057 => x"31",
          8058 => x"27",
          8059 => x"5c",
          8060 => x"82",
          8061 => x"19",
          8062 => x"ff",
          8063 => x"74",
          8064 => x"7e",
          8065 => x"ff",
          8066 => x"2a",
          8067 => x"79",
          8068 => x"87",
          8069 => x"08",
          8070 => x"98",
          8071 => x"78",
          8072 => x"3f",
          8073 => x"08",
          8074 => x"27",
          8075 => x"74",
          8076 => x"a3",
          8077 => x"1a",
          8078 => x"08",
          8079 => x"c3",
          8080 => x"e0",
          8081 => x"2e",
          8082 => x"82",
          8083 => x"1a",
          8084 => x"59",
          8085 => x"2e",
          8086 => x"77",
          8087 => x"11",
          8088 => x"55",
          8089 => x"85",
          8090 => x"31",
          8091 => x"76",
          8092 => x"81",
          8093 => x"ff",
          8094 => x"82",
          8095 => x"fe",
          8096 => x"83",
          8097 => x"56",
          8098 => x"a0",
          8099 => x"08",
          8100 => x"74",
          8101 => x"38",
          8102 => x"b8",
          8103 => x"16",
          8104 => x"89",
          8105 => x"51",
          8106 => x"3f",
          8107 => x"56",
          8108 => x"9c",
          8109 => x"19",
          8110 => x"06",
          8111 => x"31",
          8112 => x"76",
          8113 => x"7b",
          8114 => x"08",
          8115 => x"c0",
          8116 => x"e0",
          8117 => x"ff",
          8118 => x"94",
          8119 => x"ff",
          8120 => x"05",
          8121 => x"ff",
          8122 => x"7b",
          8123 => x"08",
          8124 => x"76",
          8125 => x"08",
          8126 => x"0c",
          8127 => x"f0",
          8128 => x"75",
          8129 => x"0c",
          8130 => x"04",
          8131 => x"60",
          8132 => x"40",
          8133 => x"80",
          8134 => x"3d",
          8135 => x"77",
          8136 => x"3f",
          8137 => x"08",
          8138 => x"98",
          8139 => x"91",
          8140 => x"74",
          8141 => x"38",
          8142 => x"bf",
          8143 => x"33",
          8144 => x"70",
          8145 => x"56",
          8146 => x"74",
          8147 => x"ab",
          8148 => x"82",
          8149 => x"34",
          8150 => x"9f",
          8151 => x"91",
          8152 => x"56",
          8153 => x"94",
          8154 => x"11",
          8155 => x"76",
          8156 => x"75",
          8157 => x"80",
          8158 => x"38",
          8159 => x"70",
          8160 => x"56",
          8161 => x"82",
          8162 => x"11",
          8163 => x"77",
          8164 => x"5c",
          8165 => x"38",
          8166 => x"88",
          8167 => x"74",
          8168 => x"52",
          8169 => x"18",
          8170 => x"51",
          8171 => x"82",
          8172 => x"55",
          8173 => x"08",
          8174 => x"b2",
          8175 => x"2e",
          8176 => x"74",
          8177 => x"95",
          8178 => x"19",
          8179 => x"08",
          8180 => x"88",
          8181 => x"55",
          8182 => x"9c",
          8183 => x"09",
          8184 => x"38",
          8185 => x"bd",
          8186 => x"e0",
          8187 => x"ed",
          8188 => x"08",
          8189 => x"ff",
          8190 => x"82",
          8191 => x"80",
          8192 => x"38",
          8193 => x"08",
          8194 => x"2a",
          8195 => x"80",
          8196 => x"38",
          8197 => x"8a",
          8198 => x"5b",
          8199 => x"27",
          8200 => x"7b",
          8201 => x"54",
          8202 => x"52",
          8203 => x"51",
          8204 => x"3f",
          8205 => x"08",
          8206 => x"7e",
          8207 => x"78",
          8208 => x"74",
          8209 => x"38",
          8210 => x"b4",
          8211 => x"31",
          8212 => x"05",
          8213 => x"51",
          8214 => x"3f",
          8215 => x"0b",
          8216 => x"78",
          8217 => x"80",
          8218 => x"18",
          8219 => x"08",
          8220 => x"7e",
          8221 => x"f6",
          8222 => x"98",
          8223 => x"38",
          8224 => x"12",
          8225 => x"9c",
          8226 => x"18",
          8227 => x"06",
          8228 => x"31",
          8229 => x"76",
          8230 => x"7b",
          8231 => x"08",
          8232 => x"ff",
          8233 => x"82",
          8234 => x"fd",
          8235 => x"53",
          8236 => x"18",
          8237 => x"06",
          8238 => x"51",
          8239 => x"3f",
          8240 => x"0b",
          8241 => x"7b",
          8242 => x"08",
          8243 => x"76",
          8244 => x"08",
          8245 => x"1c",
          8246 => x"08",
          8247 => x"5c",
          8248 => x"83",
          8249 => x"74",
          8250 => x"fd",
          8251 => x"18",
          8252 => x"07",
          8253 => x"19",
          8254 => x"75",
          8255 => x"0c",
          8256 => x"04",
          8257 => x"7a",
          8258 => x"05",
          8259 => x"56",
          8260 => x"82",
          8261 => x"57",
          8262 => x"08",
          8263 => x"90",
          8264 => x"86",
          8265 => x"06",
          8266 => x"73",
          8267 => x"ee",
          8268 => x"08",
          8269 => x"ff",
          8270 => x"82",
          8271 => x"57",
          8272 => x"08",
          8273 => x"a4",
          8274 => x"11",
          8275 => x"55",
          8276 => x"16",
          8277 => x"08",
          8278 => x"75",
          8279 => x"a5",
          8280 => x"08",
          8281 => x"51",
          8282 => x"3f",
          8283 => x"0a",
          8284 => x"51",
          8285 => x"3f",
          8286 => x"15",
          8287 => x"c6",
          8288 => x"81",
          8289 => x"34",
          8290 => x"bb",
          8291 => x"e0",
          8292 => x"17",
          8293 => x"06",
          8294 => x"90",
          8295 => x"82",
          8296 => x"8a",
          8297 => x"fc",
          8298 => x"70",
          8299 => x"d4",
          8300 => x"98",
          8301 => x"e0",
          8302 => x"38",
          8303 => x"05",
          8304 => x"f1",
          8305 => x"e0",
          8306 => x"82",
          8307 => x"87",
          8308 => x"98",
          8309 => x"72",
          8310 => x"0c",
          8311 => x"04",
          8312 => x"84",
          8313 => x"89",
          8314 => x"80",
          8315 => x"98",
          8316 => x"38",
          8317 => x"08",
          8318 => x"34",
          8319 => x"82",
          8320 => x"83",
          8321 => x"ee",
          8322 => x"53",
          8323 => x"05",
          8324 => x"51",
          8325 => x"82",
          8326 => x"55",
          8327 => x"08",
          8328 => x"76",
          8329 => x"94",
          8330 => x"51",
          8331 => x"82",
          8332 => x"55",
          8333 => x"08",
          8334 => x"80",
          8335 => x"70",
          8336 => x"56",
          8337 => x"89",
          8338 => x"98",
          8339 => x"b2",
          8340 => x"05",
          8341 => x"2a",
          8342 => x"51",
          8343 => x"80",
          8344 => x"76",
          8345 => x"52",
          8346 => x"3f",
          8347 => x"08",
          8348 => x"8e",
          8349 => x"98",
          8350 => x"09",
          8351 => x"38",
          8352 => x"82",
          8353 => x"94",
          8354 => x"ff",
          8355 => x"80",
          8356 => x"80",
          8357 => x"5b",
          8358 => x"34",
          8359 => x"df",
          8360 => x"05",
          8361 => x"3d",
          8362 => x"3f",
          8363 => x"08",
          8364 => x"98",
          8365 => x"38",
          8366 => x"3d",
          8367 => x"98",
          8368 => x"d8",
          8369 => x"58",
          8370 => x"08",
          8371 => x"2e",
          8372 => x"a0",
          8373 => x"3d",
          8374 => x"c4",
          8375 => x"e0",
          8376 => x"82",
          8377 => x"82",
          8378 => x"d9",
          8379 => x"7b",
          8380 => x"ea",
          8381 => x"98",
          8382 => x"e0",
          8383 => x"d8",
          8384 => x"3d",
          8385 => x"51",
          8386 => x"82",
          8387 => x"80",
          8388 => x"76",
          8389 => x"c3",
          8390 => x"e0",
          8391 => x"82",
          8392 => x"82",
          8393 => x"52",
          8394 => x"b6",
          8395 => x"98",
          8396 => x"e0",
          8397 => x"38",
          8398 => x"08",
          8399 => x"c8",
          8400 => x"82",
          8401 => x"2e",
          8402 => x"52",
          8403 => x"e8",
          8404 => x"98",
          8405 => x"e0",
          8406 => x"2e",
          8407 => x"84",
          8408 => x"06",
          8409 => x"57",
          8410 => x"76",
          8411 => x"80",
          8412 => x"b8",
          8413 => x"51",
          8414 => x"76",
          8415 => x"11",
          8416 => x"51",
          8417 => x"73",
          8418 => x"38",
          8419 => x"05",
          8420 => x"81",
          8421 => x"56",
          8422 => x"f5",
          8423 => x"54",
          8424 => x"81",
          8425 => x"80",
          8426 => x"78",
          8427 => x"55",
          8428 => x"e1",
          8429 => x"ff",
          8430 => x"58",
          8431 => x"74",
          8432 => x"75",
          8433 => x"18",
          8434 => x"08",
          8435 => x"af",
          8436 => x"f4",
          8437 => x"2e",
          8438 => x"8d",
          8439 => x"80",
          8440 => x"11",
          8441 => x"74",
          8442 => x"82",
          8443 => x"70",
          8444 => x"d2",
          8445 => x"08",
          8446 => x"5c",
          8447 => x"73",
          8448 => x"38",
          8449 => x"1a",
          8450 => x"55",
          8451 => x"38",
          8452 => x"73",
          8453 => x"38",
          8454 => x"76",
          8455 => x"74",
          8456 => x"33",
          8457 => x"05",
          8458 => x"15",
          8459 => x"ba",
          8460 => x"05",
          8461 => x"ff",
          8462 => x"06",
          8463 => x"57",
          8464 => x"e0",
          8465 => x"81",
          8466 => x"73",
          8467 => x"81",
          8468 => x"7a",
          8469 => x"38",
          8470 => x"76",
          8471 => x"0c",
          8472 => x"0d",
          8473 => x"0d",
          8474 => x"3d",
          8475 => x"71",
          8476 => x"eb",
          8477 => x"e0",
          8478 => x"82",
          8479 => x"82",
          8480 => x"15",
          8481 => x"82",
          8482 => x"15",
          8483 => x"76",
          8484 => x"90",
          8485 => x"81",
          8486 => x"06",
          8487 => x"72",
          8488 => x"56",
          8489 => x"54",
          8490 => x"17",
          8491 => x"78",
          8492 => x"38",
          8493 => x"22",
          8494 => x"59",
          8495 => x"78",
          8496 => x"76",
          8497 => x"51",
          8498 => x"3f",
          8499 => x"08",
          8500 => x"54",
          8501 => x"53",
          8502 => x"3f",
          8503 => x"08",
          8504 => x"38",
          8505 => x"75",
          8506 => x"18",
          8507 => x"31",
          8508 => x"57",
          8509 => x"b2",
          8510 => x"08",
          8511 => x"38",
          8512 => x"51",
          8513 => x"3f",
          8514 => x"08",
          8515 => x"98",
          8516 => x"81",
          8517 => x"e0",
          8518 => x"2e",
          8519 => x"82",
          8520 => x"88",
          8521 => x"98",
          8522 => x"80",
          8523 => x"38",
          8524 => x"80",
          8525 => x"77",
          8526 => x"08",
          8527 => x"0c",
          8528 => x"70",
          8529 => x"81",
          8530 => x"5a",
          8531 => x"2e",
          8532 => x"52",
          8533 => x"bb",
          8534 => x"e0",
          8535 => x"82",
          8536 => x"95",
          8537 => x"98",
          8538 => x"39",
          8539 => x"51",
          8540 => x"3f",
          8541 => x"08",
          8542 => x"2e",
          8543 => x"74",
          8544 => x"79",
          8545 => x"14",
          8546 => x"38",
          8547 => x"0c",
          8548 => x"94",
          8549 => x"94",
          8550 => x"83",
          8551 => x"72",
          8552 => x"38",
          8553 => x"51",
          8554 => x"3f",
          8555 => x"08",
          8556 => x"0b",
          8557 => x"82",
          8558 => x"39",
          8559 => x"16",
          8560 => x"bb",
          8561 => x"2a",
          8562 => x"08",
          8563 => x"15",
          8564 => x"15",
          8565 => x"90",
          8566 => x"16",
          8567 => x"33",
          8568 => x"53",
          8569 => x"34",
          8570 => x"06",
          8571 => x"2e",
          8572 => x"9c",
          8573 => x"85",
          8574 => x"16",
          8575 => x"72",
          8576 => x"0c",
          8577 => x"04",
          8578 => x"79",
          8579 => x"75",
          8580 => x"8b",
          8581 => x"89",
          8582 => x"52",
          8583 => x"05",
          8584 => x"3f",
          8585 => x"08",
          8586 => x"98",
          8587 => x"38",
          8588 => x"7a",
          8589 => x"d4",
          8590 => x"e0",
          8591 => x"82",
          8592 => x"80",
          8593 => x"16",
          8594 => x"2b",
          8595 => x"74",
          8596 => x"86",
          8597 => x"84",
          8598 => x"06",
          8599 => x"73",
          8600 => x"38",
          8601 => x"52",
          8602 => x"e0",
          8603 => x"98",
          8604 => x"0c",
          8605 => x"14",
          8606 => x"23",
          8607 => x"51",
          8608 => x"3f",
          8609 => x"08",
          8610 => x"2e",
          8611 => x"85",
          8612 => x"86",
          8613 => x"2e",
          8614 => x"76",
          8615 => x"73",
          8616 => x"0c",
          8617 => x"04",
          8618 => x"76",
          8619 => x"05",
          8620 => x"53",
          8621 => x"82",
          8622 => x"87",
          8623 => x"98",
          8624 => x"86",
          8625 => x"fb",
          8626 => x"79",
          8627 => x"05",
          8628 => x"56",
          8629 => x"3f",
          8630 => x"08",
          8631 => x"98",
          8632 => x"38",
          8633 => x"82",
          8634 => x"52",
          8635 => x"bb",
          8636 => x"e0",
          8637 => x"80",
          8638 => x"e0",
          8639 => x"73",
          8640 => x"3f",
          8641 => x"08",
          8642 => x"98",
          8643 => x"09",
          8644 => x"38",
          8645 => x"39",
          8646 => x"08",
          8647 => x"52",
          8648 => x"f6",
          8649 => x"73",
          8650 => x"8c",
          8651 => x"98",
          8652 => x"70",
          8653 => x"07",
          8654 => x"82",
          8655 => x"06",
          8656 => x"54",
          8657 => x"98",
          8658 => x"0d",
          8659 => x"0d",
          8660 => x"53",
          8661 => x"53",
          8662 => x"56",
          8663 => x"82",
          8664 => x"55",
          8665 => x"08",
          8666 => x"52",
          8667 => x"a6",
          8668 => x"98",
          8669 => x"e0",
          8670 => x"38",
          8671 => x"05",
          8672 => x"2b",
          8673 => x"80",
          8674 => x"86",
          8675 => x"76",
          8676 => x"38",
          8677 => x"51",
          8678 => x"74",
          8679 => x"0c",
          8680 => x"04",
          8681 => x"63",
          8682 => x"80",
          8683 => x"ec",
          8684 => x"3d",
          8685 => x"3f",
          8686 => x"08",
          8687 => x"98",
          8688 => x"38",
          8689 => x"73",
          8690 => x"08",
          8691 => x"13",
          8692 => x"58",
          8693 => x"26",
          8694 => x"7c",
          8695 => x"39",
          8696 => x"ce",
          8697 => x"81",
          8698 => x"e0",
          8699 => x"33",
          8700 => x"81",
          8701 => x"06",
          8702 => x"82",
          8703 => x"76",
          8704 => x"f0",
          8705 => x"af",
          8706 => x"e0",
          8707 => x"2e",
          8708 => x"e0",
          8709 => x"2e",
          8710 => x"e0",
          8711 => x"70",
          8712 => x"08",
          8713 => x"7a",
          8714 => x"7f",
          8715 => x"54",
          8716 => x"77",
          8717 => x"80",
          8718 => x"15",
          8719 => x"98",
          8720 => x"75",
          8721 => x"52",
          8722 => x"52",
          8723 => x"8e",
          8724 => x"98",
          8725 => x"e0",
          8726 => x"d6",
          8727 => x"33",
          8728 => x"1a",
          8729 => x"54",
          8730 => x"09",
          8731 => x"38",
          8732 => x"ff",
          8733 => x"82",
          8734 => x"83",
          8735 => x"70",
          8736 => x"25",
          8737 => x"59",
          8738 => x"9b",
          8739 => x"51",
          8740 => x"3f",
          8741 => x"08",
          8742 => x"70",
          8743 => x"25",
          8744 => x"59",
          8745 => x"75",
          8746 => x"7a",
          8747 => x"ff",
          8748 => x"7c",
          8749 => x"94",
          8750 => x"11",
          8751 => x"56",
          8752 => x"15",
          8753 => x"e0",
          8754 => x"3d",
          8755 => x"3d",
          8756 => x"3d",
          8757 => x"70",
          8758 => x"95",
          8759 => x"98",
          8760 => x"e0",
          8761 => x"aa",
          8762 => x"33",
          8763 => x"a2",
          8764 => x"33",
          8765 => x"70",
          8766 => x"55",
          8767 => x"73",
          8768 => x"90",
          8769 => x"08",
          8770 => x"18",
          8771 => x"82",
          8772 => x"38",
          8773 => x"08",
          8774 => x"08",
          8775 => x"ff",
          8776 => x"82",
          8777 => x"74",
          8778 => x"56",
          8779 => x"98",
          8780 => x"76",
          8781 => x"c6",
          8782 => x"98",
          8783 => x"09",
          8784 => x"38",
          8785 => x"e0",
          8786 => x"2e",
          8787 => x"85",
          8788 => x"a4",
          8789 => x"38",
          8790 => x"e0",
          8791 => x"15",
          8792 => x"38",
          8793 => x"53",
          8794 => x"08",
          8795 => x"ff",
          8796 => x"82",
          8797 => x"56",
          8798 => x"8c",
          8799 => x"17",
          8800 => x"07",
          8801 => x"18",
          8802 => x"2e",
          8803 => x"91",
          8804 => x"55",
          8805 => x"98",
          8806 => x"0d",
          8807 => x"0d",
          8808 => x"3d",
          8809 => x"52",
          8810 => x"d9",
          8811 => x"e0",
          8812 => x"82",
          8813 => x"81",
          8814 => x"46",
          8815 => x"52",
          8816 => x"52",
          8817 => x"3f",
          8818 => x"08",
          8819 => x"98",
          8820 => x"38",
          8821 => x"05",
          8822 => x"2a",
          8823 => x"51",
          8824 => x"55",
          8825 => x"38",
          8826 => x"54",
          8827 => x"81",
          8828 => x"80",
          8829 => x"70",
          8830 => x"54",
          8831 => x"81",
          8832 => x"52",
          8833 => x"ba",
          8834 => x"e0",
          8835 => x"84",
          8836 => x"06",
          8837 => x"73",
          8838 => x"d6",
          8839 => x"82",
          8840 => x"98",
          8841 => x"81",
          8842 => x"5a",
          8843 => x"08",
          8844 => x"8a",
          8845 => x"54",
          8846 => x"3f",
          8847 => x"08",
          8848 => x"98",
          8849 => x"38",
          8850 => x"08",
          8851 => x"ff",
          8852 => x"82",
          8853 => x"55",
          8854 => x"08",
          8855 => x"55",
          8856 => x"82",
          8857 => x"84",
          8858 => x"82",
          8859 => x"80",
          8860 => x"51",
          8861 => x"82",
          8862 => x"82",
          8863 => x"30",
          8864 => x"98",
          8865 => x"25",
          8866 => x"75",
          8867 => x"38",
          8868 => x"90",
          8869 => x"75",
          8870 => x"ff",
          8871 => x"82",
          8872 => x"55",
          8873 => x"78",
          8874 => x"f9",
          8875 => x"98",
          8876 => x"82",
          8877 => x"a2",
          8878 => x"e8",
          8879 => x"53",
          8880 => x"bc",
          8881 => x"3d",
          8882 => x"3f",
          8883 => x"08",
          8884 => x"98",
          8885 => x"38",
          8886 => x"52",
          8887 => x"52",
          8888 => x"3f",
          8889 => x"08",
          8890 => x"98",
          8891 => x"88",
          8892 => x"39",
          8893 => x"08",
          8894 => x"81",
          8895 => x"38",
          8896 => x"05",
          8897 => x"2a",
          8898 => x"55",
          8899 => x"81",
          8900 => x"5a",
          8901 => x"3d",
          8902 => x"ff",
          8903 => x"82",
          8904 => x"75",
          8905 => x"e0",
          8906 => x"38",
          8907 => x"e0",
          8908 => x"2e",
          8909 => x"83",
          8910 => x"82",
          8911 => x"ff",
          8912 => x"06",
          8913 => x"54",
          8914 => x"73",
          8915 => x"82",
          8916 => x"52",
          8917 => x"b2",
          8918 => x"e0",
          8919 => x"82",
          8920 => x"81",
          8921 => x"53",
          8922 => x"19",
          8923 => x"c6",
          8924 => x"ae",
          8925 => x"34",
          8926 => x"0b",
          8927 => x"34",
          8928 => x"0a",
          8929 => x"19",
          8930 => x"d8",
          8931 => x"78",
          8932 => x"51",
          8933 => x"3f",
          8934 => x"b8",
          8935 => x"d8",
          8936 => x"a3",
          8937 => x"54",
          8938 => x"d9",
          8939 => x"53",
          8940 => x"11",
          8941 => x"b7",
          8942 => x"54",
          8943 => x"15",
          8944 => x"ff",
          8945 => x"82",
          8946 => x"54",
          8947 => x"08",
          8948 => x"88",
          8949 => x"64",
          8950 => x"ff",
          8951 => x"75",
          8952 => x"78",
          8953 => x"9d",
          8954 => x"90",
          8955 => x"34",
          8956 => x"0b",
          8957 => x"78",
          8958 => x"a9",
          8959 => x"98",
          8960 => x"39",
          8961 => x"52",
          8962 => x"ac",
          8963 => x"82",
          8964 => x"9a",
          8965 => x"d8",
          8966 => x"3d",
          8967 => x"d1",
          8968 => x"53",
          8969 => x"fc",
          8970 => x"3d",
          8971 => x"3f",
          8972 => x"08",
          8973 => x"98",
          8974 => x"38",
          8975 => x"3d",
          8976 => x"3d",
          8977 => x"c8",
          8978 => x"e0",
          8979 => x"82",
          8980 => x"82",
          8981 => x"81",
          8982 => x"81",
          8983 => x"86",
          8984 => x"af",
          8985 => x"a5",
          8986 => x"aa",
          8987 => x"05",
          8988 => x"9f",
          8989 => x"77",
          8990 => x"70",
          8991 => x"a2",
          8992 => x"3d",
          8993 => x"51",
          8994 => x"82",
          8995 => x"55",
          8996 => x"08",
          8997 => x"a1",
          8998 => x"09",
          8999 => x"38",
          9000 => x"08",
          9001 => x"88",
          9002 => x"39",
          9003 => x"08",
          9004 => x"81",
          9005 => x"38",
          9006 => x"bd",
          9007 => x"e0",
          9008 => x"82",
          9009 => x"81",
          9010 => x"56",
          9011 => x"3d",
          9012 => x"52",
          9013 => x"ff",
          9014 => x"02",
          9015 => x"8b",
          9016 => x"16",
          9017 => x"2a",
          9018 => x"51",
          9019 => x"89",
          9020 => x"07",
          9021 => x"17",
          9022 => x"81",
          9023 => x"34",
          9024 => x"70",
          9025 => x"81",
          9026 => x"55",
          9027 => x"80",
          9028 => x"64",
          9029 => x"38",
          9030 => x"51",
          9031 => x"3f",
          9032 => x"08",
          9033 => x"ff",
          9034 => x"82",
          9035 => x"98",
          9036 => x"80",
          9037 => x"e0",
          9038 => x"78",
          9039 => x"9e",
          9040 => x"98",
          9041 => x"d8",
          9042 => x"55",
          9043 => x"08",
          9044 => x"81",
          9045 => x"73",
          9046 => x"81",
          9047 => x"63",
          9048 => x"76",
          9049 => x"9d",
          9050 => x"81",
          9051 => x"34",
          9052 => x"e0",
          9053 => x"38",
          9054 => x"a5",
          9055 => x"98",
          9056 => x"e0",
          9057 => x"38",
          9058 => x"a3",
          9059 => x"e0",
          9060 => x"74",
          9061 => x"0c",
          9062 => x"04",
          9063 => x"02",
          9064 => x"33",
          9065 => x"80",
          9066 => x"57",
          9067 => x"96",
          9068 => x"52",
          9069 => x"d1",
          9070 => x"e0",
          9071 => x"82",
          9072 => x"80",
          9073 => x"5a",
          9074 => x"3d",
          9075 => x"c5",
          9076 => x"e0",
          9077 => x"82",
          9078 => x"b8",
          9079 => x"cf",
          9080 => x"a0",
          9081 => x"55",
          9082 => x"75",
          9083 => x"71",
          9084 => x"33",
          9085 => x"74",
          9086 => x"57",
          9087 => x"8b",
          9088 => x"54",
          9089 => x"15",
          9090 => x"ff",
          9091 => x"82",
          9092 => x"55",
          9093 => x"98",
          9094 => x"0d",
          9095 => x"0d",
          9096 => x"53",
          9097 => x"05",
          9098 => x"51",
          9099 => x"82",
          9100 => x"55",
          9101 => x"08",
          9102 => x"76",
          9103 => x"94",
          9104 => x"51",
          9105 => x"82",
          9106 => x"55",
          9107 => x"08",
          9108 => x"80",
          9109 => x"81",
          9110 => x"86",
          9111 => x"38",
          9112 => x"86",
          9113 => x"90",
          9114 => x"54",
          9115 => x"ff",
          9116 => x"76",
          9117 => x"83",
          9118 => x"51",
          9119 => x"3f",
          9120 => x"08",
          9121 => x"e0",
          9122 => x"3d",
          9123 => x"3d",
          9124 => x"5c",
          9125 => x"99",
          9126 => x"52",
          9127 => x"cf",
          9128 => x"e0",
          9129 => x"e0",
          9130 => x"70",
          9131 => x"08",
          9132 => x"51",
          9133 => x"80",
          9134 => x"38",
          9135 => x"06",
          9136 => x"80",
          9137 => x"38",
          9138 => x"5f",
          9139 => x"3d",
          9140 => x"ff",
          9141 => x"82",
          9142 => x"57",
          9143 => x"08",
          9144 => x"74",
          9145 => x"ff",
          9146 => x"82",
          9147 => x"57",
          9148 => x"08",
          9149 => x"e0",
          9150 => x"e0",
          9151 => x"5b",
          9152 => x"18",
          9153 => x"18",
          9154 => x"74",
          9155 => x"81",
          9156 => x"78",
          9157 => x"8b",
          9158 => x"54",
          9159 => x"75",
          9160 => x"38",
          9161 => x"1b",
          9162 => x"55",
          9163 => x"2e",
          9164 => x"39",
          9165 => x"09",
          9166 => x"38",
          9167 => x"80",
          9168 => x"70",
          9169 => x"25",
          9170 => x"80",
          9171 => x"38",
          9172 => x"bc",
          9173 => x"11",
          9174 => x"ff",
          9175 => x"82",
          9176 => x"57",
          9177 => x"08",
          9178 => x"70",
          9179 => x"80",
          9180 => x"83",
          9181 => x"80",
          9182 => x"84",
          9183 => x"a7",
          9184 => x"b8",
          9185 => x"9b",
          9186 => x"e0",
          9187 => x"0c",
          9188 => x"98",
          9189 => x"0d",
          9190 => x"0d",
          9191 => x"3d",
          9192 => x"52",
          9193 => x"cd",
          9194 => x"e0",
          9195 => x"e0",
          9196 => x"54",
          9197 => x"08",
          9198 => x"8b",
          9199 => x"8a",
          9200 => x"58",
          9201 => x"3f",
          9202 => x"33",
          9203 => x"9f",
          9204 => x"86",
          9205 => x"9d",
          9206 => x"9c",
          9207 => x"e0",
          9208 => x"ff",
          9209 => x"c4",
          9210 => x"98",
          9211 => x"c0",
          9212 => x"52",
          9213 => x"08",
          9214 => x"3f",
          9215 => x"08",
          9216 => x"06",
          9217 => x"2e",
          9218 => x"52",
          9219 => x"51",
          9220 => x"3f",
          9221 => x"08",
          9222 => x"ff",
          9223 => x"38",
          9224 => x"88",
          9225 => x"8a",
          9226 => x"38",
          9227 => x"e7",
          9228 => x"75",
          9229 => x"74",
          9230 => x"73",
          9231 => x"05",
          9232 => x"16",
          9233 => x"70",
          9234 => x"34",
          9235 => x"70",
          9236 => x"56",
          9237 => x"fe",
          9238 => x"3d",
          9239 => x"55",
          9240 => x"2e",
          9241 => x"75",
          9242 => x"38",
          9243 => x"55",
          9244 => x"33",
          9245 => x"a0",
          9246 => x"06",
          9247 => x"16",
          9248 => x"38",
          9249 => x"42",
          9250 => x"3d",
          9251 => x"ff",
          9252 => x"82",
          9253 => x"54",
          9254 => x"08",
          9255 => x"81",
          9256 => x"ff",
          9257 => x"82",
          9258 => x"54",
          9259 => x"08",
          9260 => x"80",
          9261 => x"54",
          9262 => x"80",
          9263 => x"e0",
          9264 => x"2e",
          9265 => x"80",
          9266 => x"54",
          9267 => x"80",
          9268 => x"52",
          9269 => x"ab",
          9270 => x"e0",
          9271 => x"82",
          9272 => x"b1",
          9273 => x"82",
          9274 => x"52",
          9275 => x"99",
          9276 => x"54",
          9277 => x"15",
          9278 => x"77",
          9279 => x"ff",
          9280 => x"78",
          9281 => x"83",
          9282 => x"51",
          9283 => x"3f",
          9284 => x"08",
          9285 => x"74",
          9286 => x"0c",
          9287 => x"04",
          9288 => x"60",
          9289 => x"05",
          9290 => x"33",
          9291 => x"05",
          9292 => x"40",
          9293 => x"b9",
          9294 => x"98",
          9295 => x"e0",
          9296 => x"bd",
          9297 => x"33",
          9298 => x"b5",
          9299 => x"2e",
          9300 => x"1a",
          9301 => x"90",
          9302 => x"33",
          9303 => x"70",
          9304 => x"55",
          9305 => x"38",
          9306 => x"97",
          9307 => x"82",
          9308 => x"58",
          9309 => x"7e",
          9310 => x"70",
          9311 => x"55",
          9312 => x"56",
          9313 => x"cb",
          9314 => x"7d",
          9315 => x"70",
          9316 => x"2a",
          9317 => x"08",
          9318 => x"08",
          9319 => x"5d",
          9320 => x"77",
          9321 => x"9c",
          9322 => x"26",
          9323 => x"57",
          9324 => x"59",
          9325 => x"52",
          9326 => x"9c",
          9327 => x"15",
          9328 => x"9c",
          9329 => x"26",
          9330 => x"55",
          9331 => x"08",
          9332 => x"99",
          9333 => x"98",
          9334 => x"ff",
          9335 => x"e0",
          9336 => x"38",
          9337 => x"75",
          9338 => x"81",
          9339 => x"93",
          9340 => x"80",
          9341 => x"2e",
          9342 => x"ff",
          9343 => x"58",
          9344 => x"7d",
          9345 => x"38",
          9346 => x"55",
          9347 => x"b4",
          9348 => x"56",
          9349 => x"09",
          9350 => x"38",
          9351 => x"53",
          9352 => x"51",
          9353 => x"3f",
          9354 => x"08",
          9355 => x"98",
          9356 => x"38",
          9357 => x"ff",
          9358 => x"5c",
          9359 => x"84",
          9360 => x"5c",
          9361 => x"12",
          9362 => x"80",
          9363 => x"78",
          9364 => x"7c",
          9365 => x"90",
          9366 => x"c0",
          9367 => x"90",
          9368 => x"15",
          9369 => x"94",
          9370 => x"54",
          9371 => x"91",
          9372 => x"31",
          9373 => x"84",
          9374 => x"07",
          9375 => x"16",
          9376 => x"73",
          9377 => x"0c",
          9378 => x"04",
          9379 => x"6c",
          9380 => x"05",
          9381 => x"33",
          9382 => x"45",
          9383 => x"d1",
          9384 => x"80",
          9385 => x"98",
          9386 => x"a0",
          9387 => x"98",
          9388 => x"82",
          9389 => x"70",
          9390 => x"74",
          9391 => x"38",
          9392 => x"82",
          9393 => x"82",
          9394 => x"05",
          9395 => x"11",
          9396 => x"8d",
          9397 => x"41",
          9398 => x"7f",
          9399 => x"ac",
          9400 => x"98",
          9401 => x"06",
          9402 => x"56",
          9403 => x"74",
          9404 => x"76",
          9405 => x"81",
          9406 => x"8a",
          9407 => x"cc",
          9408 => x"fc",
          9409 => x"52",
          9410 => x"92",
          9411 => x"e0",
          9412 => x"38",
          9413 => x"80",
          9414 => x"74",
          9415 => x"26",
          9416 => x"15",
          9417 => x"74",
          9418 => x"38",
          9419 => x"80",
          9420 => x"84",
          9421 => x"92",
          9422 => x"80",
          9423 => x"38",
          9424 => x"06",
          9425 => x"2e",
          9426 => x"56",
          9427 => x"78",
          9428 => x"89",
          9429 => x"2b",
          9430 => x"43",
          9431 => x"38",
          9432 => x"30",
          9433 => x"77",
          9434 => x"91",
          9435 => x"dc",
          9436 => x"2e",
          9437 => x"81",
          9438 => x"7a",
          9439 => x"ff",
          9440 => x"81",
          9441 => x"98",
          9442 => x"38",
          9443 => x"51",
          9444 => x"3f",
          9445 => x"08",
          9446 => x"06",
          9447 => x"74",
          9448 => x"2e",
          9449 => x"8b",
          9450 => x"90",
          9451 => x"b2",
          9452 => x"57",
          9453 => x"8b",
          9454 => x"b6",
          9455 => x"92",
          9456 => x"e0",
          9457 => x"ba",
          9458 => x"ff",
          9459 => x"82",
          9460 => x"48",
          9461 => x"3d",
          9462 => x"81",
          9463 => x"ff",
          9464 => x"81",
          9465 => x"98",
          9466 => x"38",
          9467 => x"70",
          9468 => x"e0",
          9469 => x"51",
          9470 => x"38",
          9471 => x"55",
          9472 => x"75",
          9473 => x"38",
          9474 => x"48",
          9475 => x"ff",
          9476 => x"b8",
          9477 => x"78",
          9478 => x"8a",
          9479 => x"81",
          9480 => x"06",
          9481 => x"80",
          9482 => x"62",
          9483 => x"74",
          9484 => x"8d",
          9485 => x"06",
          9486 => x"2e",
          9487 => x"62",
          9488 => x"93",
          9489 => x"74",
          9490 => x"80",
          9491 => x"7d",
          9492 => x"81",
          9493 => x"38",
          9494 => x"67",
          9495 => x"81",
          9496 => x"dc",
          9497 => x"74",
          9498 => x"38",
          9499 => x"98",
          9500 => x"dc",
          9501 => x"82",
          9502 => x"57",
          9503 => x"80",
          9504 => x"76",
          9505 => x"38",
          9506 => x"51",
          9507 => x"3f",
          9508 => x"08",
          9509 => x"87",
          9510 => x"2a",
          9511 => x"5c",
          9512 => x"e0",
          9513 => x"80",
          9514 => x"46",
          9515 => x"0a",
          9516 => x"ec",
          9517 => x"39",
          9518 => x"67",
          9519 => x"81",
          9520 => x"cc",
          9521 => x"74",
          9522 => x"38",
          9523 => x"98",
          9524 => x"cc",
          9525 => x"82",
          9526 => x"57",
          9527 => x"80",
          9528 => x"76",
          9529 => x"38",
          9530 => x"51",
          9531 => x"3f",
          9532 => x"08",
          9533 => x"57",
          9534 => x"08",
          9535 => x"96",
          9536 => x"82",
          9537 => x"10",
          9538 => x"08",
          9539 => x"72",
          9540 => x"59",
          9541 => x"ff",
          9542 => x"5d",
          9543 => x"46",
          9544 => x"11",
          9545 => x"70",
          9546 => x"71",
          9547 => x"06",
          9548 => x"52",
          9549 => x"41",
          9550 => x"09",
          9551 => x"38",
          9552 => x"18",
          9553 => x"39",
          9554 => x"79",
          9555 => x"70",
          9556 => x"58",
          9557 => x"76",
          9558 => x"38",
          9559 => x"7d",
          9560 => x"70",
          9561 => x"55",
          9562 => x"3f",
          9563 => x"08",
          9564 => x"2e",
          9565 => x"9b",
          9566 => x"98",
          9567 => x"f5",
          9568 => x"38",
          9569 => x"38",
          9570 => x"59",
          9571 => x"38",
          9572 => x"7d",
          9573 => x"81",
          9574 => x"38",
          9575 => x"0b",
          9576 => x"08",
          9577 => x"78",
          9578 => x"1a",
          9579 => x"c0",
          9580 => x"74",
          9581 => x"39",
          9582 => x"55",
          9583 => x"8f",
          9584 => x"fd",
          9585 => x"e0",
          9586 => x"f5",
          9587 => x"78",
          9588 => x"79",
          9589 => x"80",
          9590 => x"f1",
          9591 => x"39",
          9592 => x"81",
          9593 => x"06",
          9594 => x"55",
          9595 => x"27",
          9596 => x"81",
          9597 => x"56",
          9598 => x"38",
          9599 => x"80",
          9600 => x"ff",
          9601 => x"8b",
          9602 => x"e4",
          9603 => x"ff",
          9604 => x"84",
          9605 => x"1b",
          9606 => x"aa",
          9607 => x"1c",
          9608 => x"ff",
          9609 => x"8e",
          9610 => x"8e",
          9611 => x"0b",
          9612 => x"7d",
          9613 => x"30",
          9614 => x"84",
          9615 => x"51",
          9616 => x"51",
          9617 => x"3f",
          9618 => x"83",
          9619 => x"90",
          9620 => x"ff",
          9621 => x"93",
          9622 => x"8d",
          9623 => x"39",
          9624 => x"1b",
          9625 => x"fc",
          9626 => x"95",
          9627 => x"52",
          9628 => x"ff",
          9629 => x"81",
          9630 => x"1b",
          9631 => x"c6",
          9632 => x"9c",
          9633 => x"8d",
          9634 => x"83",
          9635 => x"06",
          9636 => x"82",
          9637 => x"52",
          9638 => x"51",
          9639 => x"3f",
          9640 => x"1b",
          9641 => x"bc",
          9642 => x"ac",
          9643 => x"8d",
          9644 => x"52",
          9645 => x"ff",
          9646 => x"86",
          9647 => x"51",
          9648 => x"3f",
          9649 => x"80",
          9650 => x"a9",
          9651 => x"1c",
          9652 => x"82",
          9653 => x"80",
          9654 => x"ae",
          9655 => x"b2",
          9656 => x"1b",
          9657 => x"fc",
          9658 => x"ff",
          9659 => x"96",
          9660 => x"8c",
          9661 => x"80",
          9662 => x"34",
          9663 => x"1c",
          9664 => x"82",
          9665 => x"ab",
          9666 => x"8d",
          9667 => x"d4",
          9668 => x"fe",
          9669 => x"59",
          9670 => x"3f",
          9671 => x"53",
          9672 => x"51",
          9673 => x"3f",
          9674 => x"e0",
          9675 => x"9c",
          9676 => x"2e",
          9677 => x"80",
          9678 => x"54",
          9679 => x"7a",
          9680 => x"ff",
          9681 => x"84",
          9682 => x"52",
          9683 => x"8c",
          9684 => x"8b",
          9685 => x"52",
          9686 => x"8c",
          9687 => x"8a",
          9688 => x"52",
          9689 => x"51",
          9690 => x"3f",
          9691 => x"83",
          9692 => x"ff",
          9693 => x"82",
          9694 => x"1b",
          9695 => x"e4",
          9696 => x"d5",
          9697 => x"ff",
          9698 => x"75",
          9699 => x"53",
          9700 => x"51",
          9701 => x"3f",
          9702 => x"1f",
          9703 => x"7f",
          9704 => x"d1",
          9705 => x"80",
          9706 => x"ff",
          9707 => x"60",
          9708 => x"7d",
          9709 => x"81",
          9710 => x"f8",
          9711 => x"ff",
          9712 => x"ff",
          9713 => x"51",
          9714 => x"3f",
          9715 => x"88",
          9716 => x"39",
          9717 => x"f8",
          9718 => x"2e",
          9719 => x"55",
          9720 => x"51",
          9721 => x"3f",
          9722 => x"57",
          9723 => x"83",
          9724 => x"76",
          9725 => x"7a",
          9726 => x"ff",
          9727 => x"82",
          9728 => x"82",
          9729 => x"80",
          9730 => x"98",
          9731 => x"51",
          9732 => x"3f",
          9733 => x"78",
          9734 => x"74",
          9735 => x"18",
          9736 => x"2e",
          9737 => x"79",
          9738 => x"2e",
          9739 => x"55",
          9740 => x"62",
          9741 => x"74",
          9742 => x"75",
          9743 => x"7f",
          9744 => x"b1",
          9745 => x"98",
          9746 => x"38",
          9747 => x"78",
          9748 => x"74",
          9749 => x"57",
          9750 => x"93",
          9751 => x"67",
          9752 => x"26",
          9753 => x"57",
          9754 => x"83",
          9755 => x"64",
          9756 => x"38",
          9757 => x"53",
          9758 => x"51",
          9759 => x"3f",
          9760 => x"e0",
          9761 => x"c4",
          9762 => x"29",
          9763 => x"83",
          9764 => x"75",
          9765 => x"98",
          9766 => x"52",
          9767 => x"85",
          9768 => x"81",
          9769 => x"2a",
          9770 => x"77",
          9771 => x"84",
          9772 => x"52",
          9773 => x"89",
          9774 => x"d4",
          9775 => x"51",
          9776 => x"3f",
          9777 => x"55",
          9778 => x"81",
          9779 => x"34",
          9780 => x"16",
          9781 => x"16",
          9782 => x"16",
          9783 => x"56",
          9784 => x"52",
          9785 => x"93",
          9786 => x"0b",
          9787 => x"82",
          9788 => x"82",
          9789 => x"56",
          9790 => x"34",
          9791 => x"08",
          9792 => x"7e",
          9793 => x"1b",
          9794 => x"d8",
          9795 => x"83",
          9796 => x"ff",
          9797 => x"81",
          9798 => x"7a",
          9799 => x"ff",
          9800 => x"81",
          9801 => x"98",
          9802 => x"80",
          9803 => x"7f",
          9804 => x"a5",
          9805 => x"82",
          9806 => x"90",
          9807 => x"8e",
          9808 => x"81",
          9809 => x"82",
          9810 => x"56",
          9811 => x"98",
          9812 => x"0d",
          9813 => x"0d",
          9814 => x"59",
          9815 => x"ff",
          9816 => x"57",
          9817 => x"b4",
          9818 => x"f8",
          9819 => x"81",
          9820 => x"52",
          9821 => x"94",
          9822 => x"2e",
          9823 => x"9c",
          9824 => x"33",
          9825 => x"2e",
          9826 => x"76",
          9827 => x"58",
          9828 => x"57",
          9829 => x"09",
          9830 => x"38",
          9831 => x"78",
          9832 => x"38",
          9833 => x"82",
          9834 => x"8d",
          9835 => x"f7",
          9836 => x"02",
          9837 => x"05",
          9838 => x"77",
          9839 => x"81",
          9840 => x"8d",
          9841 => x"e7",
          9842 => x"08",
          9843 => x"24",
          9844 => x"17",
          9845 => x"8c",
          9846 => x"77",
          9847 => x"16",
          9848 => x"25",
          9849 => x"3d",
          9850 => x"75",
          9851 => x"52",
          9852 => x"ca",
          9853 => x"76",
          9854 => x"70",
          9855 => x"2a",
          9856 => x"51",
          9857 => x"84",
          9858 => x"19",
          9859 => x"8b",
          9860 => x"f9",
          9861 => x"84",
          9862 => x"56",
          9863 => x"a7",
          9864 => x"fc",
          9865 => x"53",
          9866 => x"75",
          9867 => x"dc",
          9868 => x"98",
          9869 => x"84",
          9870 => x"2e",
          9871 => x"87",
          9872 => x"08",
          9873 => x"ff",
          9874 => x"e0",
          9875 => x"3d",
          9876 => x"3d",
          9877 => x"80",
          9878 => x"52",
          9879 => x"86",
          9880 => x"74",
          9881 => x"0d",
          9882 => x"0d",
          9883 => x"05",
          9884 => x"86",
          9885 => x"54",
          9886 => x"73",
          9887 => x"fe",
          9888 => x"51",
          9889 => x"98",
          9890 => x"fd",
          9891 => x"02",
          9892 => x"05",
          9893 => x"80",
          9894 => x"ff",
          9895 => x"72",
          9896 => x"06",
          9897 => x"39",
          9898 => x"73",
          9899 => x"83",
          9900 => x"81",
          9901 => x"70",
          9902 => x"38",
          9903 => x"22",
          9904 => x"2e",
          9905 => x"12",
          9906 => x"ff",
          9907 => x"71",
          9908 => x"8d",
          9909 => x"82",
          9910 => x"70",
          9911 => x"e1",
          9912 => x"12",
          9913 => x"06",
          9914 => x"82",
          9915 => x"85",
          9916 => x"fe",
          9917 => x"92",
          9918 => x"84",
          9919 => x"22",
          9920 => x"53",
          9921 => x"26",
          9922 => x"53",
          9923 => x"83",
          9924 => x"81",
          9925 => x"70",
          9926 => x"8b",
          9927 => x"82",
          9928 => x"70",
          9929 => x"72",
          9930 => x"0c",
          9931 => x"04",
          9932 => x"77",
          9933 => x"ff",
          9934 => x"a7",
          9935 => x"ff",
          9936 => x"d5",
          9937 => x"9f",
          9938 => x"85",
          9939 => x"e0",
          9940 => x"82",
          9941 => x"70",
          9942 => x"25",
          9943 => x"07",
          9944 => x"70",
          9945 => x"75",
          9946 => x"57",
          9947 => x"2a",
          9948 => x"06",
          9949 => x"52",
          9950 => x"71",
          9951 => x"38",
          9952 => x"80",
          9953 => x"84",
          9954 => x"b8",
          9955 => x"08",
          9956 => x"31",
          9957 => x"70",
          9958 => x"51",
          9959 => x"71",
          9960 => x"06",
          9961 => x"51",
          9962 => x"f0",
          9963 => x"39",
          9964 => x"9a",
          9965 => x"51",
          9966 => x"12",
          9967 => x"88",
          9968 => x"39",
          9969 => x"51",
          9970 => x"a0",
          9971 => x"83",
          9972 => x"52",
          9973 => x"fe",
          9974 => x"10",
          9975 => x"f1",
          9976 => x"70",
          9977 => x"0c",
          9978 => x"04",
          9979 => x"ff",
          9980 => x"ff",
          9981 => x"ff",
          9982 => x"00",
          9983 => x"01",
          9984 => x"85",
          9985 => x"8c",
          9986 => x"93",
          9987 => x"9a",
          9988 => x"a1",
          9989 => x"a8",
          9990 => x"af",
          9991 => x"b6",
          9992 => x"bd",
          9993 => x"c4",
          9994 => x"cb",
          9995 => x"d1",
          9996 => x"d7",
          9997 => x"dd",
          9998 => x"e3",
          9999 => x"e9",
         10000 => x"ef",
         10001 => x"f5",
         10002 => x"fb",
         10003 => x"81",
         10004 => x"87",
         10005 => x"8d",
         10006 => x"93",
         10007 => x"99",
         10008 => x"79",
         10009 => x"79",
         10010 => x"8a",
         10011 => x"e2",
         10012 => x"61",
         10013 => x"4c",
         10014 => x"52",
         10015 => x"b3",
         10016 => x"95",
         10017 => x"2b",
         10018 => x"b1",
         10019 => x"34",
         10020 => x"4c",
         10021 => x"8a",
         10022 => x"b3",
         10023 => x"52",
         10024 => x"4c",
         10025 => x"4c",
         10026 => x"b1",
         10027 => x"2b",
         10028 => x"b3",
         10029 => x"e2",
         10030 => x"91",
         10031 => x"9f",
         10032 => x"ab",
         10033 => x"b0",
         10034 => x"b5",
         10035 => x"ba",
         10036 => x"bf",
         10037 => x"c4",
         10038 => x"ca",
         10039 => x"65",
         10040 => x"4e",
         10041 => x"4e",
         10042 => x"94",
         10043 => x"4e",
         10044 => x"4e",
         10045 => x"4e",
         10046 => x"4e",
         10047 => x"4e",
         10048 => x"4e",
         10049 => x"4e",
         10050 => x"51",
         10051 => x"4e",
         10052 => x"7c",
         10053 => x"ac",
         10054 => x"4e",
         10055 => x"4e",
         10056 => x"4e",
         10057 => x"4e",
         10058 => x"4e",
         10059 => x"4e",
         10060 => x"4e",
         10061 => x"4e",
         10062 => x"4e",
         10063 => x"4e",
         10064 => x"4e",
         10065 => x"4e",
         10066 => x"4e",
         10067 => x"4e",
         10068 => x"4e",
         10069 => x"4e",
         10070 => x"4e",
         10071 => x"4e",
         10072 => x"4e",
         10073 => x"4e",
         10074 => x"4e",
         10075 => x"4e",
         10076 => x"4e",
         10077 => x"4e",
         10078 => x"4e",
         10079 => x"4e",
         10080 => x"4e",
         10081 => x"4e",
         10082 => x"4e",
         10083 => x"4e",
         10084 => x"4e",
         10085 => x"4e",
         10086 => x"4e",
         10087 => x"4e",
         10088 => x"4e",
         10089 => x"4e",
         10090 => x"dc",
         10091 => x"4e",
         10092 => x"4e",
         10093 => x"4e",
         10094 => x"4e",
         10095 => x"4a",
         10096 => x"4e",
         10097 => x"4e",
         10098 => x"4e",
         10099 => x"4e",
         10100 => x"4e",
         10101 => x"4e",
         10102 => x"4e",
         10103 => x"4e",
         10104 => x"4e",
         10105 => x"4e",
         10106 => x"0c",
         10107 => x"73",
         10108 => x"e3",
         10109 => x"e3",
         10110 => x"e3",
         10111 => x"4e",
         10112 => x"73",
         10113 => x"4e",
         10114 => x"4e",
         10115 => x"cc",
         10116 => x"4e",
         10117 => x"4e",
         10118 => x"20",
         10119 => x"2b",
         10120 => x"4e",
         10121 => x"4e",
         10122 => x"45",
         10123 => x"4e",
         10124 => x"53",
         10125 => x"4e",
         10126 => x"4e",
         10127 => x"4a",
         10128 => x"69",
         10129 => x"00",
         10130 => x"63",
         10131 => x"00",
         10132 => x"69",
         10133 => x"00",
         10134 => x"61",
         10135 => x"00",
         10136 => x"65",
         10137 => x"00",
         10138 => x"65",
         10139 => x"00",
         10140 => x"70",
         10141 => x"00",
         10142 => x"66",
         10143 => x"00",
         10144 => x"6d",
         10145 => x"00",
         10146 => x"00",
         10147 => x"00",
         10148 => x"00",
         10149 => x"00",
         10150 => x"00",
         10151 => x"00",
         10152 => x"00",
         10153 => x"6c",
         10154 => x"00",
         10155 => x"00",
         10156 => x"74",
         10157 => x"00",
         10158 => x"65",
         10159 => x"00",
         10160 => x"6f",
         10161 => x"00",
         10162 => x"73",
         10163 => x"00",
         10164 => x"73",
         10165 => x"00",
         10166 => x"6f",
         10167 => x"00",
         10168 => x"00",
         10169 => x"6b",
         10170 => x"72",
         10171 => x"00",
         10172 => x"65",
         10173 => x"6c",
         10174 => x"72",
         10175 => x"00",
         10176 => x"6b",
         10177 => x"74",
         10178 => x"61",
         10179 => x"00",
         10180 => x"66",
         10181 => x"20",
         10182 => x"6e",
         10183 => x"00",
         10184 => x"70",
         10185 => x"20",
         10186 => x"6e",
         10187 => x"00",
         10188 => x"61",
         10189 => x"20",
         10190 => x"65",
         10191 => x"65",
         10192 => x"00",
         10193 => x"65",
         10194 => x"64",
         10195 => x"65",
         10196 => x"00",
         10197 => x"65",
         10198 => x"72",
         10199 => x"79",
         10200 => x"69",
         10201 => x"2e",
         10202 => x"00",
         10203 => x"65",
         10204 => x"6e",
         10205 => x"20",
         10206 => x"61",
         10207 => x"2e",
         10208 => x"00",
         10209 => x"69",
         10210 => x"72",
         10211 => x"20",
         10212 => x"74",
         10213 => x"65",
         10214 => x"00",
         10215 => x"76",
         10216 => x"75",
         10217 => x"72",
         10218 => x"20",
         10219 => x"61",
         10220 => x"2e",
         10221 => x"00",
         10222 => x"6b",
         10223 => x"74",
         10224 => x"61",
         10225 => x"64",
         10226 => x"00",
         10227 => x"63",
         10228 => x"61",
         10229 => x"6c",
         10230 => x"69",
         10231 => x"79",
         10232 => x"6d",
         10233 => x"75",
         10234 => x"6f",
         10235 => x"69",
         10236 => x"00",
         10237 => x"6d",
         10238 => x"61",
         10239 => x"74",
         10240 => x"00",
         10241 => x"65",
         10242 => x"2c",
         10243 => x"65",
         10244 => x"69",
         10245 => x"63",
         10246 => x"65",
         10247 => x"64",
         10248 => x"00",
         10249 => x"65",
         10250 => x"20",
         10251 => x"6b",
         10252 => x"00",
         10253 => x"75",
         10254 => x"63",
         10255 => x"74",
         10256 => x"6d",
         10257 => x"2e",
         10258 => x"00",
         10259 => x"20",
         10260 => x"79",
         10261 => x"65",
         10262 => x"69",
         10263 => x"2e",
         10264 => x"00",
         10265 => x"61",
         10266 => x"65",
         10267 => x"69",
         10268 => x"72",
         10269 => x"74",
         10270 => x"00",
         10271 => x"63",
         10272 => x"2e",
         10273 => x"00",
         10274 => x"6e",
         10275 => x"20",
         10276 => x"6f",
         10277 => x"00",
         10278 => x"75",
         10279 => x"74",
         10280 => x"25",
         10281 => x"74",
         10282 => x"75",
         10283 => x"74",
         10284 => x"73",
         10285 => x"0a",
         10286 => x"00",
         10287 => x"64",
         10288 => x"00",
         10289 => x"6c",
         10290 => x"00",
         10291 => x"00",
         10292 => x"58",
         10293 => x"00",
         10294 => x"20",
         10295 => x"20",
         10296 => x"00",
         10297 => x"58",
         10298 => x"00",
         10299 => x"00",
         10300 => x"00",
         10301 => x"00",
         10302 => x"00",
         10303 => x"25",
         10304 => x"00",
         10305 => x"31",
         10306 => x"30",
         10307 => x"00",
         10308 => x"31",
         10309 => x"00",
         10310 => x"55",
         10311 => x"65",
         10312 => x"30",
         10313 => x"20",
         10314 => x"25",
         10315 => x"2a",
         10316 => x"00",
         10317 => x"20",
         10318 => x"65",
         10319 => x"70",
         10320 => x"61",
         10321 => x"65",
         10322 => x"00",
         10323 => x"65",
         10324 => x"6e",
         10325 => x"72",
         10326 => x"00",
         10327 => x"20",
         10328 => x"65",
         10329 => x"70",
         10330 => x"00",
         10331 => x"54",
         10332 => x"44",
         10333 => x"74",
         10334 => x"75",
         10335 => x"00",
         10336 => x"54",
         10337 => x"52",
         10338 => x"74",
         10339 => x"75",
         10340 => x"00",
         10341 => x"54",
         10342 => x"58",
         10343 => x"74",
         10344 => x"75",
         10345 => x"00",
         10346 => x"54",
         10347 => x"58",
         10348 => x"74",
         10349 => x"75",
         10350 => x"00",
         10351 => x"54",
         10352 => x"58",
         10353 => x"74",
         10354 => x"75",
         10355 => x"00",
         10356 => x"54",
         10357 => x"58",
         10358 => x"74",
         10359 => x"75",
         10360 => x"00",
         10361 => x"74",
         10362 => x"20",
         10363 => x"74",
         10364 => x"72",
         10365 => x"00",
         10366 => x"62",
         10367 => x"67",
         10368 => x"6d",
         10369 => x"2e",
         10370 => x"00",
         10371 => x"6f",
         10372 => x"63",
         10373 => x"74",
         10374 => x"00",
         10375 => x"5f",
         10376 => x"2e",
         10377 => x"00",
         10378 => x"00",
         10379 => x"6c",
         10380 => x"74",
         10381 => x"6e",
         10382 => x"61",
         10383 => x"65",
         10384 => x"20",
         10385 => x"64",
         10386 => x"20",
         10387 => x"61",
         10388 => x"69",
         10389 => x"20",
         10390 => x"75",
         10391 => x"79",
         10392 => x"00",
         10393 => x"00",
         10394 => x"61",
         10395 => x"67",
         10396 => x"2e",
         10397 => x"00",
         10398 => x"79",
         10399 => x"2e",
         10400 => x"00",
         10401 => x"70",
         10402 => x"6e",
         10403 => x"2e",
         10404 => x"00",
         10405 => x"6c",
         10406 => x"30",
         10407 => x"2d",
         10408 => x"38",
         10409 => x"25",
         10410 => x"29",
         10411 => x"00",
         10412 => x"70",
         10413 => x"6d",
         10414 => x"00",
         10415 => x"6d",
         10416 => x"74",
         10417 => x"00",
         10418 => x"6c",
         10419 => x"30",
         10420 => x"00",
         10421 => x"00",
         10422 => x"6c",
         10423 => x"30",
         10424 => x"00",
         10425 => x"6c",
         10426 => x"30",
         10427 => x"2d",
         10428 => x"00",
         10429 => x"63",
         10430 => x"6e",
         10431 => x"6f",
         10432 => x"40",
         10433 => x"38",
         10434 => x"2e",
         10435 => x"00",
         10436 => x"6c",
         10437 => x"20",
         10438 => x"65",
         10439 => x"25",
         10440 => x"78",
         10441 => x"2e",
         10442 => x"00",
         10443 => x"6c",
         10444 => x"74",
         10445 => x"65",
         10446 => x"6f",
         10447 => x"28",
         10448 => x"2e",
         10449 => x"00",
         10450 => x"74",
         10451 => x"69",
         10452 => x"61",
         10453 => x"69",
         10454 => x"69",
         10455 => x"2e",
         10456 => x"00",
         10457 => x"64",
         10458 => x"62",
         10459 => x"69",
         10460 => x"2e",
         10461 => x"00",
         10462 => x"00",
         10463 => x"00",
         10464 => x"5c",
         10465 => x"25",
         10466 => x"73",
         10467 => x"00",
         10468 => x"5c",
         10469 => x"25",
         10470 => x"00",
         10471 => x"5c",
         10472 => x"00",
         10473 => x"20",
         10474 => x"6d",
         10475 => x"2e",
         10476 => x"00",
         10477 => x"6f",
         10478 => x"65",
         10479 => x"75",
         10480 => x"64",
         10481 => x"61",
         10482 => x"74",
         10483 => x"6f",
         10484 => x"73",
         10485 => x"6d",
         10486 => x"64",
         10487 => x"00",
         10488 => x"6e",
         10489 => x"2e",
         10490 => x"00",
         10491 => x"62",
         10492 => x"67",
         10493 => x"74",
         10494 => x"75",
         10495 => x"2e",
         10496 => x"00",
         10497 => x"25",
         10498 => x"64",
         10499 => x"3a",
         10500 => x"25",
         10501 => x"64",
         10502 => x"00",
         10503 => x"20",
         10504 => x"66",
         10505 => x"72",
         10506 => x"6f",
         10507 => x"00",
         10508 => x"72",
         10509 => x"53",
         10510 => x"63",
         10511 => x"69",
         10512 => x"00",
         10513 => x"65",
         10514 => x"65",
         10515 => x"6d",
         10516 => x"6d",
         10517 => x"65",
         10518 => x"00",
         10519 => x"20",
         10520 => x"53",
         10521 => x"4d",
         10522 => x"25",
         10523 => x"3a",
         10524 => x"58",
         10525 => x"00",
         10526 => x"20",
         10527 => x"41",
         10528 => x"20",
         10529 => x"25",
         10530 => x"3a",
         10531 => x"58",
         10532 => x"00",
         10533 => x"20",
         10534 => x"4e",
         10535 => x"41",
         10536 => x"25",
         10537 => x"3a",
         10538 => x"58",
         10539 => x"00",
         10540 => x"20",
         10541 => x"4d",
         10542 => x"20",
         10543 => x"25",
         10544 => x"3a",
         10545 => x"58",
         10546 => x"00",
         10547 => x"20",
         10548 => x"20",
         10549 => x"20",
         10550 => x"25",
         10551 => x"3a",
         10552 => x"58",
         10553 => x"00",
         10554 => x"20",
         10555 => x"43",
         10556 => x"20",
         10557 => x"44",
         10558 => x"63",
         10559 => x"3d",
         10560 => x"64",
         10561 => x"00",
         10562 => x"20",
         10563 => x"45",
         10564 => x"20",
         10565 => x"54",
         10566 => x"72",
         10567 => x"3d",
         10568 => x"64",
         10569 => x"00",
         10570 => x"20",
         10571 => x"52",
         10572 => x"52",
         10573 => x"43",
         10574 => x"6e",
         10575 => x"3d",
         10576 => x"64",
         10577 => x"00",
         10578 => x"20",
         10579 => x"48",
         10580 => x"45",
         10581 => x"53",
         10582 => x"00",
         10583 => x"20",
         10584 => x"49",
         10585 => x"00",
         10586 => x"20",
         10587 => x"54",
         10588 => x"00",
         10589 => x"20",
         10590 => x"00",
         10591 => x"20",
         10592 => x"00",
         10593 => x"72",
         10594 => x"65",
         10595 => x"00",
         10596 => x"20",
         10597 => x"20",
         10598 => x"65",
         10599 => x"65",
         10600 => x"72",
         10601 => x"64",
         10602 => x"73",
         10603 => x"25",
         10604 => x"0a",
         10605 => x"00",
         10606 => x"20",
         10607 => x"20",
         10608 => x"6f",
         10609 => x"53",
         10610 => x"74",
         10611 => x"64",
         10612 => x"73",
         10613 => x"25",
         10614 => x"0a",
         10615 => x"00",
         10616 => x"20",
         10617 => x"63",
         10618 => x"74",
         10619 => x"20",
         10620 => x"72",
         10621 => x"20",
         10622 => x"20",
         10623 => x"25",
         10624 => x"0a",
         10625 => x"00",
         10626 => x"63",
         10627 => x"00",
         10628 => x"20",
         10629 => x"20",
         10630 => x"20",
         10631 => x"20",
         10632 => x"20",
         10633 => x"20",
         10634 => x"20",
         10635 => x"25",
         10636 => x"0a",
         10637 => x"00",
         10638 => x"20",
         10639 => x"74",
         10640 => x"43",
         10641 => x"6b",
         10642 => x"65",
         10643 => x"20",
         10644 => x"20",
         10645 => x"25",
         10646 => x"30",
         10647 => x"48",
         10648 => x"00",
         10649 => x"20",
         10650 => x"41",
         10651 => x"6c",
         10652 => x"20",
         10653 => x"71",
         10654 => x"20",
         10655 => x"20",
         10656 => x"25",
         10657 => x"30",
         10658 => x"48",
         10659 => x"00",
         10660 => x"20",
         10661 => x"68",
         10662 => x"65",
         10663 => x"52",
         10664 => x"43",
         10665 => x"6b",
         10666 => x"65",
         10667 => x"25",
         10668 => x"30",
         10669 => x"48",
         10670 => x"00",
         10671 => x"6c",
         10672 => x"00",
         10673 => x"69",
         10674 => x"00",
         10675 => x"78",
         10676 => x"00",
         10677 => x"00",
         10678 => x"6d",
         10679 => x"00",
         10680 => x"6e",
         10681 => x"00",
         10682 => x"44",
         10683 => x"00",
         10684 => x"02",
         10685 => x"40",
         10686 => x"00",
         10687 => x"03",
         10688 => x"3c",
         10689 => x"00",
         10690 => x"04",
         10691 => x"38",
         10692 => x"00",
         10693 => x"05",
         10694 => x"34",
         10695 => x"00",
         10696 => x"06",
         10697 => x"30",
         10698 => x"00",
         10699 => x"07",
         10700 => x"2c",
         10701 => x"00",
         10702 => x"01",
         10703 => x"28",
         10704 => x"00",
         10705 => x"08",
         10706 => x"24",
         10707 => x"00",
         10708 => x"0b",
         10709 => x"20",
         10710 => x"00",
         10711 => x"09",
         10712 => x"1c",
         10713 => x"00",
         10714 => x"0a",
         10715 => x"18",
         10716 => x"00",
         10717 => x"0d",
         10718 => x"14",
         10719 => x"00",
         10720 => x"0c",
         10721 => x"10",
         10722 => x"00",
         10723 => x"0e",
         10724 => x"0c",
         10725 => x"00",
         10726 => x"0f",
         10727 => x"08",
         10728 => x"00",
         10729 => x"0f",
         10730 => x"04",
         10731 => x"00",
         10732 => x"10",
         10733 => x"00",
         10734 => x"00",
         10735 => x"11",
         10736 => x"fc",
         10737 => x"00",
         10738 => x"12",
         10739 => x"f8",
         10740 => x"00",
         10741 => x"13",
         10742 => x"f4",
         10743 => x"00",
         10744 => x"14",
         10745 => x"f0",
         10746 => x"00",
         10747 => x"15",
         10748 => x"00",
         10749 => x"00",
         10750 => x"00",
         10751 => x"00",
         10752 => x"7e",
         10753 => x"7e",
         10754 => x"7e",
         10755 => x"00",
         10756 => x"7e",
         10757 => x"7e",
         10758 => x"7e",
         10759 => x"00",
         10760 => x"00",
         10761 => x"00",
         10762 => x"00",
         10763 => x"00",
         10764 => x"00",
         10765 => x"00",
         10766 => x"00",
         10767 => x"00",
         10768 => x"00",
         10769 => x"00",
         10770 => x"74",
         10771 => x"00",
         10772 => x"74",
         10773 => x"00",
         10774 => x"00",
         10775 => x"6c",
         10776 => x"25",
         10777 => x"00",
         10778 => x"6c",
         10779 => x"74",
         10780 => x"65",
         10781 => x"20",
         10782 => x"20",
         10783 => x"74",
         10784 => x"20",
         10785 => x"65",
         10786 => x"20",
         10787 => x"2e",
         10788 => x"00",
         10789 => x"6e",
         10790 => x"6f",
         10791 => x"2f",
         10792 => x"61",
         10793 => x"68",
         10794 => x"6f",
         10795 => x"66",
         10796 => x"2c",
         10797 => x"73",
         10798 => x"69",
         10799 => x"00",
         10800 => x"00",
         10801 => x"3c",
         10802 => x"7f",
         10803 => x"00",
         10804 => x"3d",
         10805 => x"00",
         10806 => x"00",
         10807 => x"33",
         10808 => x"00",
         10809 => x"4d",
         10810 => x"53",
         10811 => x"00",
         10812 => x"4e",
         10813 => x"20",
         10814 => x"46",
         10815 => x"32",
         10816 => x"00",
         10817 => x"4e",
         10818 => x"20",
         10819 => x"46",
         10820 => x"20",
         10821 => x"00",
         10822 => x"c0",
         10823 => x"00",
         10824 => x"00",
         10825 => x"00",
         10826 => x"07",
         10827 => x"12",
         10828 => x"1c",
         10829 => x"00",
         10830 => x"41",
         10831 => x"80",
         10832 => x"49",
         10833 => x"8f",
         10834 => x"4f",
         10835 => x"55",
         10836 => x"9b",
         10837 => x"9f",
         10838 => x"55",
         10839 => x"a7",
         10840 => x"ab",
         10841 => x"af",
         10842 => x"b3",
         10843 => x"b7",
         10844 => x"bb",
         10845 => x"bf",
         10846 => x"c3",
         10847 => x"c7",
         10848 => x"cb",
         10849 => x"cf",
         10850 => x"d3",
         10851 => x"d7",
         10852 => x"db",
         10853 => x"df",
         10854 => x"e3",
         10855 => x"e7",
         10856 => x"eb",
         10857 => x"ef",
         10858 => x"f3",
         10859 => x"f7",
         10860 => x"fb",
         10861 => x"ff",
         10862 => x"3b",
         10863 => x"2f",
         10864 => x"3a",
         10865 => x"7c",
         10866 => x"00",
         10867 => x"04",
         10868 => x"40",
         10869 => x"00",
         10870 => x"00",
         10871 => x"02",
         10872 => x"08",
         10873 => x"20",
         10874 => x"00",
         10875 => x"fc",
         10876 => x"e2",
         10877 => x"e0",
         10878 => x"e7",
         10879 => x"eb",
         10880 => x"ef",
         10881 => x"ec",
         10882 => x"c5",
         10883 => x"e6",
         10884 => x"f4",
         10885 => x"f2",
         10886 => x"f9",
         10887 => x"d6",
         10888 => x"a2",
         10889 => x"a5",
         10890 => x"92",
         10891 => x"ed",
         10892 => x"fa",
         10893 => x"d1",
         10894 => x"ba",
         10895 => x"10",
         10896 => x"bd",
         10897 => x"a1",
         10898 => x"bb",
         10899 => x"92",
         10900 => x"02",
         10901 => x"61",
         10902 => x"56",
         10903 => x"63",
         10904 => x"57",
         10905 => x"5c",
         10906 => x"10",
         10907 => x"34",
         10908 => x"1c",
         10909 => x"3c",
         10910 => x"5f",
         10911 => x"54",
         10912 => x"66",
         10913 => x"50",
         10914 => x"67",
         10915 => x"64",
         10916 => x"59",
         10917 => x"52",
         10918 => x"6b",
         10919 => x"18",
         10920 => x"88",
         10921 => x"8c",
         10922 => x"80",
         10923 => x"df",
         10924 => x"c0",
         10925 => x"c3",
         10926 => x"c4",
         10927 => x"98",
         10928 => x"b4",
         10929 => x"c6",
         10930 => x"29",
         10931 => x"b1",
         10932 => x"64",
         10933 => x"21",
         10934 => x"48",
         10935 => x"19",
         10936 => x"1a",
         10937 => x"b2",
         10938 => x"a0",
         10939 => x"1a",
         10940 => x"17",
         10941 => x"07",
         10942 => x"01",
         10943 => x"00",
         10944 => x"32",
         10945 => x"39",
         10946 => x"4a",
         10947 => x"79",
         10948 => x"80",
         10949 => x"43",
         10950 => x"82",
         10951 => x"84",
         10952 => x"86",
         10953 => x"87",
         10954 => x"8a",
         10955 => x"8b",
         10956 => x"8e",
         10957 => x"90",
         10958 => x"91",
         10959 => x"94",
         10960 => x"96",
         10961 => x"98",
         10962 => x"3d",
         10963 => x"9c",
         10964 => x"20",
         10965 => x"a0",
         10966 => x"a2",
         10967 => x"a4",
         10968 => x"a6",
         10969 => x"a7",
         10970 => x"aa",
         10971 => x"ac",
         10972 => x"ae",
         10973 => x"af",
         10974 => x"b2",
         10975 => x"b3",
         10976 => x"b5",
         10977 => x"b8",
         10978 => x"ba",
         10979 => x"bc",
         10980 => x"be",
         10981 => x"c0",
         10982 => x"c2",
         10983 => x"c4",
         10984 => x"c4",
         10985 => x"c8",
         10986 => x"ca",
         10987 => x"ca",
         10988 => x"10",
         10989 => x"01",
         10990 => x"de",
         10991 => x"f3",
         10992 => x"f1",
         10993 => x"f4",
         10994 => x"28",
         10995 => x"12",
         10996 => x"09",
         10997 => x"3b",
         10998 => x"3d",
         10999 => x"3f",
         11000 => x"41",
         11001 => x"46",
         11002 => x"53",
         11003 => x"81",
         11004 => x"55",
         11005 => x"8a",
         11006 => x"8f",
         11007 => x"90",
         11008 => x"5d",
         11009 => x"5f",
         11010 => x"61",
         11011 => x"94",
         11012 => x"65",
         11013 => x"67",
         11014 => x"96",
         11015 => x"62",
         11016 => x"6d",
         11017 => x"9c",
         11018 => x"71",
         11019 => x"73",
         11020 => x"9f",
         11021 => x"77",
         11022 => x"79",
         11023 => x"7b",
         11024 => x"64",
         11025 => x"7f",
         11026 => x"81",
         11027 => x"a9",
         11028 => x"85",
         11029 => x"87",
         11030 => x"44",
         11031 => x"b2",
         11032 => x"8d",
         11033 => x"8f",
         11034 => x"91",
         11035 => x"7b",
         11036 => x"fd",
         11037 => x"ff",
         11038 => x"04",
         11039 => x"88",
         11040 => x"8a",
         11041 => x"11",
         11042 => x"02",
         11043 => x"a3",
         11044 => x"08",
         11045 => x"03",
         11046 => x"8e",
         11047 => x"d8",
         11048 => x"f2",
         11049 => x"f9",
         11050 => x"f4",
         11051 => x"f6",
         11052 => x"f7",
         11053 => x"fa",
         11054 => x"30",
         11055 => x"50",
         11056 => x"60",
         11057 => x"8a",
         11058 => x"c1",
         11059 => x"cf",
         11060 => x"c0",
         11061 => x"44",
         11062 => x"26",
         11063 => x"00",
         11064 => x"01",
         11065 => x"00",
         11066 => x"a0",
         11067 => x"00",
         11068 => x"10",
         11069 => x"20",
         11070 => x"30",
         11071 => x"40",
         11072 => x"51",
         11073 => x"59",
         11074 => x"5b",
         11075 => x"5d",
         11076 => x"5f",
         11077 => x"08",
         11078 => x"0e",
         11079 => x"bb",
         11080 => x"c9",
         11081 => x"cb",
         11082 => x"db",
         11083 => x"f9",
         11084 => x"eb",
         11085 => x"fb",
         11086 => x"08",
         11087 => x"08",
         11088 => x"08",
         11089 => x"04",
         11090 => x"b9",
         11091 => x"bc",
         11092 => x"01",
         11093 => x"d0",
         11094 => x"e0",
         11095 => x"e5",
         11096 => x"ec",
         11097 => x"01",
         11098 => x"4e",
         11099 => x"32",
         11100 => x"10",
         11101 => x"01",
         11102 => x"d0",
         11103 => x"30",
         11104 => x"60",
         11105 => x"67",
         11106 => x"75",
         11107 => x"80",
         11108 => x"00",
         11109 => x"41",
         11110 => x"00",
         11111 => x"00",
         11112 => x"40",
         11113 => x"00",
         11114 => x"00",
         11115 => x"00",
         11116 => x"48",
         11117 => x"00",
         11118 => x"00",
         11119 => x"00",
         11120 => x"50",
         11121 => x"00",
         11122 => x"00",
         11123 => x"00",
         11124 => x"58",
         11125 => x"00",
         11126 => x"00",
         11127 => x"00",
         11128 => x"60",
         11129 => x"00",
         11130 => x"00",
         11131 => x"00",
         11132 => x"68",
         11133 => x"00",
         11134 => x"00",
         11135 => x"00",
         11136 => x"70",
         11137 => x"00",
         11138 => x"00",
         11139 => x"00",
         11140 => x"78",
         11141 => x"00",
         11142 => x"00",
         11143 => x"00",
         11144 => x"80",
         11145 => x"00",
         11146 => x"00",
         11147 => x"00",
         11148 => x"88",
         11149 => x"00",
         11150 => x"00",
         11151 => x"00",
         11152 => x"8c",
         11153 => x"00",
         11154 => x"00",
         11155 => x"00",
         11156 => x"90",
         11157 => x"00",
         11158 => x"00",
         11159 => x"00",
         11160 => x"94",
         11161 => x"00",
         11162 => x"00",
         11163 => x"00",
         11164 => x"98",
         11165 => x"00",
         11166 => x"00",
         11167 => x"00",
         11168 => x"9c",
         11169 => x"00",
         11170 => x"00",
         11171 => x"00",
         11172 => x"a0",
         11173 => x"00",
         11174 => x"00",
         11175 => x"00",
         11176 => x"a4",
         11177 => x"00",
         11178 => x"00",
         11179 => x"00",
         11180 => x"ac",
         11181 => x"00",
         11182 => x"00",
         11183 => x"00",
         11184 => x"b0",
         11185 => x"00",
         11186 => x"00",
         11187 => x"00",
         11188 => x"b8",
         11189 => x"00",
         11190 => x"00",
         11191 => x"00",
         11192 => x"c0",
         11193 => x"00",
         11194 => x"00",
         11195 => x"00",
         11196 => x"c8",
         11197 => x"00",
         11198 => x"00",
         11199 => x"00",
         11200 => x"d0",
         11201 => x"00",
         11202 => x"00",
         11203 => x"00",
         11204 => x"d8",
         11205 => x"00",
         11206 => x"00",
         11207 => x"00",
         11208 => x"e0",
         11209 => x"00",
         11210 => x"00",
         11211 => x"00",
         11212 => x"00",
         11213 => x"00",
         11214 => x"ff",
         11215 => x"00",
         11216 => x"ff",
         11217 => x"00",
         11218 => x"ff",
         11219 => x"00",
         11220 => x"00",
         11221 => x"00",
         11222 => x"ff",
         11223 => x"00",
         11224 => x"00",
         11225 => x"00",
         11226 => x"00",
         11227 => x"00",
         11228 => x"00",
         11229 => x"00",
         11230 => x"00",
         11231 => x"01",
         11232 => x"01",
         11233 => x"01",
         11234 => x"00",
         11235 => x"00",
         11236 => x"00",
         11237 => x"00",
         11238 => x"00",
         11239 => x"00",
         11240 => x"00",
         11241 => x"00",
         11242 => x"00",
         11243 => x"00",
         11244 => x"00",
         11245 => x"00",
         11246 => x"00",
         11247 => x"00",
         11248 => x"00",
         11249 => x"00",
         11250 => x"00",
         11251 => x"00",
         11252 => x"00",
         11253 => x"00",
         11254 => x"00",
         11255 => x"00",
         11256 => x"00",
         11257 => x"00",
         11258 => x"00",
         11259 => x"48",
         11260 => x"00",
         11261 => x"50",
         11262 => x"00",
         11263 => x"58",
         11264 => x"00",
         11265 => x"00",
         11266 => x"00",
         11267 => x"02",
         11268 => x"04",
         11269 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"0b",
             2 => x"ed",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"88",
            10 => x"90",
            11 => x"88",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"93",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"82",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"80",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"80",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"06",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"0b",
           266 => x"85",
           267 => x"0b",
           268 => x"0b",
           269 => x"a6",
           270 => x"0b",
           271 => x"0b",
           272 => x"c6",
           273 => x"0b",
           274 => x"0b",
           275 => x"e6",
           276 => x"0b",
           277 => x"0b",
           278 => x"88",
           279 => x"0b",
           280 => x"0b",
           281 => x"a8",
           282 => x"0b",
           283 => x"0b",
           284 => x"c9",
           285 => x"0b",
           286 => x"0b",
           287 => x"eb",
           288 => x"0b",
           289 => x"0b",
           290 => x"8d",
           291 => x"0b",
           292 => x"0b",
           293 => x"af",
           294 => x"0b",
           295 => x"0b",
           296 => x"d1",
           297 => x"0b",
           298 => x"0b",
           299 => x"f3",
           300 => x"0b",
           301 => x"0b",
           302 => x"95",
           303 => x"0b",
           304 => x"0b",
           305 => x"b7",
           306 => x"0b",
           307 => x"0b",
           308 => x"d9",
           309 => x"0b",
           310 => x"0b",
           311 => x"fb",
           312 => x"0b",
           313 => x"0b",
           314 => x"9d",
           315 => x"0b",
           316 => x"0b",
           317 => x"bf",
           318 => x"0b",
           319 => x"0b",
           320 => x"e1",
           321 => x"0b",
           322 => x"0b",
           323 => x"83",
           324 => x"0b",
           325 => x"0b",
           326 => x"a5",
           327 => x"0b",
           328 => x"0b",
           329 => x"c7",
           330 => x"0b",
           331 => x"0b",
           332 => x"e9",
           333 => x"0b",
           334 => x"0b",
           335 => x"8b",
           336 => x"0b",
           337 => x"0b",
           338 => x"ad",
           339 => x"0b",
           340 => x"0b",
           341 => x"cf",
           342 => x"0b",
           343 => x"0b",
           344 => x"f1",
           345 => x"0b",
           346 => x"ff",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"8c",
           385 => x"e0",
           386 => x"81",
           387 => x"e0",
           388 => x"c0",
           389 => x"82",
           390 => x"b3",
           391 => x"e0",
           392 => x"c0",
           393 => x"82",
           394 => x"b0",
           395 => x"e0",
           396 => x"c0",
           397 => x"82",
           398 => x"af",
           399 => x"e0",
           400 => x"c0",
           401 => x"82",
           402 => x"94",
           403 => x"e0",
           404 => x"c0",
           405 => x"82",
           406 => x"b1",
           407 => x"e0",
           408 => x"c0",
           409 => x"82",
           410 => x"80",
           411 => x"82",
           412 => x"80",
           413 => x"04",
           414 => x"0c",
           415 => x"2d",
           416 => x"08",
           417 => x"90",
           418 => x"a4",
           419 => x"2d",
           420 => x"08",
           421 => x"90",
           422 => x"a4",
           423 => x"2d",
           424 => x"08",
           425 => x"90",
           426 => x"a4",
           427 => x"2d",
           428 => x"08",
           429 => x"90",
           430 => x"a4",
           431 => x"e7",
           432 => x"a4",
           433 => x"80",
           434 => x"e0",
           435 => x"ff",
           436 => x"e0",
           437 => x"c0",
           438 => x"82",
           439 => x"81",
           440 => x"82",
           441 => x"80",
           442 => x"04",
           443 => x"0c",
           444 => x"2d",
           445 => x"08",
           446 => x"90",
           447 => x"a4",
           448 => x"e5",
           449 => x"a4",
           450 => x"80",
           451 => x"e0",
           452 => x"f6",
           453 => x"e0",
           454 => x"c0",
           455 => x"82",
           456 => x"82",
           457 => x"82",
           458 => x"80",
           459 => x"04",
           460 => x"0c",
           461 => x"2d",
           462 => x"08",
           463 => x"90",
           464 => x"a4",
           465 => x"8c",
           466 => x"a4",
           467 => x"80",
           468 => x"e0",
           469 => x"88",
           470 => x"e0",
           471 => x"c0",
           472 => x"82",
           473 => x"82",
           474 => x"82",
           475 => x"80",
           476 => x"04",
           477 => x"0c",
           478 => x"2d",
           479 => x"08",
           480 => x"90",
           481 => x"a4",
           482 => x"88",
           483 => x"a4",
           484 => x"80",
           485 => x"e0",
           486 => x"8d",
           487 => x"e0",
           488 => x"c0",
           489 => x"82",
           490 => x"82",
           491 => x"82",
           492 => x"80",
           493 => x"04",
           494 => x"0c",
           495 => x"2d",
           496 => x"08",
           497 => x"90",
           498 => x"a4",
           499 => x"9d",
           500 => x"a4",
           501 => x"80",
           502 => x"e0",
           503 => x"98",
           504 => x"e0",
           505 => x"c0",
           506 => x"82",
           507 => x"82",
           508 => x"82",
           509 => x"80",
           510 => x"04",
           511 => x"0c",
           512 => x"2d",
           513 => x"08",
           514 => x"90",
           515 => x"a4",
           516 => x"9d",
           517 => x"a4",
           518 => x"80",
           519 => x"e0",
           520 => x"84",
           521 => x"e0",
           522 => x"c0",
           523 => x"82",
           524 => x"82",
           525 => x"82",
           526 => x"80",
           527 => x"04",
           528 => x"0c",
           529 => x"2d",
           530 => x"08",
           531 => x"90",
           532 => x"a4",
           533 => x"a4",
           534 => x"a4",
           535 => x"80",
           536 => x"e0",
           537 => x"9d",
           538 => x"e0",
           539 => x"c0",
           540 => x"82",
           541 => x"82",
           542 => x"82",
           543 => x"80",
           544 => x"04",
           545 => x"0c",
           546 => x"2d",
           547 => x"08",
           548 => x"90",
           549 => x"a4",
           550 => x"c6",
           551 => x"a4",
           552 => x"80",
           553 => x"e0",
           554 => x"a5",
           555 => x"e0",
           556 => x"c0",
           557 => x"82",
           558 => x"82",
           559 => x"82",
           560 => x"80",
           561 => x"04",
           562 => x"0c",
           563 => x"2d",
           564 => x"08",
           565 => x"90",
           566 => x"a4",
           567 => x"8b",
           568 => x"a4",
           569 => x"80",
           570 => x"e0",
           571 => x"b6",
           572 => x"e0",
           573 => x"c0",
           574 => x"82",
           575 => x"81",
           576 => x"82",
           577 => x"80",
           578 => x"04",
           579 => x"0c",
           580 => x"2d",
           581 => x"08",
           582 => x"90",
           583 => x"a4",
           584 => x"88",
           585 => x"a4",
           586 => x"80",
           587 => x"e0",
           588 => x"82",
           589 => x"e0",
           590 => x"c0",
           591 => x"82",
           592 => x"80",
           593 => x"82",
           594 => x"80",
           595 => x"04",
           596 => x"0c",
           597 => x"2d",
           598 => x"08",
           599 => x"90",
           600 => x"a4",
           601 => x"c7",
           602 => x"a4",
           603 => x"80",
           604 => x"e0",
           605 => x"b3",
           606 => x"e0",
           607 => x"c0",
           608 => x"82",
           609 => x"81",
           610 => x"82",
           611 => x"80",
           612 => x"04",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"10",
           621 => x"04",
           622 => x"81",
           623 => x"83",
           624 => x"05",
           625 => x"10",
           626 => x"72",
           627 => x"51",
           628 => x"72",
           629 => x"06",
           630 => x"72",
           631 => x"10",
           632 => x"10",
           633 => x"ed",
           634 => x"53",
           635 => x"e0",
           636 => x"fc",
           637 => x"38",
           638 => x"84",
           639 => x"0b",
           640 => x"f0",
           641 => x"51",
           642 => x"04",
           643 => x"a4",
           644 => x"e0",
           645 => x"3d",
           646 => x"a4",
           647 => x"70",
           648 => x"08",
           649 => x"82",
           650 => x"fc",
           651 => x"82",
           652 => x"88",
           653 => x"82",
           654 => x"52",
           655 => x"3f",
           656 => x"08",
           657 => x"a4",
           658 => x"0c",
           659 => x"08",
           660 => x"70",
           661 => x"0c",
           662 => x"3d",
           663 => x"a4",
           664 => x"e0",
           665 => x"82",
           666 => x"fb",
           667 => x"e0",
           668 => x"05",
           669 => x"33",
           670 => x"70",
           671 => x"51",
           672 => x"8f",
           673 => x"82",
           674 => x"8c",
           675 => x"83",
           676 => x"80",
           677 => x"a4",
           678 => x"0c",
           679 => x"82",
           680 => x"8c",
           681 => x"05",
           682 => x"08",
           683 => x"80",
           684 => x"a4",
           685 => x"0c",
           686 => x"08",
           687 => x"82",
           688 => x"fc",
           689 => x"e0",
           690 => x"05",
           691 => x"80",
           692 => x"0b",
           693 => x"08",
           694 => x"25",
           695 => x"82",
           696 => x"90",
           697 => x"a0",
           698 => x"e0",
           699 => x"82",
           700 => x"f8",
           701 => x"82",
           702 => x"f8",
           703 => x"2e",
           704 => x"8d",
           705 => x"82",
           706 => x"f4",
           707 => x"d2",
           708 => x"a4",
           709 => x"08",
           710 => x"08",
           711 => x"53",
           712 => x"34",
           713 => x"08",
           714 => x"ff",
           715 => x"a4",
           716 => x"0c",
           717 => x"08",
           718 => x"81",
           719 => x"a4",
           720 => x"0c",
           721 => x"82",
           722 => x"fc",
           723 => x"80",
           724 => x"e0",
           725 => x"05",
           726 => x"e0",
           727 => x"05",
           728 => x"e0",
           729 => x"05",
           730 => x"98",
           731 => x"0d",
           732 => x"0c",
           733 => x"a4",
           734 => x"e0",
           735 => x"3d",
           736 => x"82",
           737 => x"e5",
           738 => x"e0",
           739 => x"05",
           740 => x"a4",
           741 => x"0c",
           742 => x"82",
           743 => x"e8",
           744 => x"e0",
           745 => x"05",
           746 => x"a4",
           747 => x"0c",
           748 => x"08",
           749 => x"54",
           750 => x"08",
           751 => x"53",
           752 => x"08",
           753 => x"53",
           754 => x"8d",
           755 => x"98",
           756 => x"e0",
           757 => x"05",
           758 => x"a4",
           759 => x"08",
           760 => x"08",
           761 => x"05",
           762 => x"74",
           763 => x"a4",
           764 => x"08",
           765 => x"98",
           766 => x"3d",
           767 => x"a4",
           768 => x"e0",
           769 => x"82",
           770 => x"fb",
           771 => x"e0",
           772 => x"05",
           773 => x"a4",
           774 => x"0c",
           775 => x"08",
           776 => x"54",
           777 => x"08",
           778 => x"53",
           779 => x"08",
           780 => x"52",
           781 => x"82",
           782 => x"70",
           783 => x"08",
           784 => x"82",
           785 => x"f8",
           786 => x"82",
           787 => x"51",
           788 => x"0d",
           789 => x"0c",
           790 => x"a4",
           791 => x"e0",
           792 => x"3d",
           793 => x"82",
           794 => x"e4",
           795 => x"e0",
           796 => x"05",
           797 => x"0b",
           798 => x"82",
           799 => x"88",
           800 => x"11",
           801 => x"2a",
           802 => x"70",
           803 => x"51",
           804 => x"72",
           805 => x"38",
           806 => x"e0",
           807 => x"05",
           808 => x"39",
           809 => x"08",
           810 => x"53",
           811 => x"72",
           812 => x"08",
           813 => x"72",
           814 => x"53",
           815 => x"95",
           816 => x"e0",
           817 => x"05",
           818 => x"82",
           819 => x"8c",
           820 => x"e0",
           821 => x"05",
           822 => x"06",
           823 => x"80",
           824 => x"38",
           825 => x"08",
           826 => x"53",
           827 => x"81",
           828 => x"e0",
           829 => x"05",
           830 => x"b9",
           831 => x"38",
           832 => x"08",
           833 => x"53",
           834 => x"09",
           835 => x"c5",
           836 => x"a4",
           837 => x"33",
           838 => x"70",
           839 => x"51",
           840 => x"38",
           841 => x"08",
           842 => x"70",
           843 => x"81",
           844 => x"06",
           845 => x"53",
           846 => x"99",
           847 => x"a4",
           848 => x"22",
           849 => x"07",
           850 => x"82",
           851 => x"e4",
           852 => x"d0",
           853 => x"a4",
           854 => x"33",
           855 => x"70",
           856 => x"70",
           857 => x"11",
           858 => x"51",
           859 => x"55",
           860 => x"e0",
           861 => x"05",
           862 => x"a4",
           863 => x"33",
           864 => x"a4",
           865 => x"33",
           866 => x"11",
           867 => x"72",
           868 => x"08",
           869 => x"82",
           870 => x"e8",
           871 => x"98",
           872 => x"2c",
           873 => x"72",
           874 => x"38",
           875 => x"82",
           876 => x"e8",
           877 => x"e0",
           878 => x"05",
           879 => x"2a",
           880 => x"51",
           881 => x"fd",
           882 => x"e0",
           883 => x"05",
           884 => x"2b",
           885 => x"70",
           886 => x"88",
           887 => x"51",
           888 => x"82",
           889 => x"ec",
           890 => x"b8",
           891 => x"a4",
           892 => x"22",
           893 => x"70",
           894 => x"51",
           895 => x"2e",
           896 => x"e0",
           897 => x"05",
           898 => x"2b",
           899 => x"51",
           900 => x"8a",
           901 => x"82",
           902 => x"e8",
           903 => x"e0",
           904 => x"05",
           905 => x"82",
           906 => x"c4",
           907 => x"82",
           908 => x"c4",
           909 => x"d8",
           910 => x"38",
           911 => x"08",
           912 => x"70",
           913 => x"b9",
           914 => x"08",
           915 => x"53",
           916 => x"e0",
           917 => x"05",
           918 => x"07",
           919 => x"82",
           920 => x"e4",
           921 => x"e0",
           922 => x"05",
           923 => x"07",
           924 => x"82",
           925 => x"e4",
           926 => x"a8",
           927 => x"a4",
           928 => x"22",
           929 => x"07",
           930 => x"82",
           931 => x"e4",
           932 => x"90",
           933 => x"a4",
           934 => x"22",
           935 => x"07",
           936 => x"82",
           937 => x"e4",
           938 => x"f8",
           939 => x"a4",
           940 => x"22",
           941 => x"51",
           942 => x"e0",
           943 => x"05",
           944 => x"82",
           945 => x"e8",
           946 => x"d8",
           947 => x"a4",
           948 => x"22",
           949 => x"51",
           950 => x"e0",
           951 => x"05",
           952 => x"39",
           953 => x"e0",
           954 => x"05",
           955 => x"a4",
           956 => x"22",
           957 => x"53",
           958 => x"a4",
           959 => x"23",
           960 => x"82",
           961 => x"f8",
           962 => x"a8",
           963 => x"a4",
           964 => x"08",
           965 => x"08",
           966 => x"84",
           967 => x"a4",
           968 => x"0c",
           969 => x"53",
           970 => x"a4",
           971 => x"34",
           972 => x"08",
           973 => x"ff",
           974 => x"72",
           975 => x"08",
           976 => x"8c",
           977 => x"e0",
           978 => x"05",
           979 => x"a4",
           980 => x"08",
           981 => x"e0",
           982 => x"05",
           983 => x"82",
           984 => x"fc",
           985 => x"e0",
           986 => x"05",
           987 => x"2a",
           988 => x"51",
           989 => x"72",
           990 => x"38",
           991 => x"08",
           992 => x"70",
           993 => x"72",
           994 => x"82",
           995 => x"fc",
           996 => x"53",
           997 => x"82",
           998 => x"53",
           999 => x"a4",
          1000 => x"23",
          1001 => x"e0",
          1002 => x"05",
          1003 => x"8a",
          1004 => x"98",
          1005 => x"82",
          1006 => x"f4",
          1007 => x"e0",
          1008 => x"05",
          1009 => x"e0",
          1010 => x"05",
          1011 => x"31",
          1012 => x"82",
          1013 => x"ec",
          1014 => x"d8",
          1015 => x"a4",
          1016 => x"08",
          1017 => x"08",
          1018 => x"84",
          1019 => x"a4",
          1020 => x"0c",
          1021 => x"e0",
          1022 => x"05",
          1023 => x"a4",
          1024 => x"22",
          1025 => x"70",
          1026 => x"51",
          1027 => x"80",
          1028 => x"82",
          1029 => x"e8",
          1030 => x"98",
          1031 => x"98",
          1032 => x"e0",
          1033 => x"05",
          1034 => x"a2",
          1035 => x"e0",
          1036 => x"72",
          1037 => x"08",
          1038 => x"99",
          1039 => x"a4",
          1040 => x"08",
          1041 => x"3f",
          1042 => x"08",
          1043 => x"e0",
          1044 => x"05",
          1045 => x"a4",
          1046 => x"22",
          1047 => x"a4",
          1048 => x"22",
          1049 => x"54",
          1050 => x"e0",
          1051 => x"05",
          1052 => x"39",
          1053 => x"08",
          1054 => x"70",
          1055 => x"81",
          1056 => x"53",
          1057 => x"a4",
          1058 => x"a4",
          1059 => x"08",
          1060 => x"08",
          1061 => x"84",
          1062 => x"a4",
          1063 => x"0c",
          1064 => x"e0",
          1065 => x"05",
          1066 => x"39",
          1067 => x"08",
          1068 => x"82",
          1069 => x"90",
          1070 => x"05",
          1071 => x"08",
          1072 => x"70",
          1073 => x"a4",
          1074 => x"0c",
          1075 => x"a4",
          1076 => x"08",
          1077 => x"08",
          1078 => x"82",
          1079 => x"fc",
          1080 => x"25",
          1081 => x"e0",
          1082 => x"05",
          1083 => x"07",
          1084 => x"82",
          1085 => x"e4",
          1086 => x"e0",
          1087 => x"05",
          1088 => x"e0",
          1089 => x"05",
          1090 => x"a4",
          1091 => x"22",
          1092 => x"06",
          1093 => x"82",
          1094 => x"e4",
          1095 => x"af",
          1096 => x"82",
          1097 => x"f4",
          1098 => x"39",
          1099 => x"08",
          1100 => x"70",
          1101 => x"51",
          1102 => x"e0",
          1103 => x"05",
          1104 => x"0b",
          1105 => x"08",
          1106 => x"90",
          1107 => x"a4",
          1108 => x"23",
          1109 => x"08",
          1110 => x"70",
          1111 => x"81",
          1112 => x"53",
          1113 => x"a4",
          1114 => x"a4",
          1115 => x"08",
          1116 => x"08",
          1117 => x"84",
          1118 => x"a4",
          1119 => x"0c",
          1120 => x"e0",
          1121 => x"05",
          1122 => x"39",
          1123 => x"08",
          1124 => x"82",
          1125 => x"90",
          1126 => x"05",
          1127 => x"08",
          1128 => x"70",
          1129 => x"a4",
          1130 => x"0c",
          1131 => x"a4",
          1132 => x"08",
          1133 => x"08",
          1134 => x"82",
          1135 => x"e4",
          1136 => x"cf",
          1137 => x"72",
          1138 => x"08",
          1139 => x"82",
          1140 => x"82",
          1141 => x"f0",
          1142 => x"e0",
          1143 => x"05",
          1144 => x"a4",
          1145 => x"22",
          1146 => x"08",
          1147 => x"71",
          1148 => x"56",
          1149 => x"ca",
          1150 => x"98",
          1151 => x"75",
          1152 => x"a4",
          1153 => x"08",
          1154 => x"08",
          1155 => x"82",
          1156 => x"f0",
          1157 => x"33",
          1158 => x"73",
          1159 => x"82",
          1160 => x"f0",
          1161 => x"72",
          1162 => x"e0",
          1163 => x"05",
          1164 => x"df",
          1165 => x"53",
          1166 => x"a4",
          1167 => x"34",
          1168 => x"e0",
          1169 => x"05",
          1170 => x"33",
          1171 => x"53",
          1172 => x"a4",
          1173 => x"34",
          1174 => x"08",
          1175 => x"53",
          1176 => x"08",
          1177 => x"73",
          1178 => x"a4",
          1179 => x"08",
          1180 => x"e0",
          1181 => x"05",
          1182 => x"a4",
          1183 => x"22",
          1184 => x"e0",
          1185 => x"05",
          1186 => x"a0",
          1187 => x"e0",
          1188 => x"82",
          1189 => x"fc",
          1190 => x"82",
          1191 => x"fc",
          1192 => x"2e",
          1193 => x"b2",
          1194 => x"a4",
          1195 => x"08",
          1196 => x"54",
          1197 => x"74",
          1198 => x"51",
          1199 => x"e0",
          1200 => x"05",
          1201 => x"a4",
          1202 => x"22",
          1203 => x"51",
          1204 => x"2e",
          1205 => x"e0",
          1206 => x"05",
          1207 => x"51",
          1208 => x"e0",
          1209 => x"05",
          1210 => x"a4",
          1211 => x"22",
          1212 => x"70",
          1213 => x"51",
          1214 => x"2e",
          1215 => x"82",
          1216 => x"ec",
          1217 => x"90",
          1218 => x"a4",
          1219 => x"0c",
          1220 => x"08",
          1221 => x"90",
          1222 => x"a4",
          1223 => x"0c",
          1224 => x"08",
          1225 => x"51",
          1226 => x"2e",
          1227 => x"95",
          1228 => x"a4",
          1229 => x"08",
          1230 => x"72",
          1231 => x"08",
          1232 => x"93",
          1233 => x"a4",
          1234 => x"08",
          1235 => x"72",
          1236 => x"08",
          1237 => x"82",
          1238 => x"c8",
          1239 => x"e0",
          1240 => x"05",
          1241 => x"a4",
          1242 => x"22",
          1243 => x"70",
          1244 => x"51",
          1245 => x"2e",
          1246 => x"82",
          1247 => x"e8",
          1248 => x"98",
          1249 => x"2c",
          1250 => x"08",
          1251 => x"57",
          1252 => x"72",
          1253 => x"38",
          1254 => x"08",
          1255 => x"70",
          1256 => x"53",
          1257 => x"a4",
          1258 => x"23",
          1259 => x"e0",
          1260 => x"05",
          1261 => x"e0",
          1262 => x"05",
          1263 => x"31",
          1264 => x"82",
          1265 => x"e8",
          1266 => x"e0",
          1267 => x"05",
          1268 => x"2a",
          1269 => x"51",
          1270 => x"80",
          1271 => x"82",
          1272 => x"e8",
          1273 => x"88",
          1274 => x"2b",
          1275 => x"70",
          1276 => x"51",
          1277 => x"72",
          1278 => x"a4",
          1279 => x"22",
          1280 => x"51",
          1281 => x"e0",
          1282 => x"05",
          1283 => x"82",
          1284 => x"fc",
          1285 => x"88",
          1286 => x"2b",
          1287 => x"70",
          1288 => x"51",
          1289 => x"72",
          1290 => x"a4",
          1291 => x"22",
          1292 => x"51",
          1293 => x"e0",
          1294 => x"05",
          1295 => x"a4",
          1296 => x"22",
          1297 => x"06",
          1298 => x"b0",
          1299 => x"a4",
          1300 => x"22",
          1301 => x"54",
          1302 => x"a4",
          1303 => x"23",
          1304 => x"70",
          1305 => x"53",
          1306 => x"90",
          1307 => x"a4",
          1308 => x"08",
          1309 => x"8a",
          1310 => x"39",
          1311 => x"08",
          1312 => x"70",
          1313 => x"81",
          1314 => x"53",
          1315 => x"91",
          1316 => x"a4",
          1317 => x"08",
          1318 => x"8a",
          1319 => x"c7",
          1320 => x"a4",
          1321 => x"22",
          1322 => x"70",
          1323 => x"51",
          1324 => x"2e",
          1325 => x"e0",
          1326 => x"05",
          1327 => x"51",
          1328 => x"a3",
          1329 => x"a4",
          1330 => x"22",
          1331 => x"70",
          1332 => x"51",
          1333 => x"2e",
          1334 => x"e0",
          1335 => x"05",
          1336 => x"51",
          1337 => x"82",
          1338 => x"e4",
          1339 => x"86",
          1340 => x"06",
          1341 => x"72",
          1342 => x"38",
          1343 => x"08",
          1344 => x"52",
          1345 => x"df",
          1346 => x"a4",
          1347 => x"22",
          1348 => x"2e",
          1349 => x"94",
          1350 => x"a4",
          1351 => x"08",
          1352 => x"a4",
          1353 => x"33",
          1354 => x"3f",
          1355 => x"08",
          1356 => x"70",
          1357 => x"81",
          1358 => x"53",
          1359 => x"b0",
          1360 => x"a4",
          1361 => x"22",
          1362 => x"54",
          1363 => x"a4",
          1364 => x"23",
          1365 => x"70",
          1366 => x"53",
          1367 => x"90",
          1368 => x"a4",
          1369 => x"08",
          1370 => x"88",
          1371 => x"39",
          1372 => x"08",
          1373 => x"70",
          1374 => x"81",
          1375 => x"53",
          1376 => x"b0",
          1377 => x"a4",
          1378 => x"33",
          1379 => x"54",
          1380 => x"a4",
          1381 => x"34",
          1382 => x"70",
          1383 => x"53",
          1384 => x"90",
          1385 => x"a4",
          1386 => x"08",
          1387 => x"88",
          1388 => x"39",
          1389 => x"08",
          1390 => x"70",
          1391 => x"81",
          1392 => x"53",
          1393 => x"82",
          1394 => x"ec",
          1395 => x"11",
          1396 => x"82",
          1397 => x"ec",
          1398 => x"90",
          1399 => x"2c",
          1400 => x"73",
          1401 => x"82",
          1402 => x"88",
          1403 => x"a0",
          1404 => x"3f",
          1405 => x"e0",
          1406 => x"05",
          1407 => x"80",
          1408 => x"81",
          1409 => x"82",
          1410 => x"88",
          1411 => x"82",
          1412 => x"fc",
          1413 => x"87",
          1414 => x"ee",
          1415 => x"a4",
          1416 => x"33",
          1417 => x"f3",
          1418 => x"06",
          1419 => x"82",
          1420 => x"f4",
          1421 => x"11",
          1422 => x"82",
          1423 => x"f4",
          1424 => x"83",
          1425 => x"53",
          1426 => x"ff",
          1427 => x"38",
          1428 => x"08",
          1429 => x"52",
          1430 => x"08",
          1431 => x"70",
          1432 => x"e0",
          1433 => x"05",
          1434 => x"82",
          1435 => x"fc",
          1436 => x"86",
          1437 => x"b7",
          1438 => x"a4",
          1439 => x"33",
          1440 => x"d3",
          1441 => x"06",
          1442 => x"82",
          1443 => x"f4",
          1444 => x"11",
          1445 => x"82",
          1446 => x"f4",
          1447 => x"83",
          1448 => x"53",
          1449 => x"ff",
          1450 => x"38",
          1451 => x"08",
          1452 => x"52",
          1453 => x"08",
          1454 => x"70",
          1455 => x"86",
          1456 => x"e0",
          1457 => x"05",
          1458 => x"82",
          1459 => x"fc",
          1460 => x"b7",
          1461 => x"a4",
          1462 => x"08",
          1463 => x"2e",
          1464 => x"e0",
          1465 => x"05",
          1466 => x"e0",
          1467 => x"05",
          1468 => x"82",
          1469 => x"f0",
          1470 => x"e0",
          1471 => x"05",
          1472 => x"52",
          1473 => x"3f",
          1474 => x"e0",
          1475 => x"05",
          1476 => x"2a",
          1477 => x"51",
          1478 => x"80",
          1479 => x"38",
          1480 => x"08",
          1481 => x"ff",
          1482 => x"72",
          1483 => x"08",
          1484 => x"73",
          1485 => x"90",
          1486 => x"80",
          1487 => x"38",
          1488 => x"08",
          1489 => x"52",
          1490 => x"9b",
          1491 => x"82",
          1492 => x"88",
          1493 => x"82",
          1494 => x"f8",
          1495 => x"85",
          1496 => x"0b",
          1497 => x"08",
          1498 => x"ea",
          1499 => x"e0",
          1500 => x"05",
          1501 => x"a5",
          1502 => x"06",
          1503 => x"0b",
          1504 => x"08",
          1505 => x"80",
          1506 => x"a4",
          1507 => x"23",
          1508 => x"e0",
          1509 => x"05",
          1510 => x"82",
          1511 => x"f4",
          1512 => x"80",
          1513 => x"a4",
          1514 => x"08",
          1515 => x"a4",
          1516 => x"33",
          1517 => x"3f",
          1518 => x"82",
          1519 => x"88",
          1520 => x"11",
          1521 => x"e0",
          1522 => x"05",
          1523 => x"82",
          1524 => x"e0",
          1525 => x"e0",
          1526 => x"3d",
          1527 => x"a4",
          1528 => x"e0",
          1529 => x"82",
          1530 => x"fd",
          1531 => x"fb",
          1532 => x"82",
          1533 => x"8c",
          1534 => x"82",
          1535 => x"88",
          1536 => x"e4",
          1537 => x"e0",
          1538 => x"82",
          1539 => x"54",
          1540 => x"82",
          1541 => x"04",
          1542 => x"08",
          1543 => x"a4",
          1544 => x"0d",
          1545 => x"e0",
          1546 => x"05",
          1547 => x"fc",
          1548 => x"33",
          1549 => x"70",
          1550 => x"81",
          1551 => x"51",
          1552 => x"80",
          1553 => x"ff",
          1554 => x"a4",
          1555 => x"0c",
          1556 => x"82",
          1557 => x"88",
          1558 => x"72",
          1559 => x"a4",
          1560 => x"08",
          1561 => x"e0",
          1562 => x"05",
          1563 => x"82",
          1564 => x"fc",
          1565 => x"81",
          1566 => x"72",
          1567 => x"38",
          1568 => x"08",
          1569 => x"08",
          1570 => x"a4",
          1571 => x"33",
          1572 => x"08",
          1573 => x"2d",
          1574 => x"08",
          1575 => x"2e",
          1576 => x"ff",
          1577 => x"a4",
          1578 => x"0c",
          1579 => x"82",
          1580 => x"82",
          1581 => x"53",
          1582 => x"90",
          1583 => x"72",
          1584 => x"98",
          1585 => x"80",
          1586 => x"ff",
          1587 => x"a4",
          1588 => x"0c",
          1589 => x"08",
          1590 => x"70",
          1591 => x"08",
          1592 => x"53",
          1593 => x"08",
          1594 => x"82",
          1595 => x"87",
          1596 => x"e0",
          1597 => x"82",
          1598 => x"02",
          1599 => x"0c",
          1600 => x"80",
          1601 => x"a4",
          1602 => x"0c",
          1603 => x"08",
          1604 => x"85",
          1605 => x"81",
          1606 => x"32",
          1607 => x"51",
          1608 => x"53",
          1609 => x"8d",
          1610 => x"82",
          1611 => x"f4",
          1612 => x"f3",
          1613 => x"a4",
          1614 => x"08",
          1615 => x"82",
          1616 => x"88",
          1617 => x"05",
          1618 => x"08",
          1619 => x"53",
          1620 => x"a4",
          1621 => x"34",
          1622 => x"06",
          1623 => x"2e",
          1624 => x"e0",
          1625 => x"05",
          1626 => x"a4",
          1627 => x"08",
          1628 => x"a4",
          1629 => x"33",
          1630 => x"08",
          1631 => x"2d",
          1632 => x"08",
          1633 => x"2e",
          1634 => x"ff",
          1635 => x"a4",
          1636 => x"0c",
          1637 => x"82",
          1638 => x"f8",
          1639 => x"82",
          1640 => x"f4",
          1641 => x"82",
          1642 => x"f4",
          1643 => x"e0",
          1644 => x"3d",
          1645 => x"a4",
          1646 => x"e0",
          1647 => x"82",
          1648 => x"fe",
          1649 => x"fb",
          1650 => x"82",
          1651 => x"88",
          1652 => x"93",
          1653 => x"98",
          1654 => x"e0",
          1655 => x"84",
          1656 => x"e0",
          1657 => x"82",
          1658 => x"02",
          1659 => x"0c",
          1660 => x"82",
          1661 => x"8c",
          1662 => x"11",
          1663 => x"2a",
          1664 => x"70",
          1665 => x"51",
          1666 => x"72",
          1667 => x"38",
          1668 => x"e0",
          1669 => x"05",
          1670 => x"39",
          1671 => x"08",
          1672 => x"85",
          1673 => x"82",
          1674 => x"06",
          1675 => x"53",
          1676 => x"80",
          1677 => x"e0",
          1678 => x"05",
          1679 => x"a4",
          1680 => x"08",
          1681 => x"14",
          1682 => x"08",
          1683 => x"82",
          1684 => x"8c",
          1685 => x"08",
          1686 => x"a4",
          1687 => x"08",
          1688 => x"54",
          1689 => x"73",
          1690 => x"74",
          1691 => x"a4",
          1692 => x"08",
          1693 => x"81",
          1694 => x"0c",
          1695 => x"08",
          1696 => x"70",
          1697 => x"08",
          1698 => x"51",
          1699 => x"39",
          1700 => x"08",
          1701 => x"82",
          1702 => x"8c",
          1703 => x"82",
          1704 => x"88",
          1705 => x"81",
          1706 => x"90",
          1707 => x"54",
          1708 => x"82",
          1709 => x"53",
          1710 => x"82",
          1711 => x"8c",
          1712 => x"11",
          1713 => x"8c",
          1714 => x"e0",
          1715 => x"05",
          1716 => x"e0",
          1717 => x"05",
          1718 => x"8a",
          1719 => x"82",
          1720 => x"fc",
          1721 => x"e0",
          1722 => x"05",
          1723 => x"98",
          1724 => x"0d",
          1725 => x"0c",
          1726 => x"a4",
          1727 => x"e0",
          1728 => x"3d",
          1729 => x"a4",
          1730 => x"08",
          1731 => x"70",
          1732 => x"81",
          1733 => x"51",
          1734 => x"2e",
          1735 => x"0b",
          1736 => x"08",
          1737 => x"83",
          1738 => x"e0",
          1739 => x"05",
          1740 => x"33",
          1741 => x"70",
          1742 => x"51",
          1743 => x"80",
          1744 => x"38",
          1745 => x"08",
          1746 => x"82",
          1747 => x"88",
          1748 => x"53",
          1749 => x"70",
          1750 => x"51",
          1751 => x"14",
          1752 => x"a4",
          1753 => x"08",
          1754 => x"81",
          1755 => x"0c",
          1756 => x"08",
          1757 => x"84",
          1758 => x"82",
          1759 => x"f8",
          1760 => x"51",
          1761 => x"39",
          1762 => x"08",
          1763 => x"85",
          1764 => x"82",
          1765 => x"06",
          1766 => x"52",
          1767 => x"80",
          1768 => x"e0",
          1769 => x"05",
          1770 => x"70",
          1771 => x"a4",
          1772 => x"0c",
          1773 => x"e0",
          1774 => x"05",
          1775 => x"82",
          1776 => x"88",
          1777 => x"e0",
          1778 => x"05",
          1779 => x"85",
          1780 => x"a0",
          1781 => x"71",
          1782 => x"ff",
          1783 => x"a4",
          1784 => x"0c",
          1785 => x"82",
          1786 => x"88",
          1787 => x"08",
          1788 => x"0c",
          1789 => x"39",
          1790 => x"08",
          1791 => x"82",
          1792 => x"88",
          1793 => x"94",
          1794 => x"52",
          1795 => x"e0",
          1796 => x"82",
          1797 => x"fc",
          1798 => x"82",
          1799 => x"fc",
          1800 => x"25",
          1801 => x"82",
          1802 => x"88",
          1803 => x"e0",
          1804 => x"05",
          1805 => x"a4",
          1806 => x"08",
          1807 => x"82",
          1808 => x"f0",
          1809 => x"82",
          1810 => x"fc",
          1811 => x"2e",
          1812 => x"95",
          1813 => x"a4",
          1814 => x"08",
          1815 => x"71",
          1816 => x"08",
          1817 => x"93",
          1818 => x"a4",
          1819 => x"08",
          1820 => x"71",
          1821 => x"08",
          1822 => x"82",
          1823 => x"f4",
          1824 => x"82",
          1825 => x"ec",
          1826 => x"13",
          1827 => x"82",
          1828 => x"f8",
          1829 => x"39",
          1830 => x"08",
          1831 => x"8c",
          1832 => x"05",
          1833 => x"82",
          1834 => x"fc",
          1835 => x"81",
          1836 => x"82",
          1837 => x"f8",
          1838 => x"51",
          1839 => x"a4",
          1840 => x"08",
          1841 => x"0c",
          1842 => x"82",
          1843 => x"04",
          1844 => x"08",
          1845 => x"a4",
          1846 => x"0d",
          1847 => x"08",
          1848 => x"82",
          1849 => x"fc",
          1850 => x"e0",
          1851 => x"05",
          1852 => x"a4",
          1853 => x"0c",
          1854 => x"08",
          1855 => x"80",
          1856 => x"38",
          1857 => x"08",
          1858 => x"82",
          1859 => x"fc",
          1860 => x"81",
          1861 => x"e0",
          1862 => x"05",
          1863 => x"a4",
          1864 => x"08",
          1865 => x"e0",
          1866 => x"05",
          1867 => x"81",
          1868 => x"e0",
          1869 => x"05",
          1870 => x"a4",
          1871 => x"08",
          1872 => x"a4",
          1873 => x"0c",
          1874 => x"08",
          1875 => x"82",
          1876 => x"90",
          1877 => x"82",
          1878 => x"f8",
          1879 => x"e0",
          1880 => x"05",
          1881 => x"82",
          1882 => x"90",
          1883 => x"e0",
          1884 => x"05",
          1885 => x"82",
          1886 => x"90",
          1887 => x"e0",
          1888 => x"05",
          1889 => x"81",
          1890 => x"e0",
          1891 => x"05",
          1892 => x"82",
          1893 => x"fc",
          1894 => x"e0",
          1895 => x"05",
          1896 => x"82",
          1897 => x"f8",
          1898 => x"e0",
          1899 => x"05",
          1900 => x"a4",
          1901 => x"08",
          1902 => x"33",
          1903 => x"ae",
          1904 => x"a4",
          1905 => x"08",
          1906 => x"e0",
          1907 => x"05",
          1908 => x"a4",
          1909 => x"08",
          1910 => x"e0",
          1911 => x"05",
          1912 => x"a4",
          1913 => x"08",
          1914 => x"38",
          1915 => x"08",
          1916 => x"51",
          1917 => x"e0",
          1918 => x"05",
          1919 => x"82",
          1920 => x"f8",
          1921 => x"e0",
          1922 => x"05",
          1923 => x"71",
          1924 => x"e0",
          1925 => x"05",
          1926 => x"82",
          1927 => x"fc",
          1928 => x"ad",
          1929 => x"a4",
          1930 => x"08",
          1931 => x"98",
          1932 => x"3d",
          1933 => x"a4",
          1934 => x"e0",
          1935 => x"82",
          1936 => x"fe",
          1937 => x"e0",
          1938 => x"05",
          1939 => x"a4",
          1940 => x"0c",
          1941 => x"08",
          1942 => x"52",
          1943 => x"e0",
          1944 => x"05",
          1945 => x"82",
          1946 => x"fc",
          1947 => x"81",
          1948 => x"51",
          1949 => x"83",
          1950 => x"82",
          1951 => x"fc",
          1952 => x"05",
          1953 => x"08",
          1954 => x"82",
          1955 => x"fc",
          1956 => x"e0",
          1957 => x"05",
          1958 => x"82",
          1959 => x"51",
          1960 => x"82",
          1961 => x"04",
          1962 => x"08",
          1963 => x"a4",
          1964 => x"0d",
          1965 => x"08",
          1966 => x"82",
          1967 => x"fc",
          1968 => x"e0",
          1969 => x"05",
          1970 => x"33",
          1971 => x"08",
          1972 => x"81",
          1973 => x"a4",
          1974 => x"0c",
          1975 => x"08",
          1976 => x"53",
          1977 => x"34",
          1978 => x"08",
          1979 => x"81",
          1980 => x"a4",
          1981 => x"0c",
          1982 => x"06",
          1983 => x"2e",
          1984 => x"be",
          1985 => x"a4",
          1986 => x"08",
          1987 => x"98",
          1988 => x"3d",
          1989 => x"a4",
          1990 => x"e0",
          1991 => x"82",
          1992 => x"fd",
          1993 => x"e0",
          1994 => x"05",
          1995 => x"a4",
          1996 => x"0c",
          1997 => x"08",
          1998 => x"82",
          1999 => x"f8",
          2000 => x"e0",
          2001 => x"05",
          2002 => x"80",
          2003 => x"e0",
          2004 => x"05",
          2005 => x"82",
          2006 => x"90",
          2007 => x"e0",
          2008 => x"05",
          2009 => x"82",
          2010 => x"90",
          2011 => x"e0",
          2012 => x"05",
          2013 => x"ba",
          2014 => x"a4",
          2015 => x"08",
          2016 => x"82",
          2017 => x"f8",
          2018 => x"05",
          2019 => x"08",
          2020 => x"82",
          2021 => x"fc",
          2022 => x"52",
          2023 => x"82",
          2024 => x"fc",
          2025 => x"05",
          2026 => x"08",
          2027 => x"ff",
          2028 => x"e0",
          2029 => x"05",
          2030 => x"e0",
          2031 => x"85",
          2032 => x"e0",
          2033 => x"82",
          2034 => x"02",
          2035 => x"0c",
          2036 => x"82",
          2037 => x"90",
          2038 => x"2e",
          2039 => x"82",
          2040 => x"8c",
          2041 => x"71",
          2042 => x"a4",
          2043 => x"08",
          2044 => x"e0",
          2045 => x"05",
          2046 => x"a4",
          2047 => x"08",
          2048 => x"81",
          2049 => x"54",
          2050 => x"71",
          2051 => x"80",
          2052 => x"e0",
          2053 => x"05",
          2054 => x"33",
          2055 => x"08",
          2056 => x"81",
          2057 => x"a4",
          2058 => x"0c",
          2059 => x"06",
          2060 => x"8d",
          2061 => x"82",
          2062 => x"fc",
          2063 => x"9b",
          2064 => x"a4",
          2065 => x"08",
          2066 => x"e0",
          2067 => x"05",
          2068 => x"a4",
          2069 => x"08",
          2070 => x"38",
          2071 => x"82",
          2072 => x"90",
          2073 => x"2e",
          2074 => x"82",
          2075 => x"88",
          2076 => x"33",
          2077 => x"8d",
          2078 => x"82",
          2079 => x"fc",
          2080 => x"d7",
          2081 => x"a4",
          2082 => x"08",
          2083 => x"e0",
          2084 => x"05",
          2085 => x"a4",
          2086 => x"08",
          2087 => x"52",
          2088 => x"81",
          2089 => x"a4",
          2090 => x"0c",
          2091 => x"e0",
          2092 => x"05",
          2093 => x"82",
          2094 => x"8c",
          2095 => x"33",
          2096 => x"70",
          2097 => x"08",
          2098 => x"53",
          2099 => x"53",
          2100 => x"0b",
          2101 => x"08",
          2102 => x"82",
          2103 => x"fc",
          2104 => x"e0",
          2105 => x"3d",
          2106 => x"a4",
          2107 => x"e0",
          2108 => x"82",
          2109 => x"fa",
          2110 => x"e0",
          2111 => x"05",
          2112 => x"e0",
          2113 => x"05",
          2114 => x"8d",
          2115 => x"98",
          2116 => x"e0",
          2117 => x"05",
          2118 => x"a4",
          2119 => x"08",
          2120 => x"53",
          2121 => x"ec",
          2122 => x"e0",
          2123 => x"82",
          2124 => x"fc",
          2125 => x"82",
          2126 => x"fc",
          2127 => x"38",
          2128 => x"e0",
          2129 => x"05",
          2130 => x"82",
          2131 => x"fc",
          2132 => x"e0",
          2133 => x"05",
          2134 => x"80",
          2135 => x"e0",
          2136 => x"05",
          2137 => x"e0",
          2138 => x"05",
          2139 => x"e0",
          2140 => x"05",
          2141 => x"a2",
          2142 => x"98",
          2143 => x"e0",
          2144 => x"05",
          2145 => x"e0",
          2146 => x"05",
          2147 => x"98",
          2148 => x"0d",
          2149 => x"0c",
          2150 => x"a4",
          2151 => x"e0",
          2152 => x"3d",
          2153 => x"a4",
          2154 => x"08",
          2155 => x"08",
          2156 => x"82",
          2157 => x"8c",
          2158 => x"38",
          2159 => x"e0",
          2160 => x"05",
          2161 => x"39",
          2162 => x"08",
          2163 => x"52",
          2164 => x"e0",
          2165 => x"05",
          2166 => x"82",
          2167 => x"f8",
          2168 => x"81",
          2169 => x"51",
          2170 => x"9f",
          2171 => x"a4",
          2172 => x"08",
          2173 => x"e0",
          2174 => x"05",
          2175 => x"a4",
          2176 => x"08",
          2177 => x"38",
          2178 => x"82",
          2179 => x"f8",
          2180 => x"05",
          2181 => x"08",
          2182 => x"82",
          2183 => x"f8",
          2184 => x"e0",
          2185 => x"05",
          2186 => x"82",
          2187 => x"fc",
          2188 => x"82",
          2189 => x"fc",
          2190 => x"e0",
          2191 => x"3d",
          2192 => x"a4",
          2193 => x"e0",
          2194 => x"82",
          2195 => x"fe",
          2196 => x"e0",
          2197 => x"05",
          2198 => x"a4",
          2199 => x"0c",
          2200 => x"08",
          2201 => x"80",
          2202 => x"38",
          2203 => x"08",
          2204 => x"81",
          2205 => x"a4",
          2206 => x"0c",
          2207 => x"08",
          2208 => x"ff",
          2209 => x"a4",
          2210 => x"0c",
          2211 => x"08",
          2212 => x"80",
          2213 => x"82",
          2214 => x"8c",
          2215 => x"70",
          2216 => x"08",
          2217 => x"52",
          2218 => x"34",
          2219 => x"08",
          2220 => x"81",
          2221 => x"a4",
          2222 => x"0c",
          2223 => x"82",
          2224 => x"88",
          2225 => x"82",
          2226 => x"51",
          2227 => x"82",
          2228 => x"04",
          2229 => x"08",
          2230 => x"a4",
          2231 => x"0d",
          2232 => x"08",
          2233 => x"52",
          2234 => x"08",
          2235 => x"51",
          2236 => x"e0",
          2237 => x"82",
          2238 => x"53",
          2239 => x"82",
          2240 => x"04",
          2241 => x"08",
          2242 => x"a4",
          2243 => x"0d",
          2244 => x"e0",
          2245 => x"05",
          2246 => x"a4",
          2247 => x"08",
          2248 => x"38",
          2249 => x"08",
          2250 => x"51",
          2251 => x"82",
          2252 => x"70",
          2253 => x"08",
          2254 => x"52",
          2255 => x"e0",
          2256 => x"05",
          2257 => x"a4",
          2258 => x"0c",
          2259 => x"08",
          2260 => x"80",
          2261 => x"82",
          2262 => x"88",
          2263 => x"83",
          2264 => x"e0",
          2265 => x"e0",
          2266 => x"05",
          2267 => x"82",
          2268 => x"e0",
          2269 => x"97",
          2270 => x"a4",
          2271 => x"08",
          2272 => x"08",
          2273 => x"31",
          2274 => x"08",
          2275 => x"82",
          2276 => x"e0",
          2277 => x"e0",
          2278 => x"05",
          2279 => x"a4",
          2280 => x"08",
          2281 => x"71",
          2282 => x"08",
          2283 => x"27",
          2284 => x"0b",
          2285 => x"08",
          2286 => x"82",
          2287 => x"e0",
          2288 => x"05",
          2289 => x"52",
          2290 => x"a4",
          2291 => x"08",
          2292 => x"06",
          2293 => x"e0",
          2294 => x"05",
          2295 => x"e0",
          2296 => x"05",
          2297 => x"af",
          2298 => x"a4",
          2299 => x"08",
          2300 => x"e0",
          2301 => x"05",
          2302 => x"a4",
          2303 => x"08",
          2304 => x"08",
          2305 => x"2a",
          2306 => x"08",
          2307 => x"82",
          2308 => x"fc",
          2309 => x"e0",
          2310 => x"05",
          2311 => x"e0",
          2312 => x"05",
          2313 => x"82",
          2314 => x"88",
          2315 => x"80",
          2316 => x"a4",
          2317 => x"0c",
          2318 => x"08",
          2319 => x"80",
          2320 => x"38",
          2321 => x"08",
          2322 => x"10",
          2323 => x"08",
          2324 => x"ff",
          2325 => x"a4",
          2326 => x"08",
          2327 => x"73",
          2328 => x"a4",
          2329 => x"0c",
          2330 => x"08",
          2331 => x"10",
          2332 => x"a4",
          2333 => x"08",
          2334 => x"a4",
          2335 => x"0c",
          2336 => x"08",
          2337 => x"82",
          2338 => x"f4",
          2339 => x"ff",
          2340 => x"a4",
          2341 => x"08",
          2342 => x"71",
          2343 => x"a4",
          2344 => x"0c",
          2345 => x"08",
          2346 => x"81",
          2347 => x"a4",
          2348 => x"0c",
          2349 => x"08",
          2350 => x"82",
          2351 => x"ec",
          2352 => x"82",
          2353 => x"f4",
          2354 => x"31",
          2355 => x"08",
          2356 => x"82",
          2357 => x"f8",
          2358 => x"05",
          2359 => x"08",
          2360 => x"51",
          2361 => x"51",
          2362 => x"fe",
          2363 => x"e0",
          2364 => x"05",
          2365 => x"82",
          2366 => x"f0",
          2367 => x"82",
          2368 => x"88",
          2369 => x"e0",
          2370 => x"05",
          2371 => x"e0",
          2372 => x"05",
          2373 => x"82",
          2374 => x"e8",
          2375 => x"e0",
          2376 => x"3d",
          2377 => x"a4",
          2378 => x"e0",
          2379 => x"82",
          2380 => x"f8",
          2381 => x"e0",
          2382 => x"05",
          2383 => x"a4",
          2384 => x"0c",
          2385 => x"08",
          2386 => x"fc",
          2387 => x"51",
          2388 => x"90",
          2389 => x"a4",
          2390 => x"0c",
          2391 => x"0b",
          2392 => x"08",
          2393 => x"82",
          2394 => x"f0",
          2395 => x"e0",
          2396 => x"05",
          2397 => x"82",
          2398 => x"f8",
          2399 => x"82",
          2400 => x"fc",
          2401 => x"2a",
          2402 => x"08",
          2403 => x"82",
          2404 => x"f8",
          2405 => x"e0",
          2406 => x"05",
          2407 => x"a4",
          2408 => x"08",
          2409 => x"06",
          2410 => x"8c",
          2411 => x"82",
          2412 => x"ec",
          2413 => x"39",
          2414 => x"e0",
          2415 => x"05",
          2416 => x"a4",
          2417 => x"08",
          2418 => x"08",
          2419 => x"88",
          2420 => x"a4",
          2421 => x"08",
          2422 => x"a4",
          2423 => x"08",
          2424 => x"e0",
          2425 => x"05",
          2426 => x"a4",
          2427 => x"08",
          2428 => x"08",
          2429 => x"05",
          2430 => x"08",
          2431 => x"82",
          2432 => x"fc",
          2433 => x"f0",
          2434 => x"70",
          2435 => x"0b",
          2436 => x"08",
          2437 => x"8a",
          2438 => x"82",
          2439 => x"e8",
          2440 => x"e0",
          2441 => x"05",
          2442 => x"a4",
          2443 => x"0c",
          2444 => x"e0",
          2445 => x"05",
          2446 => x"e0",
          2447 => x"05",
          2448 => x"82",
          2449 => x"fc",
          2450 => x"e0",
          2451 => x"05",
          2452 => x"a4",
          2453 => x"08",
          2454 => x"a4",
          2455 => x"0c",
          2456 => x"08",
          2457 => x"8c",
          2458 => x"70",
          2459 => x"0b",
          2460 => x"08",
          2461 => x"8a",
          2462 => x"82",
          2463 => x"e4",
          2464 => x"e0",
          2465 => x"05",
          2466 => x"a4",
          2467 => x"0c",
          2468 => x"e0",
          2469 => x"05",
          2470 => x"e0",
          2471 => x"05",
          2472 => x"82",
          2473 => x"fc",
          2474 => x"e0",
          2475 => x"05",
          2476 => x"a4",
          2477 => x"08",
          2478 => x"a4",
          2479 => x"0c",
          2480 => x"e0",
          2481 => x"05",
          2482 => x"e0",
          2483 => x"05",
          2484 => x"70",
          2485 => x"81",
          2486 => x"70",
          2487 => x"e0",
          2488 => x"05",
          2489 => x"70",
          2490 => x"0c",
          2491 => x"51",
          2492 => x"53",
          2493 => x"0d",
          2494 => x"0c",
          2495 => x"a4",
          2496 => x"e0",
          2497 => x"3d",
          2498 => x"a4",
          2499 => x"08",
          2500 => x"a4",
          2501 => x"08",
          2502 => x"3f",
          2503 => x"08",
          2504 => x"a4",
          2505 => x"08",
          2506 => x"a4",
          2507 => x"08",
          2508 => x"82",
          2509 => x"51",
          2510 => x"3d",
          2511 => x"a4",
          2512 => x"e0",
          2513 => x"82",
          2514 => x"fe",
          2515 => x"e0",
          2516 => x"05",
          2517 => x"e0",
          2518 => x"05",
          2519 => x"3f",
          2520 => x"08",
          2521 => x"98",
          2522 => x"3d",
          2523 => x"a4",
          2524 => x"e0",
          2525 => x"82",
          2526 => x"f6",
          2527 => x"0b",
          2528 => x"08",
          2529 => x"82",
          2530 => x"8c",
          2531 => x"2e",
          2532 => x"e0",
          2533 => x"05",
          2534 => x"8e",
          2535 => x"98",
          2536 => x"e0",
          2537 => x"05",
          2538 => x"39",
          2539 => x"08",
          2540 => x"82",
          2541 => x"e4",
          2542 => x"e0",
          2543 => x"05",
          2544 => x"a3",
          2545 => x"a4",
          2546 => x"08",
          2547 => x"3f",
          2548 => x"08",
          2549 => x"08",
          2550 => x"71",
          2551 => x"a4",
          2552 => x"0c",
          2553 => x"82",
          2554 => x"e4",
          2555 => x"e0",
          2556 => x"05",
          2557 => x"e0",
          2558 => x"05",
          2559 => x"a4",
          2560 => x"08",
          2561 => x"08",
          2562 => x"82",
          2563 => x"fc",
          2564 => x"05",
          2565 => x"e0",
          2566 => x"05",
          2567 => x"38",
          2568 => x"08",
          2569 => x"70",
          2570 => x"08",
          2571 => x"52",
          2572 => x"82",
          2573 => x"fc",
          2574 => x"05",
          2575 => x"e0",
          2576 => x"05",
          2577 => x"81",
          2578 => x"80",
          2579 => x"a4",
          2580 => x"0c",
          2581 => x"82",
          2582 => x"f8",
          2583 => x"05",
          2584 => x"08",
          2585 => x"82",
          2586 => x"88",
          2587 => x"e0",
          2588 => x"05",
          2589 => x"e0",
          2590 => x"05",
          2591 => x"a4",
          2592 => x"08",
          2593 => x"08",
          2594 => x"31",
          2595 => x"08",
          2596 => x"71",
          2597 => x"a4",
          2598 => x"0c",
          2599 => x"82",
          2600 => x"f0",
          2601 => x"e0",
          2602 => x"05",
          2603 => x"81",
          2604 => x"e0",
          2605 => x"05",
          2606 => x"e0",
          2607 => x"05",
          2608 => x"82",
          2609 => x"88",
          2610 => x"2a",
          2611 => x"82",
          2612 => x"f4",
          2613 => x"e0",
          2614 => x"05",
          2615 => x"82",
          2616 => x"f0",
          2617 => x"82",
          2618 => x"88",
          2619 => x"e0",
          2620 => x"05",
          2621 => x"a4",
          2622 => x"08",
          2623 => x"82",
          2624 => x"fc",
          2625 => x"05",
          2626 => x"82",
          2627 => x"ec",
          2628 => x"e0",
          2629 => x"05",
          2630 => x"82",
          2631 => x"f0",
          2632 => x"e0",
          2633 => x"05",
          2634 => x"a4",
          2635 => x"08",
          2636 => x"a4",
          2637 => x"08",
          2638 => x"e0",
          2639 => x"05",
          2640 => x"a4",
          2641 => x"08",
          2642 => x"e0",
          2643 => x"05",
          2644 => x"55",
          2645 => x"53",
          2646 => x"39",
          2647 => x"08",
          2648 => x"70",
          2649 => x"08",
          2650 => x"52",
          2651 => x"08",
          2652 => x"82",
          2653 => x"8c",
          2654 => x"e0",
          2655 => x"82",
          2656 => x"02",
          2657 => x"0c",
          2658 => x"9f",
          2659 => x"a4",
          2660 => x"0c",
          2661 => x"08",
          2662 => x"82",
          2663 => x"fc",
          2664 => x"82",
          2665 => x"f8",
          2666 => x"e0",
          2667 => x"05",
          2668 => x"a4",
          2669 => x"08",
          2670 => x"a4",
          2671 => x"0c",
          2672 => x"08",
          2673 => x"82",
          2674 => x"f8",
          2675 => x"70",
          2676 => x"08",
          2677 => x"31",
          2678 => x"08",
          2679 => x"82",
          2680 => x"8c",
          2681 => x"e0",
          2682 => x"05",
          2683 => x"82",
          2684 => x"f4",
          2685 => x"82",
          2686 => x"8c",
          2687 => x"e0",
          2688 => x"05",
          2689 => x"a4",
          2690 => x"08",
          2691 => x"a4",
          2692 => x"0c",
          2693 => x"08",
          2694 => x"54",
          2695 => x"08",
          2696 => x"53",
          2697 => x"ac",
          2698 => x"98",
          2699 => x"e0",
          2700 => x"05",
          2701 => x"82",
          2702 => x"f8",
          2703 => x"70",
          2704 => x"0c",
          2705 => x"87",
          2706 => x"e0",
          2707 => x"82",
          2708 => x"02",
          2709 => x"0c",
          2710 => x"80",
          2711 => x"a4",
          2712 => x"34",
          2713 => x"08",
          2714 => x"53",
          2715 => x"82",
          2716 => x"88",
          2717 => x"08",
          2718 => x"33",
          2719 => x"e0",
          2720 => x"05",
          2721 => x"ff",
          2722 => x"a0",
          2723 => x"06",
          2724 => x"e0",
          2725 => x"05",
          2726 => x"81",
          2727 => x"53",
          2728 => x"e0",
          2729 => x"05",
          2730 => x"ad",
          2731 => x"06",
          2732 => x"0b",
          2733 => x"08",
          2734 => x"82",
          2735 => x"88",
          2736 => x"08",
          2737 => x"0c",
          2738 => x"53",
          2739 => x"e0",
          2740 => x"05",
          2741 => x"a4",
          2742 => x"33",
          2743 => x"2e",
          2744 => x"81",
          2745 => x"e0",
          2746 => x"05",
          2747 => x"81",
          2748 => x"70",
          2749 => x"72",
          2750 => x"a4",
          2751 => x"34",
          2752 => x"08",
          2753 => x"82",
          2754 => x"e8",
          2755 => x"e0",
          2756 => x"05",
          2757 => x"2e",
          2758 => x"e0",
          2759 => x"05",
          2760 => x"2e",
          2761 => x"cd",
          2762 => x"82",
          2763 => x"f4",
          2764 => x"e0",
          2765 => x"05",
          2766 => x"81",
          2767 => x"70",
          2768 => x"72",
          2769 => x"a4",
          2770 => x"34",
          2771 => x"82",
          2772 => x"a4",
          2773 => x"34",
          2774 => x"08",
          2775 => x"70",
          2776 => x"71",
          2777 => x"51",
          2778 => x"82",
          2779 => x"f8",
          2780 => x"fe",
          2781 => x"a4",
          2782 => x"33",
          2783 => x"26",
          2784 => x"0b",
          2785 => x"08",
          2786 => x"83",
          2787 => x"e0",
          2788 => x"05",
          2789 => x"73",
          2790 => x"82",
          2791 => x"f8",
          2792 => x"72",
          2793 => x"38",
          2794 => x"0b",
          2795 => x"08",
          2796 => x"82",
          2797 => x"0b",
          2798 => x"08",
          2799 => x"b2",
          2800 => x"a4",
          2801 => x"33",
          2802 => x"27",
          2803 => x"e0",
          2804 => x"05",
          2805 => x"b9",
          2806 => x"8d",
          2807 => x"82",
          2808 => x"ec",
          2809 => x"a5",
          2810 => x"82",
          2811 => x"f4",
          2812 => x"0b",
          2813 => x"08",
          2814 => x"82",
          2815 => x"f8",
          2816 => x"a0",
          2817 => x"cf",
          2818 => x"a4",
          2819 => x"33",
          2820 => x"73",
          2821 => x"82",
          2822 => x"f8",
          2823 => x"11",
          2824 => x"82",
          2825 => x"f8",
          2826 => x"e0",
          2827 => x"05",
          2828 => x"51",
          2829 => x"e0",
          2830 => x"05",
          2831 => x"a4",
          2832 => x"33",
          2833 => x"27",
          2834 => x"e0",
          2835 => x"05",
          2836 => x"51",
          2837 => x"e0",
          2838 => x"05",
          2839 => x"a4",
          2840 => x"33",
          2841 => x"26",
          2842 => x"0b",
          2843 => x"08",
          2844 => x"81",
          2845 => x"e0",
          2846 => x"05",
          2847 => x"a4",
          2848 => x"33",
          2849 => x"74",
          2850 => x"80",
          2851 => x"a4",
          2852 => x"0c",
          2853 => x"82",
          2854 => x"f4",
          2855 => x"82",
          2856 => x"fc",
          2857 => x"82",
          2858 => x"f8",
          2859 => x"12",
          2860 => x"08",
          2861 => x"82",
          2862 => x"88",
          2863 => x"08",
          2864 => x"0c",
          2865 => x"51",
          2866 => x"72",
          2867 => x"a4",
          2868 => x"34",
          2869 => x"82",
          2870 => x"f0",
          2871 => x"72",
          2872 => x"38",
          2873 => x"08",
          2874 => x"30",
          2875 => x"08",
          2876 => x"82",
          2877 => x"8c",
          2878 => x"e0",
          2879 => x"05",
          2880 => x"53",
          2881 => x"e0",
          2882 => x"05",
          2883 => x"a4",
          2884 => x"08",
          2885 => x"0c",
          2886 => x"82",
          2887 => x"04",
          2888 => x"08",
          2889 => x"a4",
          2890 => x"0d",
          2891 => x"e0",
          2892 => x"05",
          2893 => x"a4",
          2894 => x"08",
          2895 => x"0c",
          2896 => x"08",
          2897 => x"70",
          2898 => x"72",
          2899 => x"82",
          2900 => x"f8",
          2901 => x"81",
          2902 => x"72",
          2903 => x"81",
          2904 => x"82",
          2905 => x"88",
          2906 => x"08",
          2907 => x"0c",
          2908 => x"82",
          2909 => x"f8",
          2910 => x"72",
          2911 => x"81",
          2912 => x"81",
          2913 => x"a4",
          2914 => x"34",
          2915 => x"08",
          2916 => x"70",
          2917 => x"71",
          2918 => x"51",
          2919 => x"82",
          2920 => x"f8",
          2921 => x"e0",
          2922 => x"05",
          2923 => x"b0",
          2924 => x"06",
          2925 => x"82",
          2926 => x"88",
          2927 => x"08",
          2928 => x"0c",
          2929 => x"53",
          2930 => x"e0",
          2931 => x"05",
          2932 => x"a4",
          2933 => x"33",
          2934 => x"08",
          2935 => x"82",
          2936 => x"e8",
          2937 => x"e2",
          2938 => x"82",
          2939 => x"e8",
          2940 => x"f8",
          2941 => x"80",
          2942 => x"0b",
          2943 => x"08",
          2944 => x"82",
          2945 => x"88",
          2946 => x"08",
          2947 => x"0c",
          2948 => x"53",
          2949 => x"e0",
          2950 => x"05",
          2951 => x"39",
          2952 => x"e0",
          2953 => x"05",
          2954 => x"a4",
          2955 => x"08",
          2956 => x"05",
          2957 => x"08",
          2958 => x"33",
          2959 => x"08",
          2960 => x"80",
          2961 => x"e0",
          2962 => x"05",
          2963 => x"a0",
          2964 => x"81",
          2965 => x"a4",
          2966 => x"0c",
          2967 => x"82",
          2968 => x"f8",
          2969 => x"af",
          2970 => x"38",
          2971 => x"08",
          2972 => x"53",
          2973 => x"83",
          2974 => x"80",
          2975 => x"a4",
          2976 => x"0c",
          2977 => x"88",
          2978 => x"a4",
          2979 => x"34",
          2980 => x"e0",
          2981 => x"05",
          2982 => x"73",
          2983 => x"82",
          2984 => x"f8",
          2985 => x"72",
          2986 => x"38",
          2987 => x"0b",
          2988 => x"08",
          2989 => x"82",
          2990 => x"0b",
          2991 => x"08",
          2992 => x"80",
          2993 => x"a4",
          2994 => x"0c",
          2995 => x"08",
          2996 => x"53",
          2997 => x"81",
          2998 => x"e0",
          2999 => x"05",
          3000 => x"e0",
          3001 => x"38",
          3002 => x"08",
          3003 => x"e0",
          3004 => x"72",
          3005 => x"08",
          3006 => x"82",
          3007 => x"f8",
          3008 => x"11",
          3009 => x"82",
          3010 => x"f8",
          3011 => x"e0",
          3012 => x"05",
          3013 => x"73",
          3014 => x"82",
          3015 => x"f8",
          3016 => x"11",
          3017 => x"82",
          3018 => x"f8",
          3019 => x"e0",
          3020 => x"05",
          3021 => x"89",
          3022 => x"80",
          3023 => x"a4",
          3024 => x"0c",
          3025 => x"82",
          3026 => x"f8",
          3027 => x"e0",
          3028 => x"05",
          3029 => x"72",
          3030 => x"38",
          3031 => x"e0",
          3032 => x"05",
          3033 => x"39",
          3034 => x"08",
          3035 => x"70",
          3036 => x"08",
          3037 => x"29",
          3038 => x"08",
          3039 => x"70",
          3040 => x"a4",
          3041 => x"0c",
          3042 => x"08",
          3043 => x"70",
          3044 => x"71",
          3045 => x"51",
          3046 => x"53",
          3047 => x"e0",
          3048 => x"05",
          3049 => x"39",
          3050 => x"08",
          3051 => x"53",
          3052 => x"90",
          3053 => x"a4",
          3054 => x"08",
          3055 => x"a4",
          3056 => x"0c",
          3057 => x"08",
          3058 => x"82",
          3059 => x"fc",
          3060 => x"0c",
          3061 => x"82",
          3062 => x"ec",
          3063 => x"e0",
          3064 => x"05",
          3065 => x"98",
          3066 => x"0d",
          3067 => x"0c",
          3068 => x"0d",
          3069 => x"70",
          3070 => x"74",
          3071 => x"df",
          3072 => x"77",
          3073 => x"85",
          3074 => x"80",
          3075 => x"33",
          3076 => x"2e",
          3077 => x"86",
          3078 => x"55",
          3079 => x"57",
          3080 => x"82",
          3081 => x"70",
          3082 => x"dc",
          3083 => x"e0",
          3084 => x"e0",
          3085 => x"75",
          3086 => x"52",
          3087 => x"3f",
          3088 => x"08",
          3089 => x"16",
          3090 => x"81",
          3091 => x"38",
          3092 => x"81",
          3093 => x"54",
          3094 => x"c4",
          3095 => x"73",
          3096 => x"0c",
          3097 => x"04",
          3098 => x"82",
          3099 => x"04",
          3100 => x"73",
          3101 => x"26",
          3102 => x"71",
          3103 => x"b7",
          3104 => x"71",
          3105 => x"bd",
          3106 => x"80",
          3107 => x"f0",
          3108 => x"39",
          3109 => x"51",
          3110 => x"82",
          3111 => x"80",
          3112 => x"be",
          3113 => x"e4",
          3114 => x"b0",
          3115 => x"39",
          3116 => x"51",
          3117 => x"82",
          3118 => x"80",
          3119 => x"be",
          3120 => x"c8",
          3121 => x"84",
          3122 => x"39",
          3123 => x"51",
          3124 => x"bf",
          3125 => x"39",
          3126 => x"51",
          3127 => x"bf",
          3128 => x"39",
          3129 => x"51",
          3130 => x"c0",
          3131 => x"39",
          3132 => x"51",
          3133 => x"c0",
          3134 => x"39",
          3135 => x"51",
          3136 => x"c0",
          3137 => x"39",
          3138 => x"51",
          3139 => x"83",
          3140 => x"fb",
          3141 => x"79",
          3142 => x"87",
          3143 => x"38",
          3144 => x"87",
          3145 => x"90",
          3146 => x"52",
          3147 => x"a4",
          3148 => x"98",
          3149 => x"51",
          3150 => x"82",
          3151 => x"54",
          3152 => x"52",
          3153 => x"51",
          3154 => x"3f",
          3155 => x"04",
          3156 => x"66",
          3157 => x"80",
          3158 => x"5b",
          3159 => x"78",
          3160 => x"07",
          3161 => x"57",
          3162 => x"56",
          3163 => x"26",
          3164 => x"56",
          3165 => x"70",
          3166 => x"51",
          3167 => x"74",
          3168 => x"81",
          3169 => x"8c",
          3170 => x"56",
          3171 => x"3f",
          3172 => x"08",
          3173 => x"98",
          3174 => x"82",
          3175 => x"87",
          3176 => x"0c",
          3177 => x"08",
          3178 => x"d4",
          3179 => x"80",
          3180 => x"75",
          3181 => x"d5",
          3182 => x"98",
          3183 => x"e0",
          3184 => x"38",
          3185 => x"80",
          3186 => x"74",
          3187 => x"59",
          3188 => x"96",
          3189 => x"51",
          3190 => x"3f",
          3191 => x"78",
          3192 => x"7b",
          3193 => x"2a",
          3194 => x"57",
          3195 => x"80",
          3196 => x"82",
          3197 => x"87",
          3198 => x"08",
          3199 => x"fe",
          3200 => x"56",
          3201 => x"98",
          3202 => x"0d",
          3203 => x"0d",
          3204 => x"05",
          3205 => x"58",
          3206 => x"80",
          3207 => x"7a",
          3208 => x"3f",
          3209 => x"08",
          3210 => x"80",
          3211 => x"76",
          3212 => x"38",
          3213 => x"fb",
          3214 => x"55",
          3215 => x"e0",
          3216 => x"52",
          3217 => x"2d",
          3218 => x"08",
          3219 => x"78",
          3220 => x"e0",
          3221 => x"3d",
          3222 => x"3d",
          3223 => x"63",
          3224 => x"80",
          3225 => x"73",
          3226 => x"41",
          3227 => x"5e",
          3228 => x"a4",
          3229 => x"3f",
          3230 => x"08",
          3231 => x"53",
          3232 => x"a8",
          3233 => x"90",
          3234 => x"d0",
          3235 => x"86",
          3236 => x"82",
          3237 => x"58",
          3238 => x"c1",
          3239 => x"ae",
          3240 => x"c1",
          3241 => x"ae",
          3242 => x"55",
          3243 => x"81",
          3244 => x"90",
          3245 => x"7b",
          3246 => x"38",
          3247 => x"74",
          3248 => x"7a",
          3249 => x"72",
          3250 => x"c1",
          3251 => x"ae",
          3252 => x"39",
          3253 => x"51",
          3254 => x"3f",
          3255 => x"80",
          3256 => x"19",
          3257 => x"27",
          3258 => x"08",
          3259 => x"c4",
          3260 => x"99",
          3261 => x"82",
          3262 => x"ff",
          3263 => x"84",
          3264 => x"39",
          3265 => x"72",
          3266 => x"38",
          3267 => x"82",
          3268 => x"ff",
          3269 => x"89",
          3270 => x"ec",
          3271 => x"ed",
          3272 => x"55",
          3273 => x"08",
          3274 => x"cd",
          3275 => x"fc",
          3276 => x"f0",
          3277 => x"d5",
          3278 => x"74",
          3279 => x"c6",
          3280 => x"70",
          3281 => x"80",
          3282 => x"27",
          3283 => x"56",
          3284 => x"74",
          3285 => x"81",
          3286 => x"06",
          3287 => x"06",
          3288 => x"80",
          3289 => x"73",
          3290 => x"8a",
          3291 => x"fc",
          3292 => x"51",
          3293 => x"fb",
          3294 => x"a0",
          3295 => x"3f",
          3296 => x"ff",
          3297 => x"c1",
          3298 => x"8c",
          3299 => x"78",
          3300 => x"80",
          3301 => x"3f",
          3302 => x"08",
          3303 => x"98",
          3304 => x"76",
          3305 => x"81",
          3306 => x"80",
          3307 => x"3f",
          3308 => x"08",
          3309 => x"98",
          3310 => x"32",
          3311 => x"9b",
          3312 => x"70",
          3313 => x"75",
          3314 => x"58",
          3315 => x"51",
          3316 => x"24",
          3317 => x"9b",
          3318 => x"38",
          3319 => x"72",
          3320 => x"b4",
          3321 => x"72",
          3322 => x"0c",
          3323 => x"04",
          3324 => x"02",
          3325 => x"55",
          3326 => x"be",
          3327 => x"f8",
          3328 => x"fc",
          3329 => x"85",
          3330 => x"e8",
          3331 => x"d8",
          3332 => x"84",
          3333 => x"90",
          3334 => x"e9",
          3335 => x"c2",
          3336 => x"ab",
          3337 => x"80",
          3338 => x"a2",
          3339 => x"3d",
          3340 => x"3d",
          3341 => x"96",
          3342 => x"a6",
          3343 => x"51",
          3344 => x"82",
          3345 => x"9a",
          3346 => x"51",
          3347 => x"72",
          3348 => x"81",
          3349 => x"71",
          3350 => x"38",
          3351 => x"a1",
          3352 => x"cc",
          3353 => x"3f",
          3354 => x"95",
          3355 => x"2a",
          3356 => x"51",
          3357 => x"2e",
          3358 => x"51",
          3359 => x"82",
          3360 => x"9a",
          3361 => x"51",
          3362 => x"72",
          3363 => x"81",
          3364 => x"71",
          3365 => x"38",
          3366 => x"e5",
          3367 => x"ec",
          3368 => x"3f",
          3369 => x"d9",
          3370 => x"2a",
          3371 => x"51",
          3372 => x"2e",
          3373 => x"51",
          3374 => x"82",
          3375 => x"99",
          3376 => x"51",
          3377 => x"72",
          3378 => x"81",
          3379 => x"71",
          3380 => x"38",
          3381 => x"a9",
          3382 => x"94",
          3383 => x"3f",
          3384 => x"9d",
          3385 => x"2a",
          3386 => x"51",
          3387 => x"2e",
          3388 => x"51",
          3389 => x"82",
          3390 => x"99",
          3391 => x"51",
          3392 => x"72",
          3393 => x"81",
          3394 => x"71",
          3395 => x"38",
          3396 => x"ed",
          3397 => x"bc",
          3398 => x"3f",
          3399 => x"e1",
          3400 => x"2a",
          3401 => x"51",
          3402 => x"2e",
          3403 => x"51",
          3404 => x"82",
          3405 => x"98",
          3406 => x"51",
          3407 => x"a4",
          3408 => x"3d",
          3409 => x"3d",
          3410 => x"84",
          3411 => x"33",
          3412 => x"56",
          3413 => x"51",
          3414 => x"0b",
          3415 => x"9c",
          3416 => x"a9",
          3417 => x"82",
          3418 => x"82",
          3419 => x"81",
          3420 => x"82",
          3421 => x"30",
          3422 => x"98",
          3423 => x"25",
          3424 => x"51",
          3425 => x"0b",
          3426 => x"9c",
          3427 => x"82",
          3428 => x"54",
          3429 => x"09",
          3430 => x"38",
          3431 => x"53",
          3432 => x"51",
          3433 => x"3f",
          3434 => x"08",
          3435 => x"38",
          3436 => x"08",
          3437 => x"3f",
          3438 => x"f7",
          3439 => x"97",
          3440 => x"0b",
          3441 => x"db",
          3442 => x"0b",
          3443 => x"33",
          3444 => x"2e",
          3445 => x"8c",
          3446 => x"9c",
          3447 => x"75",
          3448 => x"3f",
          3449 => x"e0",
          3450 => x"3d",
          3451 => x"3d",
          3452 => x"41",
          3453 => x"82",
          3454 => x"5f",
          3455 => x"51",
          3456 => x"3f",
          3457 => x"08",
          3458 => x"59",
          3459 => x"09",
          3460 => x"38",
          3461 => x"83",
          3462 => x"a8",
          3463 => x"d1",
          3464 => x"53",
          3465 => x"e1",
          3466 => x"89",
          3467 => x"e0",
          3468 => x"2e",
          3469 => x"c4",
          3470 => x"e5",
          3471 => x"41",
          3472 => x"e4",
          3473 => x"c5",
          3474 => x"70",
          3475 => x"f8",
          3476 => x"fd",
          3477 => x"3d",
          3478 => x"51",
          3479 => x"82",
          3480 => x"90",
          3481 => x"2c",
          3482 => x"80",
          3483 => x"a5",
          3484 => x"c2",
          3485 => x"78",
          3486 => x"d2",
          3487 => x"24",
          3488 => x"80",
          3489 => x"38",
          3490 => x"80",
          3491 => x"dc",
          3492 => x"c0",
          3493 => x"38",
          3494 => x"24",
          3495 => x"78",
          3496 => x"8c",
          3497 => x"39",
          3498 => x"2e",
          3499 => x"78",
          3500 => x"92",
          3501 => x"c3",
          3502 => x"38",
          3503 => x"2e",
          3504 => x"8a",
          3505 => x"81",
          3506 => x"8d",
          3507 => x"83",
          3508 => x"78",
          3509 => x"89",
          3510 => x"90",
          3511 => x"85",
          3512 => x"38",
          3513 => x"b5",
          3514 => x"11",
          3515 => x"05",
          3516 => x"3f",
          3517 => x"08",
          3518 => x"c5",
          3519 => x"fe",
          3520 => x"ff",
          3521 => x"ec",
          3522 => x"e0",
          3523 => x"2e",
          3524 => x"b5",
          3525 => x"11",
          3526 => x"05",
          3527 => x"3f",
          3528 => x"08",
          3529 => x"e0",
          3530 => x"82",
          3531 => x"ff",
          3532 => x"64",
          3533 => x"79",
          3534 => x"ec",
          3535 => x"78",
          3536 => x"05",
          3537 => x"7a",
          3538 => x"81",
          3539 => x"3d",
          3540 => x"53",
          3541 => x"51",
          3542 => x"82",
          3543 => x"80",
          3544 => x"38",
          3545 => x"fc",
          3546 => x"84",
          3547 => x"b0",
          3548 => x"98",
          3549 => x"fd",
          3550 => x"3d",
          3551 => x"53",
          3552 => x"51",
          3553 => x"82",
          3554 => x"80",
          3555 => x"38",
          3556 => x"51",
          3557 => x"3f",
          3558 => x"64",
          3559 => x"38",
          3560 => x"70",
          3561 => x"33",
          3562 => x"81",
          3563 => x"39",
          3564 => x"80",
          3565 => x"84",
          3566 => x"e4",
          3567 => x"98",
          3568 => x"fc",
          3569 => x"3d",
          3570 => x"53",
          3571 => x"51",
          3572 => x"82",
          3573 => x"80",
          3574 => x"38",
          3575 => x"f8",
          3576 => x"84",
          3577 => x"b8",
          3578 => x"98",
          3579 => x"fc",
          3580 => x"c5",
          3581 => x"a4",
          3582 => x"5a",
          3583 => x"a8",
          3584 => x"33",
          3585 => x"5a",
          3586 => x"2e",
          3587 => x"55",
          3588 => x"33",
          3589 => x"82",
          3590 => x"ff",
          3591 => x"81",
          3592 => x"05",
          3593 => x"39",
          3594 => x"8e",
          3595 => x"39",
          3596 => x"80",
          3597 => x"84",
          3598 => x"e4",
          3599 => x"98",
          3600 => x"38",
          3601 => x"33",
          3602 => x"2e",
          3603 => x"de",
          3604 => x"80",
          3605 => x"de",
          3606 => x"78",
          3607 => x"38",
          3608 => x"08",
          3609 => x"82",
          3610 => x"59",
          3611 => x"88",
          3612 => x"c4",
          3613 => x"39",
          3614 => x"33",
          3615 => x"2e",
          3616 => x"de",
          3617 => x"9a",
          3618 => x"fa",
          3619 => x"80",
          3620 => x"82",
          3621 => x"45",
          3622 => x"de",
          3623 => x"80",
          3624 => x"3d",
          3625 => x"53",
          3626 => x"51",
          3627 => x"82",
          3628 => x"80",
          3629 => x"de",
          3630 => x"78",
          3631 => x"38",
          3632 => x"08",
          3633 => x"39",
          3634 => x"33",
          3635 => x"2e",
          3636 => x"de",
          3637 => x"bb",
          3638 => x"fe",
          3639 => x"80",
          3640 => x"82",
          3641 => x"44",
          3642 => x"de",
          3643 => x"78",
          3644 => x"38",
          3645 => x"08",
          3646 => x"82",
          3647 => x"59",
          3648 => x"88",
          3649 => x"d8",
          3650 => x"39",
          3651 => x"08",
          3652 => x"b5",
          3653 => x"11",
          3654 => x"05",
          3655 => x"3f",
          3656 => x"08",
          3657 => x"38",
          3658 => x"5c",
          3659 => x"83",
          3660 => x"7a",
          3661 => x"30",
          3662 => x"9f",
          3663 => x"06",
          3664 => x"5a",
          3665 => x"88",
          3666 => x"2e",
          3667 => x"43",
          3668 => x"51",
          3669 => x"3f",
          3670 => x"54",
          3671 => x"52",
          3672 => x"f6",
          3673 => x"bc",
          3674 => x"39",
          3675 => x"80",
          3676 => x"84",
          3677 => x"a8",
          3678 => x"98",
          3679 => x"f9",
          3680 => x"3d",
          3681 => x"53",
          3682 => x"51",
          3683 => x"82",
          3684 => x"80",
          3685 => x"64",
          3686 => x"cf",
          3687 => x"34",
          3688 => x"45",
          3689 => x"fc",
          3690 => x"84",
          3691 => x"f0",
          3692 => x"98",
          3693 => x"f9",
          3694 => x"70",
          3695 => x"82",
          3696 => x"ff",
          3697 => x"82",
          3698 => x"53",
          3699 => x"79",
          3700 => x"8e",
          3701 => x"79",
          3702 => x"ae",
          3703 => x"38",
          3704 => x"9f",
          3705 => x"fe",
          3706 => x"ff",
          3707 => x"e6",
          3708 => x"e0",
          3709 => x"2e",
          3710 => x"59",
          3711 => x"05",
          3712 => x"64",
          3713 => x"ff",
          3714 => x"c5",
          3715 => x"bc",
          3716 => x"a6",
          3717 => x"fe",
          3718 => x"ff",
          3719 => x"e0",
          3720 => x"e0",
          3721 => x"2e",
          3722 => x"b5",
          3723 => x"11",
          3724 => x"05",
          3725 => x"3f",
          3726 => x"08",
          3727 => x"38",
          3728 => x"80",
          3729 => x"79",
          3730 => x"5b",
          3731 => x"b5",
          3732 => x"11",
          3733 => x"05",
          3734 => x"3f",
          3735 => x"08",
          3736 => x"dd",
          3737 => x"22",
          3738 => x"c5",
          3739 => x"9f",
          3740 => x"fb",
          3741 => x"80",
          3742 => x"51",
          3743 => x"3f",
          3744 => x"33",
          3745 => x"2e",
          3746 => x"78",
          3747 => x"38",
          3748 => x"42",
          3749 => x"3d",
          3750 => x"53",
          3751 => x"51",
          3752 => x"82",
          3753 => x"80",
          3754 => x"61",
          3755 => x"c2",
          3756 => x"70",
          3757 => x"23",
          3758 => x"a9",
          3759 => x"d4",
          3760 => x"d4",
          3761 => x"39",
          3762 => x"f4",
          3763 => x"84",
          3764 => x"fb",
          3765 => x"98",
          3766 => x"f6",
          3767 => x"3d",
          3768 => x"53",
          3769 => x"51",
          3770 => x"82",
          3771 => x"80",
          3772 => x"61",
          3773 => x"59",
          3774 => x"42",
          3775 => x"f0",
          3776 => x"84",
          3777 => x"c7",
          3778 => x"98",
          3779 => x"f6",
          3780 => x"70",
          3781 => x"82",
          3782 => x"ff",
          3783 => x"82",
          3784 => x"53",
          3785 => x"79",
          3786 => x"b6",
          3787 => x"79",
          3788 => x"ae",
          3789 => x"38",
          3790 => x"9b",
          3791 => x"fe",
          3792 => x"ff",
          3793 => x"de",
          3794 => x"e0",
          3795 => x"2e",
          3796 => x"61",
          3797 => x"61",
          3798 => x"ff",
          3799 => x"c5",
          3800 => x"b9",
          3801 => x"aa",
          3802 => x"ff",
          3803 => x"ff",
          3804 => x"e3",
          3805 => x"e0",
          3806 => x"2e",
          3807 => x"64",
          3808 => x"f4",
          3809 => x"85",
          3810 => x"78",
          3811 => x"ff",
          3812 => x"ff",
          3813 => x"e3",
          3814 => x"e0",
          3815 => x"2e",
          3816 => x"64",
          3817 => x"90",
          3818 => x"e1",
          3819 => x"78",
          3820 => x"98",
          3821 => x"f5",
          3822 => x"e0",
          3823 => x"82",
          3824 => x"ff",
          3825 => x"f4",
          3826 => x"c6",
          3827 => x"b8",
          3828 => x"9c",
          3829 => x"e9",
          3830 => x"e4",
          3831 => x"b8",
          3832 => x"ff",
          3833 => x"ce",
          3834 => x"39",
          3835 => x"59",
          3836 => x"f4",
          3837 => x"f8",
          3838 => x"c9",
          3839 => x"e0",
          3840 => x"82",
          3841 => x"80",
          3842 => x"38",
          3843 => x"08",
          3844 => x"ff",
          3845 => x"83",
          3846 => x"e0",
          3847 => x"7f",
          3848 => x"78",
          3849 => x"d2",
          3850 => x"98",
          3851 => x"8a",
          3852 => x"98",
          3853 => x"81",
          3854 => x"5b",
          3855 => x"b2",
          3856 => x"24",
          3857 => x"81",
          3858 => x"80",
          3859 => x"83",
          3860 => x"80",
          3861 => x"c6",
          3862 => x"55",
          3863 => x"54",
          3864 => x"c7",
          3865 => x"3d",
          3866 => x"51",
          3867 => x"3f",
          3868 => x"52",
          3869 => x"b0",
          3870 => x"ac",
          3871 => x"7b",
          3872 => x"fc",
          3873 => x"82",
          3874 => x"b5",
          3875 => x"05",
          3876 => x"e1",
          3877 => x"7b",
          3878 => x"82",
          3879 => x"b5",
          3880 => x"05",
          3881 => x"cd",
          3882 => x"b4",
          3883 => x"c8",
          3884 => x"65",
          3885 => x"90",
          3886 => x"90",
          3887 => x"b5",
          3888 => x"05",
          3889 => x"3f",
          3890 => x"08",
          3891 => x"08",
          3892 => x"70",
          3893 => x"25",
          3894 => x"5f",
          3895 => x"83",
          3896 => x"81",
          3897 => x"06",
          3898 => x"2e",
          3899 => x"1b",
          3900 => x"06",
          3901 => x"fe",
          3902 => x"81",
          3903 => x"32",
          3904 => x"89",
          3905 => x"2e",
          3906 => x"89",
          3907 => x"a4",
          3908 => x"84",
          3909 => x"b1",
          3910 => x"a5",
          3911 => x"b4",
          3912 => x"f4",
          3913 => x"39",
          3914 => x"80",
          3915 => x"c8",
          3916 => x"94",
          3917 => x"54",
          3918 => x"80",
          3919 => x"cb",
          3920 => x"e0",
          3921 => x"2b",
          3922 => x"53",
          3923 => x"52",
          3924 => x"80",
          3925 => x"e0",
          3926 => x"75",
          3927 => x"94",
          3928 => x"54",
          3929 => x"80",
          3930 => x"ca",
          3931 => x"e0",
          3932 => x"2b",
          3933 => x"53",
          3934 => x"52",
          3935 => x"d4",
          3936 => x"e0",
          3937 => x"75",
          3938 => x"83",
          3939 => x"94",
          3940 => x"80",
          3941 => x"c0",
          3942 => x"81",
          3943 => x"81",
          3944 => x"83",
          3945 => x"99",
          3946 => x"5c",
          3947 => x"0b",
          3948 => x"88",
          3949 => x"72",
          3950 => x"fc",
          3951 => x"aa",
          3952 => x"3f",
          3953 => x"51",
          3954 => x"3f",
          3955 => x"51",
          3956 => x"3f",
          3957 => x"51",
          3958 => x"81",
          3959 => x"3f",
          3960 => x"80",
          3961 => x"0d",
          3962 => x"54",
          3963 => x"52",
          3964 => x"2e",
          3965 => x"72",
          3966 => x"a0",
          3967 => x"06",
          3968 => x"13",
          3969 => x"72",
          3970 => x"a2",
          3971 => x"06",
          3972 => x"13",
          3973 => x"72",
          3974 => x"2e",
          3975 => x"9f",
          3976 => x"81",
          3977 => x"72",
          3978 => x"70",
          3979 => x"38",
          3980 => x"80",
          3981 => x"73",
          3982 => x"39",
          3983 => x"80",
          3984 => x"54",
          3985 => x"83",
          3986 => x"70",
          3987 => x"38",
          3988 => x"80",
          3989 => x"54",
          3990 => x"09",
          3991 => x"38",
          3992 => x"a2",
          3993 => x"70",
          3994 => x"07",
          3995 => x"70",
          3996 => x"38",
          3997 => x"81",
          3998 => x"71",
          3999 => x"51",
          4000 => x"98",
          4001 => x"0d",
          4002 => x"0d",
          4003 => x"08",
          4004 => x"38",
          4005 => x"05",
          4006 => x"d7",
          4007 => x"e0",
          4008 => x"38",
          4009 => x"39",
          4010 => x"82",
          4011 => x"86",
          4012 => x"fc",
          4013 => x"82",
          4014 => x"05",
          4015 => x"52",
          4016 => x"81",
          4017 => x"13",
          4018 => x"51",
          4019 => x"9e",
          4020 => x"38",
          4021 => x"51",
          4022 => x"97",
          4023 => x"38",
          4024 => x"51",
          4025 => x"bb",
          4026 => x"38",
          4027 => x"51",
          4028 => x"bb",
          4029 => x"38",
          4030 => x"55",
          4031 => x"87",
          4032 => x"d9",
          4033 => x"22",
          4034 => x"73",
          4035 => x"80",
          4036 => x"0b",
          4037 => x"9c",
          4038 => x"87",
          4039 => x"0c",
          4040 => x"87",
          4041 => x"0c",
          4042 => x"87",
          4043 => x"0c",
          4044 => x"87",
          4045 => x"0c",
          4046 => x"87",
          4047 => x"0c",
          4048 => x"87",
          4049 => x"0c",
          4050 => x"98",
          4051 => x"87",
          4052 => x"0c",
          4053 => x"c0",
          4054 => x"80",
          4055 => x"e0",
          4056 => x"3d",
          4057 => x"3d",
          4058 => x"87",
          4059 => x"5d",
          4060 => x"87",
          4061 => x"08",
          4062 => x"23",
          4063 => x"b8",
          4064 => x"82",
          4065 => x"c0",
          4066 => x"5a",
          4067 => x"34",
          4068 => x"b0",
          4069 => x"84",
          4070 => x"c0",
          4071 => x"5a",
          4072 => x"34",
          4073 => x"a8",
          4074 => x"86",
          4075 => x"c0",
          4076 => x"5c",
          4077 => x"23",
          4078 => x"a0",
          4079 => x"8a",
          4080 => x"7d",
          4081 => x"ff",
          4082 => x"7b",
          4083 => x"06",
          4084 => x"33",
          4085 => x"33",
          4086 => x"33",
          4087 => x"33",
          4088 => x"33",
          4089 => x"ff",
          4090 => x"82",
          4091 => x"ff",
          4092 => x"8f",
          4093 => x"fd",
          4094 => x"97",
          4095 => x"80",
          4096 => x"2e",
          4097 => x"83",
          4098 => x"72",
          4099 => x"30",
          4100 => x"74",
          4101 => x"51",
          4102 => x"86",
          4103 => x"3f",
          4104 => x"f0",
          4105 => x"98",
          4106 => x"70",
          4107 => x"52",
          4108 => x"09",
          4109 => x"38",
          4110 => x"81",
          4111 => x"06",
          4112 => x"54",
          4113 => x"70",
          4114 => x"25",
          4115 => x"51",
          4116 => x"ab",
          4117 => x"e0",
          4118 => x"3d",
          4119 => x"3d",
          4120 => x"83",
          4121 => x"2b",
          4122 => x"ff",
          4123 => x"e0",
          4124 => x"2b",
          4125 => x"74",
          4126 => x"56",
          4127 => x"80",
          4128 => x"72",
          4129 => x"0c",
          4130 => x"04",
          4131 => x"02",
          4132 => x"82",
          4133 => x"70",
          4134 => x"58",
          4135 => x"c0",
          4136 => x"75",
          4137 => x"38",
          4138 => x"94",
          4139 => x"70",
          4140 => x"81",
          4141 => x"52",
          4142 => x"8c",
          4143 => x"2a",
          4144 => x"51",
          4145 => x"38",
          4146 => x"70",
          4147 => x"51",
          4148 => x"8d",
          4149 => x"2a",
          4150 => x"51",
          4151 => x"be",
          4152 => x"ff",
          4153 => x"c0",
          4154 => x"70",
          4155 => x"38",
          4156 => x"90",
          4157 => x"0c",
          4158 => x"98",
          4159 => x"0d",
          4160 => x"0d",
          4161 => x"33",
          4162 => x"9f",
          4163 => x"52",
          4164 => x"b0",
          4165 => x"0d",
          4166 => x"0d",
          4167 => x"33",
          4168 => x"2e",
          4169 => x"87",
          4170 => x"8d",
          4171 => x"82",
          4172 => x"70",
          4173 => x"58",
          4174 => x"94",
          4175 => x"80",
          4176 => x"87",
          4177 => x"53",
          4178 => x"96",
          4179 => x"06",
          4180 => x"72",
          4181 => x"38",
          4182 => x"70",
          4183 => x"53",
          4184 => x"74",
          4185 => x"81",
          4186 => x"72",
          4187 => x"38",
          4188 => x"70",
          4189 => x"53",
          4190 => x"38",
          4191 => x"06",
          4192 => x"94",
          4193 => x"80",
          4194 => x"87",
          4195 => x"54",
          4196 => x"80",
          4197 => x"98",
          4198 => x"0d",
          4199 => x"0d",
          4200 => x"74",
          4201 => x"ff",
          4202 => x"57",
          4203 => x"80",
          4204 => x"81",
          4205 => x"15",
          4206 => x"33",
          4207 => x"06",
          4208 => x"58",
          4209 => x"84",
          4210 => x"2e",
          4211 => x"c0",
          4212 => x"70",
          4213 => x"2a",
          4214 => x"53",
          4215 => x"80",
          4216 => x"71",
          4217 => x"81",
          4218 => x"70",
          4219 => x"81",
          4220 => x"06",
          4221 => x"80",
          4222 => x"71",
          4223 => x"81",
          4224 => x"70",
          4225 => x"74",
          4226 => x"51",
          4227 => x"80",
          4228 => x"2e",
          4229 => x"c0",
          4230 => x"77",
          4231 => x"17",
          4232 => x"81",
          4233 => x"53",
          4234 => x"86",
          4235 => x"e0",
          4236 => x"3d",
          4237 => x"3d",
          4238 => x"b0",
          4239 => x"ff",
          4240 => x"87",
          4241 => x"51",
          4242 => x"86",
          4243 => x"94",
          4244 => x"08",
          4245 => x"70",
          4246 => x"51",
          4247 => x"2e",
          4248 => x"81",
          4249 => x"87",
          4250 => x"52",
          4251 => x"86",
          4252 => x"94",
          4253 => x"08",
          4254 => x"06",
          4255 => x"0c",
          4256 => x"0d",
          4257 => x"3f",
          4258 => x"08",
          4259 => x"82",
          4260 => x"04",
          4261 => x"82",
          4262 => x"70",
          4263 => x"52",
          4264 => x"94",
          4265 => x"80",
          4266 => x"87",
          4267 => x"52",
          4268 => x"82",
          4269 => x"06",
          4270 => x"ff",
          4271 => x"2e",
          4272 => x"81",
          4273 => x"87",
          4274 => x"52",
          4275 => x"86",
          4276 => x"94",
          4277 => x"08",
          4278 => x"70",
          4279 => x"53",
          4280 => x"e0",
          4281 => x"3d",
          4282 => x"3d",
          4283 => x"9e",
          4284 => x"9c",
          4285 => x"51",
          4286 => x"2e",
          4287 => x"87",
          4288 => x"08",
          4289 => x"0c",
          4290 => x"a8",
          4291 => x"b8",
          4292 => x"9e",
          4293 => x"de",
          4294 => x"c0",
          4295 => x"82",
          4296 => x"87",
          4297 => x"08",
          4298 => x"0c",
          4299 => x"a0",
          4300 => x"c8",
          4301 => x"9e",
          4302 => x"de",
          4303 => x"c0",
          4304 => x"82",
          4305 => x"87",
          4306 => x"08",
          4307 => x"0c",
          4308 => x"b8",
          4309 => x"d8",
          4310 => x"9e",
          4311 => x"de",
          4312 => x"c0",
          4313 => x"82",
          4314 => x"87",
          4315 => x"08",
          4316 => x"0c",
          4317 => x"80",
          4318 => x"82",
          4319 => x"87",
          4320 => x"08",
          4321 => x"0c",
          4322 => x"88",
          4323 => x"f0",
          4324 => x"9e",
          4325 => x"de",
          4326 => x"0b",
          4327 => x"34",
          4328 => x"c0",
          4329 => x"70",
          4330 => x"06",
          4331 => x"70",
          4332 => x"38",
          4333 => x"82",
          4334 => x"80",
          4335 => x"9e",
          4336 => x"88",
          4337 => x"51",
          4338 => x"80",
          4339 => x"81",
          4340 => x"de",
          4341 => x"0b",
          4342 => x"90",
          4343 => x"80",
          4344 => x"52",
          4345 => x"2e",
          4346 => x"52",
          4347 => x"fb",
          4348 => x"87",
          4349 => x"08",
          4350 => x"80",
          4351 => x"52",
          4352 => x"83",
          4353 => x"71",
          4354 => x"34",
          4355 => x"c0",
          4356 => x"70",
          4357 => x"06",
          4358 => x"70",
          4359 => x"38",
          4360 => x"82",
          4361 => x"80",
          4362 => x"9e",
          4363 => x"90",
          4364 => x"51",
          4365 => x"80",
          4366 => x"81",
          4367 => x"de",
          4368 => x"0b",
          4369 => x"90",
          4370 => x"80",
          4371 => x"52",
          4372 => x"2e",
          4373 => x"52",
          4374 => x"ff",
          4375 => x"87",
          4376 => x"08",
          4377 => x"80",
          4378 => x"52",
          4379 => x"83",
          4380 => x"71",
          4381 => x"34",
          4382 => x"c0",
          4383 => x"70",
          4384 => x"06",
          4385 => x"70",
          4386 => x"38",
          4387 => x"82",
          4388 => x"80",
          4389 => x"9e",
          4390 => x"80",
          4391 => x"51",
          4392 => x"80",
          4393 => x"81",
          4394 => x"df",
          4395 => x"0b",
          4396 => x"90",
          4397 => x"80",
          4398 => x"52",
          4399 => x"83",
          4400 => x"71",
          4401 => x"34",
          4402 => x"90",
          4403 => x"80",
          4404 => x"2a",
          4405 => x"70",
          4406 => x"34",
          4407 => x"c0",
          4408 => x"70",
          4409 => x"51",
          4410 => x"80",
          4411 => x"81",
          4412 => x"df",
          4413 => x"c0",
          4414 => x"70",
          4415 => x"70",
          4416 => x"51",
          4417 => x"df",
          4418 => x"0b",
          4419 => x"90",
          4420 => x"06",
          4421 => x"70",
          4422 => x"38",
          4423 => x"82",
          4424 => x"87",
          4425 => x"08",
          4426 => x"51",
          4427 => x"df",
          4428 => x"3d",
          4429 => x"3d",
          4430 => x"9c",
          4431 => x"cd",
          4432 => x"f8",
          4433 => x"80",
          4434 => x"82",
          4435 => x"ff",
          4436 => x"82",
          4437 => x"ff",
          4438 => x"82",
          4439 => x"54",
          4440 => x"94",
          4441 => x"d4",
          4442 => x"d8",
          4443 => x"52",
          4444 => x"51",
          4445 => x"3f",
          4446 => x"33",
          4447 => x"2e",
          4448 => x"de",
          4449 => x"de",
          4450 => x"54",
          4451 => x"f8",
          4452 => x"f9",
          4453 => x"fc",
          4454 => x"80",
          4455 => x"82",
          4456 => x"82",
          4457 => x"11",
          4458 => x"c9",
          4459 => x"88",
          4460 => x"de",
          4461 => x"73",
          4462 => x"38",
          4463 => x"08",
          4464 => x"08",
          4465 => x"82",
          4466 => x"ff",
          4467 => x"82",
          4468 => x"54",
          4469 => x"94",
          4470 => x"c4",
          4471 => x"c8",
          4472 => x"52",
          4473 => x"51",
          4474 => x"3f",
          4475 => x"33",
          4476 => x"2e",
          4477 => x"df",
          4478 => x"82",
          4479 => x"ff",
          4480 => x"82",
          4481 => x"54",
          4482 => x"8e",
          4483 => x"88",
          4484 => x"ca",
          4485 => x"87",
          4486 => x"df",
          4487 => x"73",
          4488 => x"38",
          4489 => x"33",
          4490 => x"a8",
          4491 => x"dd",
          4492 => x"f9",
          4493 => x"80",
          4494 => x"82",
          4495 => x"ff",
          4496 => x"82",
          4497 => x"54",
          4498 => x"89",
          4499 => x"dc",
          4500 => x"c4",
          4501 => x"80",
          4502 => x"80",
          4503 => x"82",
          4504 => x"ff",
          4505 => x"82",
          4506 => x"54",
          4507 => x"89",
          4508 => x"f4",
          4509 => x"a0",
          4510 => x"82",
          4511 => x"80",
          4512 => x"82",
          4513 => x"ff",
          4514 => x"82",
          4515 => x"ff",
          4516 => x"82",
          4517 => x"52",
          4518 => x"51",
          4519 => x"3f",
          4520 => x"08",
          4521 => x"b8",
          4522 => x"e1",
          4523 => x"e4",
          4524 => x"cb",
          4525 => x"86",
          4526 => x"cc",
          4527 => x"a2",
          4528 => x"de",
          4529 => x"82",
          4530 => x"ff",
          4531 => x"82",
          4532 => x"56",
          4533 => x"52",
          4534 => x"b7",
          4535 => x"e0",
          4536 => x"84",
          4537 => x"71",
          4538 => x"82",
          4539 => x"52",
          4540 => x"51",
          4541 => x"3f",
          4542 => x"33",
          4543 => x"2e",
          4544 => x"de",
          4545 => x"bd",
          4546 => x"75",
          4547 => x"c4",
          4548 => x"98",
          4549 => x"c0",
          4550 => x"31",
          4551 => x"e0",
          4552 => x"82",
          4553 => x"ff",
          4554 => x"82",
          4555 => x"54",
          4556 => x"aa",
          4557 => x"f4",
          4558 => x"84",
          4559 => x"51",
          4560 => x"3f",
          4561 => x"08",
          4562 => x"29",
          4563 => x"54",
          4564 => x"98",
          4565 => x"cd",
          4566 => x"85",
          4567 => x"51",
          4568 => x"3f",
          4569 => x"04",
          4570 => x"02",
          4571 => x"ff",
          4572 => x"84",
          4573 => x"71",
          4574 => x"b8",
          4575 => x"71",
          4576 => x"cd",
          4577 => x"39",
          4578 => x"51",
          4579 => x"cd",
          4580 => x"39",
          4581 => x"51",
          4582 => x"cd",
          4583 => x"39",
          4584 => x"51",
          4585 => x"3f",
          4586 => x"04",
          4587 => x"0c",
          4588 => x"87",
          4589 => x"0c",
          4590 => x"8c",
          4591 => x"96",
          4592 => x"fd",
          4593 => x"98",
          4594 => x"2c",
          4595 => x"70",
          4596 => x"10",
          4597 => x"2b",
          4598 => x"54",
          4599 => x"0b",
          4600 => x"12",
          4601 => x"71",
          4602 => x"38",
          4603 => x"11",
          4604 => x"84",
          4605 => x"33",
          4606 => x"52",
          4607 => x"2e",
          4608 => x"83",
          4609 => x"72",
          4610 => x"0c",
          4611 => x"04",
          4612 => x"79",
          4613 => x"a3",
          4614 => x"33",
          4615 => x"72",
          4616 => x"38",
          4617 => x"08",
          4618 => x"ff",
          4619 => x"82",
          4620 => x"52",
          4621 => x"a3",
          4622 => x"fb",
          4623 => x"88",
          4624 => x"a3",
          4625 => x"ff",
          4626 => x"74",
          4627 => x"ff",
          4628 => x"39",
          4629 => x"83",
          4630 => x"74",
          4631 => x"0d",
          4632 => x"0d",
          4633 => x"05",
          4634 => x"02",
          4635 => x"05",
          4636 => x"e8",
          4637 => x"29",
          4638 => x"05",
          4639 => x"59",
          4640 => x"59",
          4641 => x"86",
          4642 => x"9a",
          4643 => x"df",
          4644 => x"84",
          4645 => x"90",
          4646 => x"70",
          4647 => x"5a",
          4648 => x"82",
          4649 => x"75",
          4650 => x"e8",
          4651 => x"29",
          4652 => x"05",
          4653 => x"56",
          4654 => x"2e",
          4655 => x"53",
          4656 => x"51",
          4657 => x"3f",
          4658 => x"33",
          4659 => x"74",
          4660 => x"34",
          4661 => x"06",
          4662 => x"27",
          4663 => x"0b",
          4664 => x"34",
          4665 => x"b6",
          4666 => x"e4",
          4667 => x"80",
          4668 => x"82",
          4669 => x"55",
          4670 => x"8c",
          4671 => x"54",
          4672 => x"52",
          4673 => x"ec",
          4674 => x"df",
          4675 => x"8a",
          4676 => x"d6",
          4677 => x"e4",
          4678 => x"ef",
          4679 => x"3d",
          4680 => x"3d",
          4681 => x"90",
          4682 => x"72",
          4683 => x"80",
          4684 => x"71",
          4685 => x"3f",
          4686 => x"ff",
          4687 => x"54",
          4688 => x"25",
          4689 => x"0b",
          4690 => x"34",
          4691 => x"08",
          4692 => x"2e",
          4693 => x"51",
          4694 => x"3f",
          4695 => x"08",
          4696 => x"3f",
          4697 => x"df",
          4698 => x"3d",
          4699 => x"3d",
          4700 => x"80",
          4701 => x"e4",
          4702 => x"f5",
          4703 => x"e0",
          4704 => x"d3",
          4705 => x"e4",
          4706 => x"f8",
          4707 => x"70",
          4708 => x"9f",
          4709 => x"e0",
          4710 => x"2e",
          4711 => x"51",
          4712 => x"3f",
          4713 => x"08",
          4714 => x"82",
          4715 => x"25",
          4716 => x"e0",
          4717 => x"05",
          4718 => x"55",
          4719 => x"75",
          4720 => x"81",
          4721 => x"dc",
          4722 => x"80",
          4723 => x"ff",
          4724 => x"06",
          4725 => x"a6",
          4726 => x"d9",
          4727 => x"3d",
          4728 => x"08",
          4729 => x"70",
          4730 => x"52",
          4731 => x"08",
          4732 => x"f2",
          4733 => x"98",
          4734 => x"38",
          4735 => x"df",
          4736 => x"55",
          4737 => x"8b",
          4738 => x"56",
          4739 => x"3f",
          4740 => x"08",
          4741 => x"38",
          4742 => x"a8",
          4743 => x"e0",
          4744 => x"18",
          4745 => x"0b",
          4746 => x"08",
          4747 => x"82",
          4748 => x"ff",
          4749 => x"55",
          4750 => x"34",
          4751 => x"30",
          4752 => x"9f",
          4753 => x"55",
          4754 => x"85",
          4755 => x"ac",
          4756 => x"e4",
          4757 => x"08",
          4758 => x"f4",
          4759 => x"e0",
          4760 => x"2e",
          4761 => x"d0",
          4762 => x"ff",
          4763 => x"77",
          4764 => x"06",
          4765 => x"52",
          4766 => x"a8",
          4767 => x"51",
          4768 => x"3f",
          4769 => x"54",
          4770 => x"08",
          4771 => x"58",
          4772 => x"98",
          4773 => x"0d",
          4774 => x"0d",
          4775 => x"5c",
          4776 => x"57",
          4777 => x"73",
          4778 => x"81",
          4779 => x"78",
          4780 => x"56",
          4781 => x"98",
          4782 => x"70",
          4783 => x"33",
          4784 => x"73",
          4785 => x"81",
          4786 => x"75",
          4787 => x"38",
          4788 => x"88",
          4789 => x"ec",
          4790 => x"52",
          4791 => x"da",
          4792 => x"98",
          4793 => x"52",
          4794 => x"ff",
          4795 => x"82",
          4796 => x"80",
          4797 => x"15",
          4798 => x"81",
          4799 => x"74",
          4800 => x"38",
          4801 => x"e6",
          4802 => x"81",
          4803 => x"3d",
          4804 => x"f8",
          4805 => x"88",
          4806 => x"98",
          4807 => x"9a",
          4808 => x"53",
          4809 => x"51",
          4810 => x"82",
          4811 => x"81",
          4812 => x"74",
          4813 => x"54",
          4814 => x"14",
          4815 => x"06",
          4816 => x"74",
          4817 => x"38",
          4818 => x"82",
          4819 => x"8c",
          4820 => x"d3",
          4821 => x"3d",
          4822 => x"08",
          4823 => x"59",
          4824 => x"0b",
          4825 => x"82",
          4826 => x"82",
          4827 => x"55",
          4828 => x"cb",
          4829 => x"df",
          4830 => x"55",
          4831 => x"81",
          4832 => x"2e",
          4833 => x"81",
          4834 => x"55",
          4835 => x"2e",
          4836 => x"a8",
          4837 => x"3f",
          4838 => x"08",
          4839 => x"0c",
          4840 => x"08",
          4841 => x"92",
          4842 => x"76",
          4843 => x"98",
          4844 => x"de",
          4845 => x"e0",
          4846 => x"2e",
          4847 => x"d1",
          4848 => x"98",
          4849 => x"f7",
          4850 => x"98",
          4851 => x"df",
          4852 => x"80",
          4853 => x"3d",
          4854 => x"81",
          4855 => x"82",
          4856 => x"56",
          4857 => x"08",
          4858 => x"81",
          4859 => x"38",
          4860 => x"08",
          4861 => x"c2",
          4862 => x"98",
          4863 => x"0b",
          4864 => x"08",
          4865 => x"82",
          4866 => x"ff",
          4867 => x"55",
          4868 => x"34",
          4869 => x"81",
          4870 => x"75",
          4871 => x"3f",
          4872 => x"81",
          4873 => x"54",
          4874 => x"83",
          4875 => x"74",
          4876 => x"81",
          4877 => x"38",
          4878 => x"82",
          4879 => x"76",
          4880 => x"df",
          4881 => x"2e",
          4882 => x"d6",
          4883 => x"5d",
          4884 => x"a3",
          4885 => x"98",
          4886 => x"70",
          4887 => x"59",
          4888 => x"ec",
          4889 => x"ff",
          4890 => x"d4",
          4891 => x"2b",
          4892 => x"82",
          4893 => x"70",
          4894 => x"97",
          4895 => x"2c",
          4896 => x"29",
          4897 => x"05",
          4898 => x"70",
          4899 => x"51",
          4900 => x"51",
          4901 => x"81",
          4902 => x"2e",
          4903 => x"77",
          4904 => x"38",
          4905 => x"0a",
          4906 => x"0a",
          4907 => x"2c",
          4908 => x"75",
          4909 => x"38",
          4910 => x"52",
          4911 => x"83",
          4912 => x"98",
          4913 => x"06",
          4914 => x"2e",
          4915 => x"82",
          4916 => x"81",
          4917 => x"74",
          4918 => x"29",
          4919 => x"05",
          4920 => x"70",
          4921 => x"56",
          4922 => x"95",
          4923 => x"76",
          4924 => x"77",
          4925 => x"3f",
          4926 => x"08",
          4927 => x"54",
          4928 => x"d3",
          4929 => x"75",
          4930 => x"ca",
          4931 => x"55",
          4932 => x"d4",
          4933 => x"2b",
          4934 => x"82",
          4935 => x"70",
          4936 => x"98",
          4937 => x"11",
          4938 => x"82",
          4939 => x"33",
          4940 => x"51",
          4941 => x"55",
          4942 => x"09",
          4943 => x"90",
          4944 => x"f0",
          4945 => x"0c",
          4946 => x"f7",
          4947 => x"0b",
          4948 => x"34",
          4949 => x"82",
          4950 => x"75",
          4951 => x"34",
          4952 => x"34",
          4953 => x"7e",
          4954 => x"26",
          4955 => x"73",
          4956 => x"b8",
          4957 => x"73",
          4958 => x"f7",
          4959 => x"73",
          4960 => x"c9",
          4961 => x"d8",
          4962 => x"75",
          4963 => x"74",
          4964 => x"98",
          4965 => x"73",
          4966 => x"38",
          4967 => x"73",
          4968 => x"34",
          4969 => x"0a",
          4970 => x"0a",
          4971 => x"2c",
          4972 => x"33",
          4973 => x"df",
          4974 => x"dc",
          4975 => x"56",
          4976 => x"f7",
          4977 => x"1a",
          4978 => x"33",
          4979 => x"f7",
          4980 => x"73",
          4981 => x"38",
          4982 => x"73",
          4983 => x"34",
          4984 => x"33",
          4985 => x"0a",
          4986 => x"0a",
          4987 => x"2c",
          4988 => x"33",
          4989 => x"56",
          4990 => x"a8",
          4991 => x"fc",
          4992 => x"1a",
          4993 => x"54",
          4994 => x"3f",
          4995 => x"0a",
          4996 => x"0a",
          4997 => x"2c",
          4998 => x"33",
          4999 => x"73",
          5000 => x"38",
          5001 => x"33",
          5002 => x"70",
          5003 => x"f7",
          5004 => x"51",
          5005 => x"77",
          5006 => x"38",
          5007 => x"08",
          5008 => x"ff",
          5009 => x"74",
          5010 => x"29",
          5011 => x"05",
          5012 => x"82",
          5013 => x"56",
          5014 => x"75",
          5015 => x"fb",
          5016 => x"7a",
          5017 => x"81",
          5018 => x"f7",
          5019 => x"52",
          5020 => x"51",
          5021 => x"81",
          5022 => x"f7",
          5023 => x"81",
          5024 => x"55",
          5025 => x"fb",
          5026 => x"f7",
          5027 => x"05",
          5028 => x"f7",
          5029 => x"15",
          5030 => x"f7",
          5031 => x"fb",
          5032 => x"88",
          5033 => x"bf",
          5034 => x"dc",
          5035 => x"2b",
          5036 => x"82",
          5037 => x"57",
          5038 => x"74",
          5039 => x"38",
          5040 => x"81",
          5041 => x"34",
          5042 => x"08",
          5043 => x"51",
          5044 => x"3f",
          5045 => x"0a",
          5046 => x"0a",
          5047 => x"2c",
          5048 => x"33",
          5049 => x"75",
          5050 => x"38",
          5051 => x"08",
          5052 => x"ff",
          5053 => x"82",
          5054 => x"70",
          5055 => x"98",
          5056 => x"d8",
          5057 => x"56",
          5058 => x"24",
          5059 => x"82",
          5060 => x"52",
          5061 => x"95",
          5062 => x"81",
          5063 => x"81",
          5064 => x"70",
          5065 => x"f7",
          5066 => x"51",
          5067 => x"25",
          5068 => x"99",
          5069 => x"d8",
          5070 => x"54",
          5071 => x"82",
          5072 => x"52",
          5073 => x"95",
          5074 => x"f7",
          5075 => x"51",
          5076 => x"82",
          5077 => x"81",
          5078 => x"73",
          5079 => x"f7",
          5080 => x"73",
          5081 => x"38",
          5082 => x"52",
          5083 => x"f1",
          5084 => x"80",
          5085 => x"0b",
          5086 => x"34",
          5087 => x"f7",
          5088 => x"82",
          5089 => x"af",
          5090 => x"82",
          5091 => x"54",
          5092 => x"f9",
          5093 => x"fb",
          5094 => x"88",
          5095 => x"c7",
          5096 => x"dc",
          5097 => x"54",
          5098 => x"dc",
          5099 => x"ff",
          5100 => x"39",
          5101 => x"33",
          5102 => x"33",
          5103 => x"75",
          5104 => x"38",
          5105 => x"73",
          5106 => x"34",
          5107 => x"70",
          5108 => x"81",
          5109 => x"51",
          5110 => x"25",
          5111 => x"1a",
          5112 => x"33",
          5113 => x"fb",
          5114 => x"73",
          5115 => x"93",
          5116 => x"81",
          5117 => x"81",
          5118 => x"70",
          5119 => x"f7",
          5120 => x"51",
          5121 => x"24",
          5122 => x"fb",
          5123 => x"a0",
          5124 => x"d3",
          5125 => x"dc",
          5126 => x"2b",
          5127 => x"82",
          5128 => x"57",
          5129 => x"74",
          5130 => x"a1",
          5131 => x"fc",
          5132 => x"51",
          5133 => x"3f",
          5134 => x"0a",
          5135 => x"0a",
          5136 => x"2c",
          5137 => x"33",
          5138 => x"75",
          5139 => x"38",
          5140 => x"82",
          5141 => x"70",
          5142 => x"82",
          5143 => x"59",
          5144 => x"77",
          5145 => x"38",
          5146 => x"08",
          5147 => x"54",
          5148 => x"dc",
          5149 => x"70",
          5150 => x"ff",
          5151 => x"82",
          5152 => x"70",
          5153 => x"82",
          5154 => x"58",
          5155 => x"75",
          5156 => x"f7",
          5157 => x"f7",
          5158 => x"52",
          5159 => x"51",
          5160 => x"80",
          5161 => x"dc",
          5162 => x"82",
          5163 => x"f7",
          5164 => x"b0",
          5165 => x"dc",
          5166 => x"80",
          5167 => x"74",
          5168 => x"f6",
          5169 => x"98",
          5170 => x"d8",
          5171 => x"98",
          5172 => x"06",
          5173 => x"74",
          5174 => x"ff",
          5175 => x"93",
          5176 => x"39",
          5177 => x"82",
          5178 => x"fc",
          5179 => x"54",
          5180 => x"a7",
          5181 => x"ff",
          5182 => x"82",
          5183 => x"82",
          5184 => x"82",
          5185 => x"81",
          5186 => x"05",
          5187 => x"79",
          5188 => x"86",
          5189 => x"54",
          5190 => x"73",
          5191 => x"80",
          5192 => x"38",
          5193 => x"9a",
          5194 => x"39",
          5195 => x"09",
          5196 => x"38",
          5197 => x"08",
          5198 => x"2e",
          5199 => x"51",
          5200 => x"3f",
          5201 => x"08",
          5202 => x"34",
          5203 => x"08",
          5204 => x"81",
          5205 => x"52",
          5206 => x"9b",
          5207 => x"c3",
          5208 => x"29",
          5209 => x"05",
          5210 => x"54",
          5211 => x"ab",
          5212 => x"ff",
          5213 => x"82",
          5214 => x"82",
          5215 => x"82",
          5216 => x"81",
          5217 => x"05",
          5218 => x"79",
          5219 => x"8a",
          5220 => x"54",
          5221 => x"06",
          5222 => x"74",
          5223 => x"34",
          5224 => x"82",
          5225 => x"82",
          5226 => x"52",
          5227 => x"e0",
          5228 => x"39",
          5229 => x"33",
          5230 => x"06",
          5231 => x"33",
          5232 => x"74",
          5233 => x"85",
          5234 => x"fc",
          5235 => x"14",
          5236 => x"f7",
          5237 => x"1a",
          5238 => x"54",
          5239 => x"3f",
          5240 => x"82",
          5241 => x"54",
          5242 => x"f4",
          5243 => x"fb",
          5244 => x"88",
          5245 => x"ef",
          5246 => x"dc",
          5247 => x"54",
          5248 => x"dc",
          5249 => x"39",
          5250 => x"84",
          5251 => x"82",
          5252 => x"a0",
          5253 => x"e0",
          5254 => x"80",
          5255 => x"52",
          5256 => x"51",
          5257 => x"3f",
          5258 => x"08",
          5259 => x"77",
          5260 => x"57",
          5261 => x"34",
          5262 => x"08",
          5263 => x"15",
          5264 => x"15",
          5265 => x"88",
          5266 => x"86",
          5267 => x"87",
          5268 => x"e0",
          5269 => x"e0",
          5270 => x"05",
          5271 => x"07",
          5272 => x"ff",
          5273 => x"2a",
          5274 => x"56",
          5275 => x"34",
          5276 => x"34",
          5277 => x"22",
          5278 => x"82",
          5279 => x"05",
          5280 => x"55",
          5281 => x"15",
          5282 => x"15",
          5283 => x"0d",
          5284 => x"0d",
          5285 => x"51",
          5286 => x"8f",
          5287 => x"83",
          5288 => x"70",
          5289 => x"06",
          5290 => x"70",
          5291 => x"0c",
          5292 => x"04",
          5293 => x"02",
          5294 => x"02",
          5295 => x"05",
          5296 => x"82",
          5297 => x"71",
          5298 => x"11",
          5299 => x"73",
          5300 => x"81",
          5301 => x"88",
          5302 => x"a4",
          5303 => x"22",
          5304 => x"ff",
          5305 => x"88",
          5306 => x"52",
          5307 => x"5b",
          5308 => x"55",
          5309 => x"70",
          5310 => x"82",
          5311 => x"14",
          5312 => x"52",
          5313 => x"15",
          5314 => x"15",
          5315 => x"88",
          5316 => x"70",
          5317 => x"33",
          5318 => x"07",
          5319 => x"8f",
          5320 => x"51",
          5321 => x"71",
          5322 => x"ff",
          5323 => x"88",
          5324 => x"51",
          5325 => x"34",
          5326 => x"06",
          5327 => x"12",
          5328 => x"88",
          5329 => x"71",
          5330 => x"81",
          5331 => x"3d",
          5332 => x"3d",
          5333 => x"88",
          5334 => x"05",
          5335 => x"70",
          5336 => x"11",
          5337 => x"87",
          5338 => x"8b",
          5339 => x"2b",
          5340 => x"59",
          5341 => x"72",
          5342 => x"33",
          5343 => x"71",
          5344 => x"70",
          5345 => x"56",
          5346 => x"84",
          5347 => x"85",
          5348 => x"e0",
          5349 => x"14",
          5350 => x"85",
          5351 => x"8b",
          5352 => x"2b",
          5353 => x"57",
          5354 => x"86",
          5355 => x"13",
          5356 => x"2b",
          5357 => x"2a",
          5358 => x"52",
          5359 => x"34",
          5360 => x"34",
          5361 => x"08",
          5362 => x"81",
          5363 => x"88",
          5364 => x"81",
          5365 => x"70",
          5366 => x"51",
          5367 => x"71",
          5368 => x"81",
          5369 => x"3d",
          5370 => x"3d",
          5371 => x"05",
          5372 => x"88",
          5373 => x"2b",
          5374 => x"33",
          5375 => x"71",
          5376 => x"70",
          5377 => x"70",
          5378 => x"33",
          5379 => x"71",
          5380 => x"53",
          5381 => x"52",
          5382 => x"53",
          5383 => x"25",
          5384 => x"72",
          5385 => x"3f",
          5386 => x"08",
          5387 => x"33",
          5388 => x"71",
          5389 => x"83",
          5390 => x"11",
          5391 => x"12",
          5392 => x"2b",
          5393 => x"2b",
          5394 => x"06",
          5395 => x"51",
          5396 => x"53",
          5397 => x"88",
          5398 => x"72",
          5399 => x"73",
          5400 => x"82",
          5401 => x"70",
          5402 => x"81",
          5403 => x"8b",
          5404 => x"2b",
          5405 => x"57",
          5406 => x"70",
          5407 => x"33",
          5408 => x"07",
          5409 => x"ff",
          5410 => x"2a",
          5411 => x"58",
          5412 => x"34",
          5413 => x"34",
          5414 => x"04",
          5415 => x"82",
          5416 => x"02",
          5417 => x"05",
          5418 => x"2b",
          5419 => x"11",
          5420 => x"33",
          5421 => x"71",
          5422 => x"59",
          5423 => x"56",
          5424 => x"71",
          5425 => x"33",
          5426 => x"07",
          5427 => x"a2",
          5428 => x"07",
          5429 => x"53",
          5430 => x"53",
          5431 => x"70",
          5432 => x"82",
          5433 => x"70",
          5434 => x"81",
          5435 => x"8b",
          5436 => x"2b",
          5437 => x"57",
          5438 => x"82",
          5439 => x"13",
          5440 => x"2b",
          5441 => x"2a",
          5442 => x"52",
          5443 => x"34",
          5444 => x"34",
          5445 => x"08",
          5446 => x"33",
          5447 => x"71",
          5448 => x"82",
          5449 => x"52",
          5450 => x"0d",
          5451 => x"0d",
          5452 => x"88",
          5453 => x"2a",
          5454 => x"ff",
          5455 => x"57",
          5456 => x"3f",
          5457 => x"08",
          5458 => x"71",
          5459 => x"33",
          5460 => x"71",
          5461 => x"83",
          5462 => x"11",
          5463 => x"12",
          5464 => x"2b",
          5465 => x"07",
          5466 => x"51",
          5467 => x"55",
          5468 => x"80",
          5469 => x"82",
          5470 => x"75",
          5471 => x"3f",
          5472 => x"84",
          5473 => x"15",
          5474 => x"2b",
          5475 => x"07",
          5476 => x"88",
          5477 => x"55",
          5478 => x"86",
          5479 => x"81",
          5480 => x"75",
          5481 => x"82",
          5482 => x"70",
          5483 => x"33",
          5484 => x"71",
          5485 => x"70",
          5486 => x"57",
          5487 => x"72",
          5488 => x"73",
          5489 => x"82",
          5490 => x"18",
          5491 => x"86",
          5492 => x"0b",
          5493 => x"82",
          5494 => x"53",
          5495 => x"34",
          5496 => x"34",
          5497 => x"08",
          5498 => x"81",
          5499 => x"88",
          5500 => x"82",
          5501 => x"70",
          5502 => x"51",
          5503 => x"74",
          5504 => x"81",
          5505 => x"3d",
          5506 => x"3d",
          5507 => x"82",
          5508 => x"84",
          5509 => x"3f",
          5510 => x"86",
          5511 => x"fe",
          5512 => x"3d",
          5513 => x"3d",
          5514 => x"52",
          5515 => x"3f",
          5516 => x"08",
          5517 => x"06",
          5518 => x"08",
          5519 => x"85",
          5520 => x"88",
          5521 => x"5f",
          5522 => x"5a",
          5523 => x"59",
          5524 => x"80",
          5525 => x"88",
          5526 => x"33",
          5527 => x"71",
          5528 => x"70",
          5529 => x"06",
          5530 => x"83",
          5531 => x"70",
          5532 => x"53",
          5533 => x"55",
          5534 => x"8a",
          5535 => x"2e",
          5536 => x"78",
          5537 => x"15",
          5538 => x"33",
          5539 => x"07",
          5540 => x"c2",
          5541 => x"ff",
          5542 => x"38",
          5543 => x"56",
          5544 => x"2b",
          5545 => x"08",
          5546 => x"81",
          5547 => x"88",
          5548 => x"81",
          5549 => x"51",
          5550 => x"5c",
          5551 => x"2e",
          5552 => x"55",
          5553 => x"78",
          5554 => x"38",
          5555 => x"80",
          5556 => x"38",
          5557 => x"09",
          5558 => x"38",
          5559 => x"f2",
          5560 => x"39",
          5561 => x"53",
          5562 => x"51",
          5563 => x"82",
          5564 => x"70",
          5565 => x"33",
          5566 => x"71",
          5567 => x"83",
          5568 => x"5a",
          5569 => x"05",
          5570 => x"83",
          5571 => x"70",
          5572 => x"59",
          5573 => x"84",
          5574 => x"81",
          5575 => x"76",
          5576 => x"82",
          5577 => x"75",
          5578 => x"11",
          5579 => x"11",
          5580 => x"33",
          5581 => x"07",
          5582 => x"53",
          5583 => x"5a",
          5584 => x"86",
          5585 => x"87",
          5586 => x"e0",
          5587 => x"1c",
          5588 => x"85",
          5589 => x"8b",
          5590 => x"2b",
          5591 => x"5a",
          5592 => x"54",
          5593 => x"34",
          5594 => x"34",
          5595 => x"08",
          5596 => x"1d",
          5597 => x"85",
          5598 => x"88",
          5599 => x"88",
          5600 => x"5f",
          5601 => x"73",
          5602 => x"75",
          5603 => x"82",
          5604 => x"1b",
          5605 => x"73",
          5606 => x"0c",
          5607 => x"04",
          5608 => x"74",
          5609 => x"88",
          5610 => x"f4",
          5611 => x"53",
          5612 => x"8b",
          5613 => x"fc",
          5614 => x"e0",
          5615 => x"72",
          5616 => x"0c",
          5617 => x"04",
          5618 => x"64",
          5619 => x"80",
          5620 => x"82",
          5621 => x"60",
          5622 => x"06",
          5623 => x"a8",
          5624 => x"38",
          5625 => x"b8",
          5626 => x"98",
          5627 => x"c7",
          5628 => x"38",
          5629 => x"92",
          5630 => x"83",
          5631 => x"51",
          5632 => x"82",
          5633 => x"83",
          5634 => x"82",
          5635 => x"7d",
          5636 => x"2a",
          5637 => x"ff",
          5638 => x"2b",
          5639 => x"33",
          5640 => x"71",
          5641 => x"70",
          5642 => x"83",
          5643 => x"70",
          5644 => x"05",
          5645 => x"1a",
          5646 => x"12",
          5647 => x"2b",
          5648 => x"2b",
          5649 => x"53",
          5650 => x"5c",
          5651 => x"5c",
          5652 => x"73",
          5653 => x"38",
          5654 => x"ff",
          5655 => x"70",
          5656 => x"06",
          5657 => x"16",
          5658 => x"33",
          5659 => x"07",
          5660 => x"1c",
          5661 => x"12",
          5662 => x"2b",
          5663 => x"07",
          5664 => x"52",
          5665 => x"80",
          5666 => x"78",
          5667 => x"83",
          5668 => x"41",
          5669 => x"27",
          5670 => x"60",
          5671 => x"7b",
          5672 => x"06",
          5673 => x"51",
          5674 => x"7a",
          5675 => x"06",
          5676 => x"39",
          5677 => x"7a",
          5678 => x"38",
          5679 => x"aa",
          5680 => x"39",
          5681 => x"7a",
          5682 => x"c8",
          5683 => x"82",
          5684 => x"12",
          5685 => x"2b",
          5686 => x"54",
          5687 => x"80",
          5688 => x"f7",
          5689 => x"e0",
          5690 => x"ff",
          5691 => x"54",
          5692 => x"83",
          5693 => x"88",
          5694 => x"05",
          5695 => x"ff",
          5696 => x"82",
          5697 => x"14",
          5698 => x"83",
          5699 => x"59",
          5700 => x"39",
          5701 => x"7a",
          5702 => x"d4",
          5703 => x"f5",
          5704 => x"e0",
          5705 => x"82",
          5706 => x"12",
          5707 => x"2b",
          5708 => x"54",
          5709 => x"80",
          5710 => x"f6",
          5711 => x"e0",
          5712 => x"ff",
          5713 => x"54",
          5714 => x"83",
          5715 => x"88",
          5716 => x"05",
          5717 => x"ff",
          5718 => x"82",
          5719 => x"14",
          5720 => x"62",
          5721 => x"5c",
          5722 => x"ff",
          5723 => x"39",
          5724 => x"54",
          5725 => x"82",
          5726 => x"5c",
          5727 => x"08",
          5728 => x"38",
          5729 => x"52",
          5730 => x"08",
          5731 => x"8a",
          5732 => x"f7",
          5733 => x"58",
          5734 => x"99",
          5735 => x"7a",
          5736 => x"f2",
          5737 => x"19",
          5738 => x"e0",
          5739 => x"84",
          5740 => x"f9",
          5741 => x"73",
          5742 => x"0c",
          5743 => x"04",
          5744 => x"77",
          5745 => x"52",
          5746 => x"3f",
          5747 => x"08",
          5748 => x"98",
          5749 => x"8e",
          5750 => x"80",
          5751 => x"98",
          5752 => x"90",
          5753 => x"82",
          5754 => x"86",
          5755 => x"ff",
          5756 => x"8f",
          5757 => x"81",
          5758 => x"26",
          5759 => x"e0",
          5760 => x"52",
          5761 => x"98",
          5762 => x"0d",
          5763 => x"0d",
          5764 => x"33",
          5765 => x"9f",
          5766 => x"53",
          5767 => x"81",
          5768 => x"38",
          5769 => x"87",
          5770 => x"11",
          5771 => x"54",
          5772 => x"84",
          5773 => x"54",
          5774 => x"87",
          5775 => x"11",
          5776 => x"0c",
          5777 => x"c0",
          5778 => x"70",
          5779 => x"70",
          5780 => x"51",
          5781 => x"8a",
          5782 => x"98",
          5783 => x"70",
          5784 => x"08",
          5785 => x"06",
          5786 => x"38",
          5787 => x"8c",
          5788 => x"80",
          5789 => x"71",
          5790 => x"14",
          5791 => x"94",
          5792 => x"70",
          5793 => x"0c",
          5794 => x"04",
          5795 => x"60",
          5796 => x"8c",
          5797 => x"33",
          5798 => x"5b",
          5799 => x"5a",
          5800 => x"82",
          5801 => x"81",
          5802 => x"52",
          5803 => x"38",
          5804 => x"84",
          5805 => x"92",
          5806 => x"c0",
          5807 => x"87",
          5808 => x"13",
          5809 => x"57",
          5810 => x"0b",
          5811 => x"8c",
          5812 => x"0c",
          5813 => x"75",
          5814 => x"2a",
          5815 => x"51",
          5816 => x"80",
          5817 => x"7b",
          5818 => x"7b",
          5819 => x"5d",
          5820 => x"59",
          5821 => x"06",
          5822 => x"73",
          5823 => x"81",
          5824 => x"ff",
          5825 => x"72",
          5826 => x"38",
          5827 => x"8c",
          5828 => x"c3",
          5829 => x"98",
          5830 => x"71",
          5831 => x"38",
          5832 => x"2e",
          5833 => x"76",
          5834 => x"92",
          5835 => x"72",
          5836 => x"06",
          5837 => x"f7",
          5838 => x"5a",
          5839 => x"80",
          5840 => x"70",
          5841 => x"5a",
          5842 => x"80",
          5843 => x"73",
          5844 => x"06",
          5845 => x"38",
          5846 => x"fe",
          5847 => x"fc",
          5848 => x"52",
          5849 => x"83",
          5850 => x"71",
          5851 => x"e0",
          5852 => x"3d",
          5853 => x"3d",
          5854 => x"64",
          5855 => x"bf",
          5856 => x"40",
          5857 => x"59",
          5858 => x"58",
          5859 => x"82",
          5860 => x"81",
          5861 => x"52",
          5862 => x"09",
          5863 => x"b1",
          5864 => x"84",
          5865 => x"92",
          5866 => x"c0",
          5867 => x"87",
          5868 => x"13",
          5869 => x"56",
          5870 => x"87",
          5871 => x"0c",
          5872 => x"82",
          5873 => x"58",
          5874 => x"84",
          5875 => x"06",
          5876 => x"71",
          5877 => x"38",
          5878 => x"05",
          5879 => x"0c",
          5880 => x"73",
          5881 => x"81",
          5882 => x"71",
          5883 => x"38",
          5884 => x"8c",
          5885 => x"d0",
          5886 => x"98",
          5887 => x"71",
          5888 => x"38",
          5889 => x"2e",
          5890 => x"76",
          5891 => x"92",
          5892 => x"72",
          5893 => x"06",
          5894 => x"f7",
          5895 => x"59",
          5896 => x"1a",
          5897 => x"06",
          5898 => x"59",
          5899 => x"80",
          5900 => x"73",
          5901 => x"06",
          5902 => x"38",
          5903 => x"fe",
          5904 => x"fc",
          5905 => x"52",
          5906 => x"83",
          5907 => x"71",
          5908 => x"e0",
          5909 => x"3d",
          5910 => x"3d",
          5911 => x"84",
          5912 => x"33",
          5913 => x"a7",
          5914 => x"54",
          5915 => x"fa",
          5916 => x"e0",
          5917 => x"06",
          5918 => x"72",
          5919 => x"85",
          5920 => x"98",
          5921 => x"56",
          5922 => x"80",
          5923 => x"76",
          5924 => x"74",
          5925 => x"c0",
          5926 => x"54",
          5927 => x"2e",
          5928 => x"d4",
          5929 => x"2e",
          5930 => x"80",
          5931 => x"08",
          5932 => x"70",
          5933 => x"51",
          5934 => x"2e",
          5935 => x"c0",
          5936 => x"52",
          5937 => x"87",
          5938 => x"08",
          5939 => x"38",
          5940 => x"87",
          5941 => x"14",
          5942 => x"70",
          5943 => x"52",
          5944 => x"96",
          5945 => x"92",
          5946 => x"0a",
          5947 => x"39",
          5948 => x"0c",
          5949 => x"39",
          5950 => x"54",
          5951 => x"98",
          5952 => x"0d",
          5953 => x"0d",
          5954 => x"33",
          5955 => x"88",
          5956 => x"e0",
          5957 => x"51",
          5958 => x"04",
          5959 => x"75",
          5960 => x"82",
          5961 => x"90",
          5962 => x"2b",
          5963 => x"33",
          5964 => x"88",
          5965 => x"71",
          5966 => x"98",
          5967 => x"54",
          5968 => x"85",
          5969 => x"ff",
          5970 => x"02",
          5971 => x"05",
          5972 => x"70",
          5973 => x"05",
          5974 => x"88",
          5975 => x"72",
          5976 => x"0d",
          5977 => x"0d",
          5978 => x"52",
          5979 => x"81",
          5980 => x"70",
          5981 => x"70",
          5982 => x"05",
          5983 => x"88",
          5984 => x"72",
          5985 => x"54",
          5986 => x"2a",
          5987 => x"34",
          5988 => x"04",
          5989 => x"76",
          5990 => x"54",
          5991 => x"2e",
          5992 => x"70",
          5993 => x"33",
          5994 => x"05",
          5995 => x"11",
          5996 => x"84",
          5997 => x"fe",
          5998 => x"77",
          5999 => x"53",
          6000 => x"81",
          6001 => x"ff",
          6002 => x"f4",
          6003 => x"0d",
          6004 => x"0d",
          6005 => x"56",
          6006 => x"70",
          6007 => x"33",
          6008 => x"05",
          6009 => x"71",
          6010 => x"56",
          6011 => x"72",
          6012 => x"38",
          6013 => x"e2",
          6014 => x"e0",
          6015 => x"3d",
          6016 => x"3d",
          6017 => x"54",
          6018 => x"71",
          6019 => x"38",
          6020 => x"70",
          6021 => x"f3",
          6022 => x"82",
          6023 => x"84",
          6024 => x"80",
          6025 => x"98",
          6026 => x"3d",
          6027 => x"08",
          6028 => x"05",
          6029 => x"54",
          6030 => x"e7",
          6031 => x"82",
          6032 => x"a2",
          6033 => x"2e",
          6034 => x"b5",
          6035 => x"80",
          6036 => x"82",
          6037 => x"83",
          6038 => x"53",
          6039 => x"86",
          6040 => x"0c",
          6041 => x"82",
          6042 => x"87",
          6043 => x"f7",
          6044 => x"56",
          6045 => x"17",
          6046 => x"74",
          6047 => x"d6",
          6048 => x"b4",
          6049 => x"b8",
          6050 => x"81",
          6051 => x"59",
          6052 => x"82",
          6053 => x"7a",
          6054 => x"06",
          6055 => x"e0",
          6056 => x"17",
          6057 => x"08",
          6058 => x"08",
          6059 => x"08",
          6060 => x"74",
          6061 => x"38",
          6062 => x"55",
          6063 => x"09",
          6064 => x"38",
          6065 => x"18",
          6066 => x"81",
          6067 => x"f9",
          6068 => x"39",
          6069 => x"82",
          6070 => x"8b",
          6071 => x"fa",
          6072 => x"7a",
          6073 => x"57",
          6074 => x"08",
          6075 => x"75",
          6076 => x"3f",
          6077 => x"08",
          6078 => x"98",
          6079 => x"81",
          6080 => x"b8",
          6081 => x"16",
          6082 => x"80",
          6083 => x"98",
          6084 => x"85",
          6085 => x"81",
          6086 => x"17",
          6087 => x"e0",
          6088 => x"3d",
          6089 => x"3d",
          6090 => x"52",
          6091 => x"3f",
          6092 => x"08",
          6093 => x"98",
          6094 => x"38",
          6095 => x"74",
          6096 => x"81",
          6097 => x"38",
          6098 => x"59",
          6099 => x"09",
          6100 => x"e3",
          6101 => x"53",
          6102 => x"08",
          6103 => x"70",
          6104 => x"d3",
          6105 => x"d5",
          6106 => x"17",
          6107 => x"3f",
          6108 => x"a4",
          6109 => x"51",
          6110 => x"86",
          6111 => x"f2",
          6112 => x"17",
          6113 => x"3f",
          6114 => x"52",
          6115 => x"51",
          6116 => x"90",
          6117 => x"84",
          6118 => x"fb",
          6119 => x"17",
          6120 => x"70",
          6121 => x"79",
          6122 => x"52",
          6123 => x"51",
          6124 => x"77",
          6125 => x"80",
          6126 => x"81",
          6127 => x"f9",
          6128 => x"e0",
          6129 => x"2e",
          6130 => x"58",
          6131 => x"98",
          6132 => x"0d",
          6133 => x"0d",
          6134 => x"9c",
          6135 => x"05",
          6136 => x"80",
          6137 => x"27",
          6138 => x"14",
          6139 => x"29",
          6140 => x"05",
          6141 => x"82",
          6142 => x"87",
          6143 => x"f9",
          6144 => x"7a",
          6145 => x"54",
          6146 => x"27",
          6147 => x"76",
          6148 => x"27",
          6149 => x"ff",
          6150 => x"58",
          6151 => x"80",
          6152 => x"82",
          6153 => x"72",
          6154 => x"38",
          6155 => x"72",
          6156 => x"8e",
          6157 => x"39",
          6158 => x"17",
          6159 => x"a8",
          6160 => x"53",
          6161 => x"fd",
          6162 => x"e0",
          6163 => x"9f",
          6164 => x"ff",
          6165 => x"11",
          6166 => x"70",
          6167 => x"18",
          6168 => x"76",
          6169 => x"53",
          6170 => x"82",
          6171 => x"80",
          6172 => x"83",
          6173 => x"b8",
          6174 => x"88",
          6175 => x"79",
          6176 => x"84",
          6177 => x"58",
          6178 => x"80",
          6179 => x"9f",
          6180 => x"80",
          6181 => x"88",
          6182 => x"08",
          6183 => x"51",
          6184 => x"82",
          6185 => x"80",
          6186 => x"10",
          6187 => x"74",
          6188 => x"51",
          6189 => x"82",
          6190 => x"83",
          6191 => x"58",
          6192 => x"87",
          6193 => x"08",
          6194 => x"51",
          6195 => x"82",
          6196 => x"9b",
          6197 => x"2b",
          6198 => x"74",
          6199 => x"51",
          6200 => x"82",
          6201 => x"f0",
          6202 => x"83",
          6203 => x"77",
          6204 => x"0c",
          6205 => x"04",
          6206 => x"7a",
          6207 => x"58",
          6208 => x"81",
          6209 => x"9e",
          6210 => x"17",
          6211 => x"96",
          6212 => x"53",
          6213 => x"81",
          6214 => x"79",
          6215 => x"72",
          6216 => x"38",
          6217 => x"72",
          6218 => x"b8",
          6219 => x"39",
          6220 => x"17",
          6221 => x"a8",
          6222 => x"53",
          6223 => x"fb",
          6224 => x"e0",
          6225 => x"82",
          6226 => x"81",
          6227 => x"83",
          6228 => x"b8",
          6229 => x"78",
          6230 => x"56",
          6231 => x"76",
          6232 => x"38",
          6233 => x"9f",
          6234 => x"33",
          6235 => x"07",
          6236 => x"74",
          6237 => x"83",
          6238 => x"89",
          6239 => x"08",
          6240 => x"51",
          6241 => x"82",
          6242 => x"59",
          6243 => x"08",
          6244 => x"74",
          6245 => x"16",
          6246 => x"84",
          6247 => x"76",
          6248 => x"88",
          6249 => x"81",
          6250 => x"8f",
          6251 => x"53",
          6252 => x"80",
          6253 => x"88",
          6254 => x"08",
          6255 => x"51",
          6256 => x"82",
          6257 => x"59",
          6258 => x"08",
          6259 => x"77",
          6260 => x"06",
          6261 => x"83",
          6262 => x"05",
          6263 => x"f6",
          6264 => x"39",
          6265 => x"a8",
          6266 => x"52",
          6267 => x"ef",
          6268 => x"98",
          6269 => x"e0",
          6270 => x"38",
          6271 => x"06",
          6272 => x"83",
          6273 => x"18",
          6274 => x"54",
          6275 => x"f6",
          6276 => x"e0",
          6277 => x"0a",
          6278 => x"52",
          6279 => x"c5",
          6280 => x"83",
          6281 => x"82",
          6282 => x"8a",
          6283 => x"f8",
          6284 => x"7c",
          6285 => x"59",
          6286 => x"81",
          6287 => x"38",
          6288 => x"08",
          6289 => x"73",
          6290 => x"38",
          6291 => x"52",
          6292 => x"a4",
          6293 => x"98",
          6294 => x"e0",
          6295 => x"f2",
          6296 => x"82",
          6297 => x"39",
          6298 => x"e6",
          6299 => x"98",
          6300 => x"de",
          6301 => x"78",
          6302 => x"3f",
          6303 => x"08",
          6304 => x"98",
          6305 => x"80",
          6306 => x"e0",
          6307 => x"2e",
          6308 => x"e0",
          6309 => x"2e",
          6310 => x"53",
          6311 => x"51",
          6312 => x"82",
          6313 => x"c5",
          6314 => x"08",
          6315 => x"18",
          6316 => x"57",
          6317 => x"90",
          6318 => x"94",
          6319 => x"16",
          6320 => x"54",
          6321 => x"34",
          6322 => x"78",
          6323 => x"38",
          6324 => x"82",
          6325 => x"8a",
          6326 => x"f6",
          6327 => x"7e",
          6328 => x"5b",
          6329 => x"38",
          6330 => x"58",
          6331 => x"88",
          6332 => x"08",
          6333 => x"38",
          6334 => x"39",
          6335 => x"51",
          6336 => x"81",
          6337 => x"e0",
          6338 => x"82",
          6339 => x"e0",
          6340 => x"82",
          6341 => x"ff",
          6342 => x"38",
          6343 => x"82",
          6344 => x"26",
          6345 => x"79",
          6346 => x"08",
          6347 => x"73",
          6348 => x"b9",
          6349 => x"2e",
          6350 => x"80",
          6351 => x"1a",
          6352 => x"08",
          6353 => x"38",
          6354 => x"52",
          6355 => x"af",
          6356 => x"82",
          6357 => x"81",
          6358 => x"06",
          6359 => x"e0",
          6360 => x"82",
          6361 => x"09",
          6362 => x"72",
          6363 => x"70",
          6364 => x"e0",
          6365 => x"51",
          6366 => x"73",
          6367 => x"82",
          6368 => x"80",
          6369 => x"90",
          6370 => x"81",
          6371 => x"38",
          6372 => x"08",
          6373 => x"73",
          6374 => x"75",
          6375 => x"77",
          6376 => x"56",
          6377 => x"76",
          6378 => x"82",
          6379 => x"26",
          6380 => x"75",
          6381 => x"f8",
          6382 => x"e0",
          6383 => x"2e",
          6384 => x"59",
          6385 => x"08",
          6386 => x"81",
          6387 => x"82",
          6388 => x"59",
          6389 => x"08",
          6390 => x"70",
          6391 => x"25",
          6392 => x"51",
          6393 => x"73",
          6394 => x"75",
          6395 => x"81",
          6396 => x"38",
          6397 => x"f5",
          6398 => x"75",
          6399 => x"f9",
          6400 => x"e0",
          6401 => x"e0",
          6402 => x"70",
          6403 => x"08",
          6404 => x"51",
          6405 => x"80",
          6406 => x"73",
          6407 => x"38",
          6408 => x"52",
          6409 => x"d0",
          6410 => x"98",
          6411 => x"a5",
          6412 => x"18",
          6413 => x"08",
          6414 => x"18",
          6415 => x"74",
          6416 => x"38",
          6417 => x"18",
          6418 => x"33",
          6419 => x"73",
          6420 => x"97",
          6421 => x"74",
          6422 => x"38",
          6423 => x"55",
          6424 => x"e0",
          6425 => x"85",
          6426 => x"75",
          6427 => x"e0",
          6428 => x"3d",
          6429 => x"3d",
          6430 => x"52",
          6431 => x"3f",
          6432 => x"08",
          6433 => x"82",
          6434 => x"80",
          6435 => x"52",
          6436 => x"c1",
          6437 => x"98",
          6438 => x"98",
          6439 => x"0c",
          6440 => x"53",
          6441 => x"15",
          6442 => x"f2",
          6443 => x"56",
          6444 => x"16",
          6445 => x"22",
          6446 => x"27",
          6447 => x"54",
          6448 => x"76",
          6449 => x"33",
          6450 => x"3f",
          6451 => x"08",
          6452 => x"38",
          6453 => x"76",
          6454 => x"70",
          6455 => x"9f",
          6456 => x"56",
          6457 => x"e0",
          6458 => x"3d",
          6459 => x"3d",
          6460 => x"71",
          6461 => x"57",
          6462 => x"0a",
          6463 => x"38",
          6464 => x"53",
          6465 => x"38",
          6466 => x"0c",
          6467 => x"54",
          6468 => x"75",
          6469 => x"73",
          6470 => x"ac",
          6471 => x"73",
          6472 => x"85",
          6473 => x"0b",
          6474 => x"5a",
          6475 => x"27",
          6476 => x"ac",
          6477 => x"18",
          6478 => x"39",
          6479 => x"70",
          6480 => x"58",
          6481 => x"b2",
          6482 => x"76",
          6483 => x"3f",
          6484 => x"08",
          6485 => x"98",
          6486 => x"bd",
          6487 => x"82",
          6488 => x"27",
          6489 => x"16",
          6490 => x"98",
          6491 => x"38",
          6492 => x"39",
          6493 => x"55",
          6494 => x"52",
          6495 => x"d5",
          6496 => x"98",
          6497 => x"0c",
          6498 => x"0c",
          6499 => x"53",
          6500 => x"80",
          6501 => x"85",
          6502 => x"94",
          6503 => x"2a",
          6504 => x"0c",
          6505 => x"06",
          6506 => x"9c",
          6507 => x"58",
          6508 => x"98",
          6509 => x"0d",
          6510 => x"0d",
          6511 => x"90",
          6512 => x"05",
          6513 => x"f0",
          6514 => x"27",
          6515 => x"0b",
          6516 => x"98",
          6517 => x"84",
          6518 => x"2e",
          6519 => x"76",
          6520 => x"58",
          6521 => x"38",
          6522 => x"15",
          6523 => x"08",
          6524 => x"38",
          6525 => x"88",
          6526 => x"53",
          6527 => x"81",
          6528 => x"c0",
          6529 => x"22",
          6530 => x"89",
          6531 => x"72",
          6532 => x"74",
          6533 => x"f3",
          6534 => x"e0",
          6535 => x"82",
          6536 => x"82",
          6537 => x"27",
          6538 => x"81",
          6539 => x"98",
          6540 => x"80",
          6541 => x"16",
          6542 => x"98",
          6543 => x"ca",
          6544 => x"38",
          6545 => x"0c",
          6546 => x"dd",
          6547 => x"08",
          6548 => x"f9",
          6549 => x"e0",
          6550 => x"87",
          6551 => x"98",
          6552 => x"80",
          6553 => x"55",
          6554 => x"08",
          6555 => x"38",
          6556 => x"e0",
          6557 => x"2e",
          6558 => x"e0",
          6559 => x"75",
          6560 => x"3f",
          6561 => x"08",
          6562 => x"94",
          6563 => x"52",
          6564 => x"c1",
          6565 => x"98",
          6566 => x"0c",
          6567 => x"0c",
          6568 => x"05",
          6569 => x"80",
          6570 => x"e0",
          6571 => x"3d",
          6572 => x"3d",
          6573 => x"71",
          6574 => x"57",
          6575 => x"51",
          6576 => x"82",
          6577 => x"54",
          6578 => x"08",
          6579 => x"82",
          6580 => x"56",
          6581 => x"52",
          6582 => x"83",
          6583 => x"98",
          6584 => x"e0",
          6585 => x"d2",
          6586 => x"98",
          6587 => x"08",
          6588 => x"54",
          6589 => x"e5",
          6590 => x"06",
          6591 => x"58",
          6592 => x"08",
          6593 => x"38",
          6594 => x"75",
          6595 => x"80",
          6596 => x"81",
          6597 => x"7a",
          6598 => x"06",
          6599 => x"39",
          6600 => x"08",
          6601 => x"76",
          6602 => x"3f",
          6603 => x"08",
          6604 => x"98",
          6605 => x"ff",
          6606 => x"84",
          6607 => x"06",
          6608 => x"54",
          6609 => x"98",
          6610 => x"0d",
          6611 => x"0d",
          6612 => x"52",
          6613 => x"3f",
          6614 => x"08",
          6615 => x"06",
          6616 => x"51",
          6617 => x"83",
          6618 => x"06",
          6619 => x"14",
          6620 => x"3f",
          6621 => x"08",
          6622 => x"07",
          6623 => x"e0",
          6624 => x"3d",
          6625 => x"3d",
          6626 => x"70",
          6627 => x"06",
          6628 => x"53",
          6629 => x"af",
          6630 => x"33",
          6631 => x"83",
          6632 => x"06",
          6633 => x"90",
          6634 => x"15",
          6635 => x"3f",
          6636 => x"04",
          6637 => x"75",
          6638 => x"8b",
          6639 => x"2a",
          6640 => x"29",
          6641 => x"81",
          6642 => x"71",
          6643 => x"ff",
          6644 => x"56",
          6645 => x"72",
          6646 => x"82",
          6647 => x"85",
          6648 => x"f2",
          6649 => x"62",
          6650 => x"79",
          6651 => x"81",
          6652 => x"5d",
          6653 => x"80",
          6654 => x"38",
          6655 => x"52",
          6656 => x"db",
          6657 => x"98",
          6658 => x"e0",
          6659 => x"eb",
          6660 => x"08",
          6661 => x"55",
          6662 => x"84",
          6663 => x"39",
          6664 => x"bf",
          6665 => x"ff",
          6666 => x"72",
          6667 => x"82",
          6668 => x"56",
          6669 => x"2e",
          6670 => x"83",
          6671 => x"82",
          6672 => x"53",
          6673 => x"09",
          6674 => x"38",
          6675 => x"73",
          6676 => x"99",
          6677 => x"98",
          6678 => x"06",
          6679 => x"88",
          6680 => x"06",
          6681 => x"56",
          6682 => x"87",
          6683 => x"5c",
          6684 => x"76",
          6685 => x"81",
          6686 => x"38",
          6687 => x"70",
          6688 => x"53",
          6689 => x"92",
          6690 => x"33",
          6691 => x"06",
          6692 => x"08",
          6693 => x"56",
          6694 => x"7c",
          6695 => x"06",
          6696 => x"8d",
          6697 => x"7c",
          6698 => x"81",
          6699 => x"38",
          6700 => x"9a",
          6701 => x"e8",
          6702 => x"e0",
          6703 => x"ff",
          6704 => x"72",
          6705 => x"74",
          6706 => x"bf",
          6707 => x"f3",
          6708 => x"81",
          6709 => x"82",
          6710 => x"33",
          6711 => x"e8",
          6712 => x"e0",
          6713 => x"ff",
          6714 => x"77",
          6715 => x"38",
          6716 => x"26",
          6717 => x"73",
          6718 => x"59",
          6719 => x"23",
          6720 => x"8b",
          6721 => x"ff",
          6722 => x"81",
          6723 => x"81",
          6724 => x"77",
          6725 => x"74",
          6726 => x"2a",
          6727 => x"51",
          6728 => x"80",
          6729 => x"73",
          6730 => x"92",
          6731 => x"1a",
          6732 => x"23",
          6733 => x"81",
          6734 => x"53",
          6735 => x"ff",
          6736 => x"9d",
          6737 => x"38",
          6738 => x"e8",
          6739 => x"98",
          6740 => x"06",
          6741 => x"2e",
          6742 => x"0b",
          6743 => x"a0",
          6744 => x"78",
          6745 => x"3f",
          6746 => x"08",
          6747 => x"98",
          6748 => x"98",
          6749 => x"84",
          6750 => x"80",
          6751 => x"0c",
          6752 => x"98",
          6753 => x"0d",
          6754 => x"0d",
          6755 => x"40",
          6756 => x"78",
          6757 => x"3f",
          6758 => x"08",
          6759 => x"98",
          6760 => x"38",
          6761 => x"5f",
          6762 => x"ac",
          6763 => x"19",
          6764 => x"51",
          6765 => x"82",
          6766 => x"58",
          6767 => x"08",
          6768 => x"9c",
          6769 => x"33",
          6770 => x"86",
          6771 => x"82",
          6772 => x"17",
          6773 => x"70",
          6774 => x"56",
          6775 => x"1a",
          6776 => x"e5",
          6777 => x"38",
          6778 => x"70",
          6779 => x"54",
          6780 => x"8e",
          6781 => x"b2",
          6782 => x"2e",
          6783 => x"81",
          6784 => x"19",
          6785 => x"2a",
          6786 => x"51",
          6787 => x"82",
          6788 => x"86",
          6789 => x"06",
          6790 => x"80",
          6791 => x"8d",
          6792 => x"81",
          6793 => x"90",
          6794 => x"1d",
          6795 => x"5e",
          6796 => x"09",
          6797 => x"b9",
          6798 => x"33",
          6799 => x"2e",
          6800 => x"81",
          6801 => x"1f",
          6802 => x"52",
          6803 => x"3f",
          6804 => x"08",
          6805 => x"06",
          6806 => x"95",
          6807 => x"70",
          6808 => x"29",
          6809 => x"56",
          6810 => x"5a",
          6811 => x"1b",
          6812 => x"51",
          6813 => x"82",
          6814 => x"83",
          6815 => x"56",
          6816 => x"b1",
          6817 => x"fe",
          6818 => x"38",
          6819 => x"e1",
          6820 => x"e0",
          6821 => x"10",
          6822 => x"53",
          6823 => x"59",
          6824 => x"8d",
          6825 => x"e0",
          6826 => x"09",
          6827 => x"c1",
          6828 => x"8b",
          6829 => x"ff",
          6830 => x"81",
          6831 => x"81",
          6832 => x"7b",
          6833 => x"38",
          6834 => x"86",
          6835 => x"06",
          6836 => x"79",
          6837 => x"38",
          6838 => x"8b",
          6839 => x"1d",
          6840 => x"54",
          6841 => x"ff",
          6842 => x"ff",
          6843 => x"84",
          6844 => x"54",
          6845 => x"39",
          6846 => x"76",
          6847 => x"3f",
          6848 => x"08",
          6849 => x"54",
          6850 => x"bb",
          6851 => x"33",
          6852 => x"73",
          6853 => x"53",
          6854 => x"9c",
          6855 => x"e5",
          6856 => x"e0",
          6857 => x"2e",
          6858 => x"ff",
          6859 => x"ac",
          6860 => x"52",
          6861 => x"81",
          6862 => x"98",
          6863 => x"e0",
          6864 => x"2e",
          6865 => x"77",
          6866 => x"0c",
          6867 => x"04",
          6868 => x"64",
          6869 => x"12",
          6870 => x"06",
          6871 => x"86",
          6872 => x"b5",
          6873 => x"1d",
          6874 => x"56",
          6875 => x"80",
          6876 => x"81",
          6877 => x"16",
          6878 => x"55",
          6879 => x"8c",
          6880 => x"70",
          6881 => x"70",
          6882 => x"e4",
          6883 => x"80",
          6884 => x"81",
          6885 => x"80",
          6886 => x"38",
          6887 => x"ab",
          6888 => x"5b",
          6889 => x"7b",
          6890 => x"53",
          6891 => x"51",
          6892 => x"85",
          6893 => x"c6",
          6894 => x"77",
          6895 => x"ff",
          6896 => x"55",
          6897 => x"b4",
          6898 => x"ff",
          6899 => x"19",
          6900 => x"57",
          6901 => x"76",
          6902 => x"81",
          6903 => x"2a",
          6904 => x"51",
          6905 => x"73",
          6906 => x"38",
          6907 => x"a1",
          6908 => x"17",
          6909 => x"25",
          6910 => x"39",
          6911 => x"02",
          6912 => x"05",
          6913 => x"b0",
          6914 => x"54",
          6915 => x"84",
          6916 => x"54",
          6917 => x"ff",
          6918 => x"76",
          6919 => x"58",
          6920 => x"38",
          6921 => x"05",
          6922 => x"fe",
          6923 => x"77",
          6924 => x"78",
          6925 => x"a0",
          6926 => x"74",
          6927 => x"52",
          6928 => x"3f",
          6929 => x"08",
          6930 => x"38",
          6931 => x"74",
          6932 => x"38",
          6933 => x"81",
          6934 => x"77",
          6935 => x"74",
          6936 => x"51",
          6937 => x"94",
          6938 => x"eb",
          6939 => x"15",
          6940 => x"58",
          6941 => x"87",
          6942 => x"81",
          6943 => x"70",
          6944 => x"57",
          6945 => x"87",
          6946 => x"38",
          6947 => x"f9",
          6948 => x"98",
          6949 => x"81",
          6950 => x"e3",
          6951 => x"84",
          6952 => x"7a",
          6953 => x"82",
          6954 => x"e0",
          6955 => x"82",
          6956 => x"84",
          6957 => x"06",
          6958 => x"02",
          6959 => x"33",
          6960 => x"02",
          6961 => x"33",
          6962 => x"70",
          6963 => x"55",
          6964 => x"73",
          6965 => x"38",
          6966 => x"1d",
          6967 => x"f4",
          6968 => x"98",
          6969 => x"78",
          6970 => x"f3",
          6971 => x"e0",
          6972 => x"82",
          6973 => x"82",
          6974 => x"19",
          6975 => x"2e",
          6976 => x"78",
          6977 => x"1b",
          6978 => x"53",
          6979 => x"ef",
          6980 => x"e0",
          6981 => x"82",
          6982 => x"81",
          6983 => x"1a",
          6984 => x"3f",
          6985 => x"08",
          6986 => x"5d",
          6987 => x"52",
          6988 => x"ab",
          6989 => x"98",
          6990 => x"e0",
          6991 => x"d7",
          6992 => x"08",
          6993 => x"7a",
          6994 => x"5a",
          6995 => x"8d",
          6996 => x"0b",
          6997 => x"82",
          6998 => x"8c",
          6999 => x"e0",
          7000 => x"9a",
          7001 => x"df",
          7002 => x"29",
          7003 => x"55",
          7004 => x"ff",
          7005 => x"38",
          7006 => x"70",
          7007 => x"57",
          7008 => x"52",
          7009 => x"17",
          7010 => x"51",
          7011 => x"73",
          7012 => x"ff",
          7013 => x"17",
          7014 => x"27",
          7015 => x"83",
          7016 => x"8b",
          7017 => x"1b",
          7018 => x"54",
          7019 => x"77",
          7020 => x"58",
          7021 => x"81",
          7022 => x"34",
          7023 => x"51",
          7024 => x"82",
          7025 => x"57",
          7026 => x"08",
          7027 => x"ff",
          7028 => x"fe",
          7029 => x"1a",
          7030 => x"51",
          7031 => x"82",
          7032 => x"57",
          7033 => x"08",
          7034 => x"53",
          7035 => x"08",
          7036 => x"08",
          7037 => x"3f",
          7038 => x"1a",
          7039 => x"08",
          7040 => x"3f",
          7041 => x"ab",
          7042 => x"06",
          7043 => x"8c",
          7044 => x"0b",
          7045 => x"76",
          7046 => x"e0",
          7047 => x"3d",
          7048 => x"3d",
          7049 => x"08",
          7050 => x"ac",
          7051 => x"59",
          7052 => x"ff",
          7053 => x"72",
          7054 => x"ed",
          7055 => x"e0",
          7056 => x"82",
          7057 => x"80",
          7058 => x"15",
          7059 => x"51",
          7060 => x"82",
          7061 => x"54",
          7062 => x"08",
          7063 => x"15",
          7064 => x"73",
          7065 => x"83",
          7066 => x"15",
          7067 => x"a2",
          7068 => x"98",
          7069 => x"51",
          7070 => x"82",
          7071 => x"54",
          7072 => x"08",
          7073 => x"38",
          7074 => x"09",
          7075 => x"38",
          7076 => x"82",
          7077 => x"88",
          7078 => x"f4",
          7079 => x"60",
          7080 => x"59",
          7081 => x"96",
          7082 => x"1c",
          7083 => x"83",
          7084 => x"1c",
          7085 => x"81",
          7086 => x"70",
          7087 => x"05",
          7088 => x"57",
          7089 => x"57",
          7090 => x"81",
          7091 => x"10",
          7092 => x"81",
          7093 => x"53",
          7094 => x"80",
          7095 => x"70",
          7096 => x"06",
          7097 => x"8f",
          7098 => x"38",
          7099 => x"df",
          7100 => x"96",
          7101 => x"79",
          7102 => x"54",
          7103 => x"7a",
          7104 => x"07",
          7105 => x"84",
          7106 => x"98",
          7107 => x"ff",
          7108 => x"ff",
          7109 => x"38",
          7110 => x"a5",
          7111 => x"2a",
          7112 => x"34",
          7113 => x"34",
          7114 => x"39",
          7115 => x"30",
          7116 => x"80",
          7117 => x"25",
          7118 => x"54",
          7119 => x"85",
          7120 => x"9a",
          7121 => x"34",
          7122 => x"17",
          7123 => x"8c",
          7124 => x"10",
          7125 => x"51",
          7126 => x"fe",
          7127 => x"30",
          7128 => x"70",
          7129 => x"59",
          7130 => x"17",
          7131 => x"80",
          7132 => x"34",
          7133 => x"1a",
          7134 => x"9c",
          7135 => x"70",
          7136 => x"5b",
          7137 => x"a0",
          7138 => x"74",
          7139 => x"81",
          7140 => x"81",
          7141 => x"89",
          7142 => x"70",
          7143 => x"25",
          7144 => x"76",
          7145 => x"38",
          7146 => x"8b",
          7147 => x"70",
          7148 => x"34",
          7149 => x"74",
          7150 => x"05",
          7151 => x"17",
          7152 => x"27",
          7153 => x"77",
          7154 => x"53",
          7155 => x"14",
          7156 => x"33",
          7157 => x"87",
          7158 => x"38",
          7159 => x"19",
          7160 => x"80",
          7161 => x"73",
          7162 => x"55",
          7163 => x"80",
          7164 => x"38",
          7165 => x"19",
          7166 => x"33",
          7167 => x"54",
          7168 => x"26",
          7169 => x"1c",
          7170 => x"33",
          7171 => x"79",
          7172 => x"72",
          7173 => x"85",
          7174 => x"2a",
          7175 => x"06",
          7176 => x"2e",
          7177 => x"15",
          7178 => x"ff",
          7179 => x"74",
          7180 => x"05",
          7181 => x"19",
          7182 => x"19",
          7183 => x"59",
          7184 => x"ff",
          7185 => x"17",
          7186 => x"80",
          7187 => x"34",
          7188 => x"8c",
          7189 => x"53",
          7190 => x"72",
          7191 => x"9c",
          7192 => x"8b",
          7193 => x"19",
          7194 => x"08",
          7195 => x"53",
          7196 => x"82",
          7197 => x"78",
          7198 => x"51",
          7199 => x"82",
          7200 => x"86",
          7201 => x"13",
          7202 => x"3f",
          7203 => x"08",
          7204 => x"8e",
          7205 => x"f0",
          7206 => x"70",
          7207 => x"80",
          7208 => x"51",
          7209 => x"af",
          7210 => x"81",
          7211 => x"dc",
          7212 => x"74",
          7213 => x"38",
          7214 => x"08",
          7215 => x"aa",
          7216 => x"44",
          7217 => x"33",
          7218 => x"73",
          7219 => x"81",
          7220 => x"81",
          7221 => x"dc",
          7222 => x"70",
          7223 => x"07",
          7224 => x"73",
          7225 => x"88",
          7226 => x"70",
          7227 => x"73",
          7228 => x"38",
          7229 => x"ab",
          7230 => x"52",
          7231 => x"ee",
          7232 => x"98",
          7233 => x"e1",
          7234 => x"7d",
          7235 => x"08",
          7236 => x"59",
          7237 => x"05",
          7238 => x"3f",
          7239 => x"08",
          7240 => x"b1",
          7241 => x"ff",
          7242 => x"98",
          7243 => x"38",
          7244 => x"82",
          7245 => x"90",
          7246 => x"73",
          7247 => x"19",
          7248 => x"98",
          7249 => x"ff",
          7250 => x"32",
          7251 => x"73",
          7252 => x"25",
          7253 => x"55",
          7254 => x"38",
          7255 => x"2e",
          7256 => x"80",
          7257 => x"38",
          7258 => x"d1",
          7259 => x"92",
          7260 => x"98",
          7261 => x"38",
          7262 => x"26",
          7263 => x"78",
          7264 => x"75",
          7265 => x"19",
          7266 => x"39",
          7267 => x"80",
          7268 => x"56",
          7269 => x"af",
          7270 => x"06",
          7271 => x"57",
          7272 => x"32",
          7273 => x"80",
          7274 => x"51",
          7275 => x"dc",
          7276 => x"9f",
          7277 => x"2b",
          7278 => x"2e",
          7279 => x"8c",
          7280 => x"54",
          7281 => x"a5",
          7282 => x"39",
          7283 => x"09",
          7284 => x"c9",
          7285 => x"22",
          7286 => x"2e",
          7287 => x"80",
          7288 => x"22",
          7289 => x"2e",
          7290 => x"b6",
          7291 => x"1a",
          7292 => x"23",
          7293 => x"1f",
          7294 => x"54",
          7295 => x"83",
          7296 => x"73",
          7297 => x"05",
          7298 => x"18",
          7299 => x"27",
          7300 => x"a0",
          7301 => x"ab",
          7302 => x"c4",
          7303 => x"2e",
          7304 => x"10",
          7305 => x"55",
          7306 => x"16",
          7307 => x"32",
          7308 => x"9f",
          7309 => x"53",
          7310 => x"75",
          7311 => x"38",
          7312 => x"ff",
          7313 => x"e0",
          7314 => x"7a",
          7315 => x"80",
          7316 => x"8d",
          7317 => x"85",
          7318 => x"83",
          7319 => x"99",
          7320 => x"22",
          7321 => x"ff",
          7322 => x"5d",
          7323 => x"09",
          7324 => x"38",
          7325 => x"10",
          7326 => x"51",
          7327 => x"a0",
          7328 => x"7c",
          7329 => x"83",
          7330 => x"54",
          7331 => x"09",
          7332 => x"38",
          7333 => x"57",
          7334 => x"aa",
          7335 => x"fe",
          7336 => x"51",
          7337 => x"2e",
          7338 => x"10",
          7339 => x"55",
          7340 => x"78",
          7341 => x"38",
          7342 => x"22",
          7343 => x"ae",
          7344 => x"06",
          7345 => x"53",
          7346 => x"1e",
          7347 => x"3f",
          7348 => x"5c",
          7349 => x"10",
          7350 => x"81",
          7351 => x"54",
          7352 => x"82",
          7353 => x"a0",
          7354 => x"75",
          7355 => x"30",
          7356 => x"51",
          7357 => x"79",
          7358 => x"73",
          7359 => x"38",
          7360 => x"57",
          7361 => x"54",
          7362 => x"78",
          7363 => x"81",
          7364 => x"32",
          7365 => x"72",
          7366 => x"70",
          7367 => x"51",
          7368 => x"80",
          7369 => x"7e",
          7370 => x"ae",
          7371 => x"2e",
          7372 => x"83",
          7373 => x"79",
          7374 => x"38",
          7375 => x"58",
          7376 => x"2b",
          7377 => x"5d",
          7378 => x"39",
          7379 => x"27",
          7380 => x"82",
          7381 => x"b5",
          7382 => x"80",
          7383 => x"82",
          7384 => x"83",
          7385 => x"70",
          7386 => x"81",
          7387 => x"56",
          7388 => x"8c",
          7389 => x"ff",
          7390 => x"b8",
          7391 => x"54",
          7392 => x"27",
          7393 => x"1f",
          7394 => x"26",
          7395 => x"83",
          7396 => x"57",
          7397 => x"7d",
          7398 => x"76",
          7399 => x"55",
          7400 => x"81",
          7401 => x"c3",
          7402 => x"2e",
          7403 => x"52",
          7404 => x"51",
          7405 => x"82",
          7406 => x"80",
          7407 => x"80",
          7408 => x"07",
          7409 => x"39",
          7410 => x"54",
          7411 => x"85",
          7412 => x"07",
          7413 => x"16",
          7414 => x"26",
          7415 => x"81",
          7416 => x"70",
          7417 => x"06",
          7418 => x"7d",
          7419 => x"54",
          7420 => x"81",
          7421 => x"de",
          7422 => x"33",
          7423 => x"e5",
          7424 => x"06",
          7425 => x"0b",
          7426 => x"7e",
          7427 => x"81",
          7428 => x"7b",
          7429 => x"fc",
          7430 => x"8c",
          7431 => x"8c",
          7432 => x"7b",
          7433 => x"73",
          7434 => x"81",
          7435 => x"76",
          7436 => x"76",
          7437 => x"81",
          7438 => x"73",
          7439 => x"81",
          7440 => x"80",
          7441 => x"76",
          7442 => x"7b",
          7443 => x"81",
          7444 => x"73",
          7445 => x"38",
          7446 => x"57",
          7447 => x"34",
          7448 => x"a5",
          7449 => x"98",
          7450 => x"33",
          7451 => x"e0",
          7452 => x"2e",
          7453 => x"e0",
          7454 => x"2e",
          7455 => x"80",
          7456 => x"85",
          7457 => x"06",
          7458 => x"57",
          7459 => x"80",
          7460 => x"74",
          7461 => x"73",
          7462 => x"ed",
          7463 => x"0b",
          7464 => x"80",
          7465 => x"39",
          7466 => x"54",
          7467 => x"85",
          7468 => x"74",
          7469 => x"81",
          7470 => x"73",
          7471 => x"1e",
          7472 => x"2a",
          7473 => x"51",
          7474 => x"80",
          7475 => x"90",
          7476 => x"ff",
          7477 => x"b8",
          7478 => x"51",
          7479 => x"82",
          7480 => x"88",
          7481 => x"a1",
          7482 => x"e0",
          7483 => x"3d",
          7484 => x"3d",
          7485 => x"ff",
          7486 => x"71",
          7487 => x"5c",
          7488 => x"80",
          7489 => x"38",
          7490 => x"05",
          7491 => x"9f",
          7492 => x"71",
          7493 => x"38",
          7494 => x"71",
          7495 => x"81",
          7496 => x"38",
          7497 => x"11",
          7498 => x"06",
          7499 => x"70",
          7500 => x"38",
          7501 => x"81",
          7502 => x"05",
          7503 => x"76",
          7504 => x"38",
          7505 => x"d2",
          7506 => x"77",
          7507 => x"57",
          7508 => x"05",
          7509 => x"70",
          7510 => x"33",
          7511 => x"53",
          7512 => x"99",
          7513 => x"e0",
          7514 => x"ff",
          7515 => x"ff",
          7516 => x"70",
          7517 => x"38",
          7518 => x"81",
          7519 => x"51",
          7520 => x"9f",
          7521 => x"72",
          7522 => x"81",
          7523 => x"70",
          7524 => x"72",
          7525 => x"32",
          7526 => x"72",
          7527 => x"73",
          7528 => x"53",
          7529 => x"70",
          7530 => x"38",
          7531 => x"19",
          7532 => x"75",
          7533 => x"38",
          7534 => x"83",
          7535 => x"74",
          7536 => x"59",
          7537 => x"39",
          7538 => x"33",
          7539 => x"e0",
          7540 => x"3d",
          7541 => x"3d",
          7542 => x"80",
          7543 => x"34",
          7544 => x"17",
          7545 => x"75",
          7546 => x"3f",
          7547 => x"e0",
          7548 => x"80",
          7549 => x"16",
          7550 => x"3f",
          7551 => x"08",
          7552 => x"06",
          7553 => x"73",
          7554 => x"2e",
          7555 => x"80",
          7556 => x"0b",
          7557 => x"56",
          7558 => x"e9",
          7559 => x"06",
          7560 => x"57",
          7561 => x"32",
          7562 => x"80",
          7563 => x"51",
          7564 => x"8a",
          7565 => x"e8",
          7566 => x"06",
          7567 => x"53",
          7568 => x"52",
          7569 => x"51",
          7570 => x"82",
          7571 => x"55",
          7572 => x"08",
          7573 => x"38",
          7574 => x"d1",
          7575 => x"8a",
          7576 => x"ed",
          7577 => x"98",
          7578 => x"e0",
          7579 => x"2e",
          7580 => x"55",
          7581 => x"98",
          7582 => x"0d",
          7583 => x"0d",
          7584 => x"05",
          7585 => x"33",
          7586 => x"75",
          7587 => x"fc",
          7588 => x"e0",
          7589 => x"8b",
          7590 => x"82",
          7591 => x"24",
          7592 => x"82",
          7593 => x"84",
          7594 => x"e0",
          7595 => x"55",
          7596 => x"73",
          7597 => x"b1",
          7598 => x"0c",
          7599 => x"06",
          7600 => x"57",
          7601 => x"ae",
          7602 => x"33",
          7603 => x"3f",
          7604 => x"08",
          7605 => x"70",
          7606 => x"55",
          7607 => x"76",
          7608 => x"83",
          7609 => x"2a",
          7610 => x"51",
          7611 => x"72",
          7612 => x"86",
          7613 => x"74",
          7614 => x"59",
          7615 => x"19",
          7616 => x"34",
          7617 => x"14",
          7618 => x"81",
          7619 => x"98",
          7620 => x"06",
          7621 => x"54",
          7622 => x"72",
          7623 => x"76",
          7624 => x"38",
          7625 => x"70",
          7626 => x"53",
          7627 => x"86",
          7628 => x"70",
          7629 => x"5b",
          7630 => x"82",
          7631 => x"81",
          7632 => x"76",
          7633 => x"38",
          7634 => x"81",
          7635 => x"e0",
          7636 => x"53",
          7637 => x"81",
          7638 => x"3d",
          7639 => x"83",
          7640 => x"15",
          7641 => x"53",
          7642 => x"8d",
          7643 => x"15",
          7644 => x"3f",
          7645 => x"08",
          7646 => x"70",
          7647 => x"0c",
          7648 => x"16",
          7649 => x"80",
          7650 => x"77",
          7651 => x"8d",
          7652 => x"30",
          7653 => x"72",
          7654 => x"3d",
          7655 => x"05",
          7656 => x"53",
          7657 => x"59",
          7658 => x"83",
          7659 => x"2e",
          7660 => x"52",
          7661 => x"9e",
          7662 => x"98",
          7663 => x"06",
          7664 => x"82",
          7665 => x"33",
          7666 => x"78",
          7667 => x"06",
          7668 => x"58",
          7669 => x"91",
          7670 => x"2e",
          7671 => x"16",
          7672 => x"56",
          7673 => x"c0",
          7674 => x"76",
          7675 => x"f9",
          7676 => x"76",
          7677 => x"f1",
          7678 => x"14",
          7679 => x"3f",
          7680 => x"08",
          7681 => x"06",
          7682 => x"80",
          7683 => x"06",
          7684 => x"80",
          7685 => x"c9",
          7686 => x"e0",
          7687 => x"ff",
          7688 => x"77",
          7689 => x"dc",
          7690 => x"f0",
          7691 => x"98",
          7692 => x"a0",
          7693 => x"c8",
          7694 => x"15",
          7695 => x"14",
          7696 => x"70",
          7697 => x"51",
          7698 => x"56",
          7699 => x"84",
          7700 => x"81",
          7701 => x"71",
          7702 => x"16",
          7703 => x"53",
          7704 => x"23",
          7705 => x"8b",
          7706 => x"73",
          7707 => x"80",
          7708 => x"8d",
          7709 => x"39",
          7710 => x"51",
          7711 => x"82",
          7712 => x"53",
          7713 => x"08",
          7714 => x"72",
          7715 => x"8d",
          7716 => x"d5",
          7717 => x"14",
          7718 => x"3f",
          7719 => x"08",
          7720 => x"06",
          7721 => x"38",
          7722 => x"51",
          7723 => x"82",
          7724 => x"55",
          7725 => x"51",
          7726 => x"82",
          7727 => x"83",
          7728 => x"53",
          7729 => x"80",
          7730 => x"38",
          7731 => x"78",
          7732 => x"2a",
          7733 => x"78",
          7734 => x"8d",
          7735 => x"22",
          7736 => x"31",
          7737 => x"ec",
          7738 => x"98",
          7739 => x"e0",
          7740 => x"2e",
          7741 => x"82",
          7742 => x"80",
          7743 => x"f5",
          7744 => x"83",
          7745 => x"ff",
          7746 => x"38",
          7747 => x"9f",
          7748 => x"38",
          7749 => x"39",
          7750 => x"80",
          7751 => x"38",
          7752 => x"9c",
          7753 => x"a4",
          7754 => x"1c",
          7755 => x"0c",
          7756 => x"17",
          7757 => x"76",
          7758 => x"81",
          7759 => x"80",
          7760 => x"c7",
          7761 => x"e0",
          7762 => x"ff",
          7763 => x"8d",
          7764 => x"95",
          7765 => x"91",
          7766 => x"14",
          7767 => x"3f",
          7768 => x"08",
          7769 => x"74",
          7770 => x"a2",
          7771 => x"79",
          7772 => x"f5",
          7773 => x"ac",
          7774 => x"15",
          7775 => x"2e",
          7776 => x"10",
          7777 => x"2a",
          7778 => x"05",
          7779 => x"ff",
          7780 => x"53",
          7781 => x"a0",
          7782 => x"81",
          7783 => x"0b",
          7784 => x"ff",
          7785 => x"0c",
          7786 => x"84",
          7787 => x"83",
          7788 => x"06",
          7789 => x"80",
          7790 => x"c6",
          7791 => x"e0",
          7792 => x"ff",
          7793 => x"72",
          7794 => x"81",
          7795 => x"38",
          7796 => x"73",
          7797 => x"3f",
          7798 => x"08",
          7799 => x"82",
          7800 => x"84",
          7801 => x"b6",
          7802 => x"99",
          7803 => x"98",
          7804 => x"ff",
          7805 => x"82",
          7806 => x"09",
          7807 => x"c8",
          7808 => x"51",
          7809 => x"82",
          7810 => x"84",
          7811 => x"d2",
          7812 => x"06",
          7813 => x"9c",
          7814 => x"80",
          7815 => x"98",
          7816 => x"85",
          7817 => x"09",
          7818 => x"38",
          7819 => x"51",
          7820 => x"82",
          7821 => x"94",
          7822 => x"a4",
          7823 => x"dc",
          7824 => x"98",
          7825 => x"0c",
          7826 => x"82",
          7827 => x"81",
          7828 => x"82",
          7829 => x"72",
          7830 => x"82",
          7831 => x"8c",
          7832 => x"0b",
          7833 => x"80",
          7834 => x"e0",
          7835 => x"3d",
          7836 => x"3d",
          7837 => x"89",
          7838 => x"2e",
          7839 => x"08",
          7840 => x"2e",
          7841 => x"33",
          7842 => x"2e",
          7843 => x"13",
          7844 => x"22",
          7845 => x"76",
          7846 => x"06",
          7847 => x"13",
          7848 => x"be",
          7849 => x"e0",
          7850 => x"06",
          7851 => x"38",
          7852 => x"54",
          7853 => x"80",
          7854 => x"71",
          7855 => x"82",
          7856 => x"87",
          7857 => x"fa",
          7858 => x"ab",
          7859 => x"58",
          7860 => x"05",
          7861 => x"9a",
          7862 => x"80",
          7863 => x"98",
          7864 => x"38",
          7865 => x"08",
          7866 => x"f7",
          7867 => x"08",
          7868 => x"80",
          7869 => x"80",
          7870 => x"54",
          7871 => x"84",
          7872 => x"34",
          7873 => x"75",
          7874 => x"2e",
          7875 => x"53",
          7876 => x"53",
          7877 => x"f6",
          7878 => x"e0",
          7879 => x"73",
          7880 => x"0c",
          7881 => x"04",
          7882 => x"68",
          7883 => x"80",
          7884 => x"59",
          7885 => x"78",
          7886 => x"c8",
          7887 => x"06",
          7888 => x"3d",
          7889 => x"9a",
          7890 => x"52",
          7891 => x"3f",
          7892 => x"08",
          7893 => x"98",
          7894 => x"38",
          7895 => x"52",
          7896 => x"52",
          7897 => x"3f",
          7898 => x"08",
          7899 => x"98",
          7900 => x"02",
          7901 => x"33",
          7902 => x"55",
          7903 => x"25",
          7904 => x"55",
          7905 => x"54",
          7906 => x"81",
          7907 => x"80",
          7908 => x"74",
          7909 => x"81",
          7910 => x"75",
          7911 => x"3f",
          7912 => x"08",
          7913 => x"02",
          7914 => x"91",
          7915 => x"81",
          7916 => x"82",
          7917 => x"06",
          7918 => x"80",
          7919 => x"88",
          7920 => x"39",
          7921 => x"58",
          7922 => x"38",
          7923 => x"70",
          7924 => x"54",
          7925 => x"81",
          7926 => x"52",
          7927 => x"ed",
          7928 => x"98",
          7929 => x"88",
          7930 => x"62",
          7931 => x"c2",
          7932 => x"54",
          7933 => x"15",
          7934 => x"62",
          7935 => x"d7",
          7936 => x"52",
          7937 => x"51",
          7938 => x"7a",
          7939 => x"83",
          7940 => x"80",
          7941 => x"38",
          7942 => x"08",
          7943 => x"53",
          7944 => x"3d",
          7945 => x"cc",
          7946 => x"e0",
          7947 => x"82",
          7948 => x"82",
          7949 => x"39",
          7950 => x"38",
          7951 => x"33",
          7952 => x"70",
          7953 => x"55",
          7954 => x"2e",
          7955 => x"55",
          7956 => x"77",
          7957 => x"81",
          7958 => x"73",
          7959 => x"38",
          7960 => x"54",
          7961 => x"a0",
          7962 => x"82",
          7963 => x"52",
          7964 => x"eb",
          7965 => x"98",
          7966 => x"18",
          7967 => x"55",
          7968 => x"98",
          7969 => x"38",
          7970 => x"70",
          7971 => x"54",
          7972 => x"86",
          7973 => x"c0",
          7974 => x"b4",
          7975 => x"1b",
          7976 => x"1b",
          7977 => x"70",
          7978 => x"a1",
          7979 => x"98",
          7980 => x"98",
          7981 => x"0c",
          7982 => x"52",
          7983 => x"3f",
          7984 => x"08",
          7985 => x"08",
          7986 => x"77",
          7987 => x"86",
          7988 => x"1a",
          7989 => x"1a",
          7990 => x"91",
          7991 => x"0b",
          7992 => x"80",
          7993 => x"0c",
          7994 => x"70",
          7995 => x"54",
          7996 => x"81",
          7997 => x"e0",
          7998 => x"2e",
          7999 => x"82",
          8000 => x"94",
          8001 => x"17",
          8002 => x"2b",
          8003 => x"57",
          8004 => x"52",
          8005 => x"e7",
          8006 => x"98",
          8007 => x"e0",
          8008 => x"26",
          8009 => x"55",
          8010 => x"08",
          8011 => x"81",
          8012 => x"79",
          8013 => x"31",
          8014 => x"70",
          8015 => x"25",
          8016 => x"76",
          8017 => x"81",
          8018 => x"55",
          8019 => x"38",
          8020 => x"0c",
          8021 => x"75",
          8022 => x"54",
          8023 => x"a2",
          8024 => x"7a",
          8025 => x"3f",
          8026 => x"08",
          8027 => x"55",
          8028 => x"89",
          8029 => x"98",
          8030 => x"1a",
          8031 => x"80",
          8032 => x"54",
          8033 => x"98",
          8034 => x"0d",
          8035 => x"0d",
          8036 => x"64",
          8037 => x"59",
          8038 => x"90",
          8039 => x"52",
          8040 => x"ce",
          8041 => x"98",
          8042 => x"e0",
          8043 => x"38",
          8044 => x"55",
          8045 => x"86",
          8046 => x"82",
          8047 => x"19",
          8048 => x"55",
          8049 => x"80",
          8050 => x"38",
          8051 => x"0b",
          8052 => x"82",
          8053 => x"39",
          8054 => x"1a",
          8055 => x"82",
          8056 => x"19",
          8057 => x"08",
          8058 => x"7c",
          8059 => x"74",
          8060 => x"2e",
          8061 => x"94",
          8062 => x"83",
          8063 => x"56",
          8064 => x"38",
          8065 => x"22",
          8066 => x"89",
          8067 => x"55",
          8068 => x"75",
          8069 => x"19",
          8070 => x"39",
          8071 => x"52",
          8072 => x"db",
          8073 => x"98",
          8074 => x"75",
          8075 => x"38",
          8076 => x"ff",
          8077 => x"98",
          8078 => x"19",
          8079 => x"51",
          8080 => x"82",
          8081 => x"80",
          8082 => x"38",
          8083 => x"08",
          8084 => x"2a",
          8085 => x"80",
          8086 => x"38",
          8087 => x"8a",
          8088 => x"5c",
          8089 => x"27",
          8090 => x"7a",
          8091 => x"54",
          8092 => x"52",
          8093 => x"51",
          8094 => x"3f",
          8095 => x"08",
          8096 => x"7e",
          8097 => x"56",
          8098 => x"2e",
          8099 => x"16",
          8100 => x"55",
          8101 => x"95",
          8102 => x"53",
          8103 => x"b4",
          8104 => x"31",
          8105 => x"05",
          8106 => x"e8",
          8107 => x"2b",
          8108 => x"76",
          8109 => x"94",
          8110 => x"ff",
          8111 => x"71",
          8112 => x"7b",
          8113 => x"38",
          8114 => x"19",
          8115 => x"51",
          8116 => x"82",
          8117 => x"fd",
          8118 => x"53",
          8119 => x"83",
          8120 => x"b8",
          8121 => x"51",
          8122 => x"3f",
          8123 => x"7e",
          8124 => x"0c",
          8125 => x"1b",
          8126 => x"1c",
          8127 => x"fd",
          8128 => x"56",
          8129 => x"98",
          8130 => x"0d",
          8131 => x"0d",
          8132 => x"64",
          8133 => x"58",
          8134 => x"90",
          8135 => x"52",
          8136 => x"ce",
          8137 => x"98",
          8138 => x"e0",
          8139 => x"38",
          8140 => x"55",
          8141 => x"86",
          8142 => x"83",
          8143 => x"18",
          8144 => x"2a",
          8145 => x"51",
          8146 => x"56",
          8147 => x"83",
          8148 => x"39",
          8149 => x"19",
          8150 => x"83",
          8151 => x"0b",
          8152 => x"81",
          8153 => x"39",
          8154 => x"7c",
          8155 => x"74",
          8156 => x"38",
          8157 => x"7b",
          8158 => x"f3",
          8159 => x"08",
          8160 => x"06",
          8161 => x"82",
          8162 => x"8a",
          8163 => x"05",
          8164 => x"06",
          8165 => x"bf",
          8166 => x"38",
          8167 => x"55",
          8168 => x"7a",
          8169 => x"98",
          8170 => x"77",
          8171 => x"3f",
          8172 => x"08",
          8173 => x"98",
          8174 => x"82",
          8175 => x"81",
          8176 => x"38",
          8177 => x"ff",
          8178 => x"98",
          8179 => x"18",
          8180 => x"74",
          8181 => x"7e",
          8182 => x"08",
          8183 => x"2e",
          8184 => x"8e",
          8185 => x"ff",
          8186 => x"82",
          8187 => x"fe",
          8188 => x"18",
          8189 => x"51",
          8190 => x"3f",
          8191 => x"08",
          8192 => x"d0",
          8193 => x"98",
          8194 => x"89",
          8195 => x"78",
          8196 => x"d7",
          8197 => x"7f",
          8198 => x"58",
          8199 => x"75",
          8200 => x"75",
          8201 => x"78",
          8202 => x"7c",
          8203 => x"33",
          8204 => x"c2",
          8205 => x"98",
          8206 => x"38",
          8207 => x"08",
          8208 => x"56",
          8209 => x"9c",
          8210 => x"53",
          8211 => x"77",
          8212 => x"7d",
          8213 => x"16",
          8214 => x"b8",
          8215 => x"80",
          8216 => x"34",
          8217 => x"56",
          8218 => x"8c",
          8219 => x"19",
          8220 => x"38",
          8221 => x"bb",
          8222 => x"e0",
          8223 => x"de",
          8224 => x"b4",
          8225 => x"76",
          8226 => x"94",
          8227 => x"ff",
          8228 => x"71",
          8229 => x"7b",
          8230 => x"38",
          8231 => x"18",
          8232 => x"51",
          8233 => x"3f",
          8234 => x"08",
          8235 => x"75",
          8236 => x"94",
          8237 => x"ff",
          8238 => x"05",
          8239 => x"d4",
          8240 => x"81",
          8241 => x"34",
          8242 => x"7e",
          8243 => x"0c",
          8244 => x"1a",
          8245 => x"94",
          8246 => x"1b",
          8247 => x"5e",
          8248 => x"27",
          8249 => x"55",
          8250 => x"0c",
          8251 => x"90",
          8252 => x"c0",
          8253 => x"90",
          8254 => x"56",
          8255 => x"98",
          8256 => x"0d",
          8257 => x"0d",
          8258 => x"fc",
          8259 => x"52",
          8260 => x"3f",
          8261 => x"08",
          8262 => x"98",
          8263 => x"38",
          8264 => x"70",
          8265 => x"81",
          8266 => x"55",
          8267 => x"80",
          8268 => x"16",
          8269 => x"51",
          8270 => x"3f",
          8271 => x"08",
          8272 => x"98",
          8273 => x"38",
          8274 => x"8b",
          8275 => x"07",
          8276 => x"8b",
          8277 => x"16",
          8278 => x"52",
          8279 => x"cc",
          8280 => x"16",
          8281 => x"15",
          8282 => x"f9",
          8283 => x"b2",
          8284 => x"15",
          8285 => x"ed",
          8286 => x"92",
          8287 => x"b7",
          8288 => x"54",
          8289 => x"15",
          8290 => x"ff",
          8291 => x"82",
          8292 => x"90",
          8293 => x"bf",
          8294 => x"73",
          8295 => x"76",
          8296 => x"0c",
          8297 => x"04",
          8298 => x"76",
          8299 => x"fe",
          8300 => x"e0",
          8301 => x"82",
          8302 => x"9c",
          8303 => x"fc",
          8304 => x"51",
          8305 => x"82",
          8306 => x"53",
          8307 => x"08",
          8308 => x"e0",
          8309 => x"0c",
          8310 => x"98",
          8311 => x"0d",
          8312 => x"0d",
          8313 => x"e6",
          8314 => x"52",
          8315 => x"e0",
          8316 => x"8b",
          8317 => x"98",
          8318 => x"f4",
          8319 => x"71",
          8320 => x"0c",
          8321 => x"04",
          8322 => x"80",
          8323 => x"cc",
          8324 => x"3d",
          8325 => x"3f",
          8326 => x"08",
          8327 => x"98",
          8328 => x"38",
          8329 => x"52",
          8330 => x"05",
          8331 => x"3f",
          8332 => x"08",
          8333 => x"98",
          8334 => x"02",
          8335 => x"33",
          8336 => x"55",
          8337 => x"25",
          8338 => x"7a",
          8339 => x"54",
          8340 => x"a2",
          8341 => x"84",
          8342 => x"06",
          8343 => x"73",
          8344 => x"38",
          8345 => x"70",
          8346 => x"e1",
          8347 => x"98",
          8348 => x"0c",
          8349 => x"e0",
          8350 => x"2e",
          8351 => x"83",
          8352 => x"74",
          8353 => x"0c",
          8354 => x"04",
          8355 => x"0d",
          8356 => x"08",
          8357 => x"08",
          8358 => x"7a",
          8359 => x"80",
          8360 => x"b4",
          8361 => x"e0",
          8362 => x"d1",
          8363 => x"98",
          8364 => x"e0",
          8365 => x"a1",
          8366 => x"d4",
          8367 => x"7c",
          8368 => x"80",
          8369 => x"55",
          8370 => x"3d",
          8371 => x"80",
          8372 => x"38",
          8373 => x"d3",
          8374 => x"55",
          8375 => x"82",
          8376 => x"57",
          8377 => x"08",
          8378 => x"80",
          8379 => x"52",
          8380 => x"b7",
          8381 => x"e0",
          8382 => x"82",
          8383 => x"82",
          8384 => x"da",
          8385 => x"7b",
          8386 => x"3f",
          8387 => x"08",
          8388 => x"0c",
          8389 => x"51",
          8390 => x"82",
          8391 => x"57",
          8392 => x"08",
          8393 => x"80",
          8394 => x"c9",
          8395 => x"e0",
          8396 => x"82",
          8397 => x"a7",
          8398 => x"3d",
          8399 => x"51",
          8400 => x"73",
          8401 => x"08",
          8402 => x"76",
          8403 => x"c4",
          8404 => x"e0",
          8405 => x"82",
          8406 => x"80",
          8407 => x"76",
          8408 => x"81",
          8409 => x"82",
          8410 => x"39",
          8411 => x"38",
          8412 => x"fd",
          8413 => x"74",
          8414 => x"3f",
          8415 => x"78",
          8416 => x"33",
          8417 => x"56",
          8418 => x"92",
          8419 => x"c6",
          8420 => x"16",
          8421 => x"33",
          8422 => x"73",
          8423 => x"16",
          8424 => x"26",
          8425 => x"75",
          8426 => x"38",
          8427 => x"05",
          8428 => x"80",
          8429 => x"11",
          8430 => x"18",
          8431 => x"58",
          8432 => x"34",
          8433 => x"ff",
          8434 => x"3d",
          8435 => x"58",
          8436 => x"fd",
          8437 => x"7b",
          8438 => x"06",
          8439 => x"18",
          8440 => x"08",
          8441 => x"af",
          8442 => x"0b",
          8443 => x"33",
          8444 => x"82",
          8445 => x"70",
          8446 => x"52",
          8447 => x"56",
          8448 => x"8d",
          8449 => x"70",
          8450 => x"51",
          8451 => x"f5",
          8452 => x"54",
          8453 => x"a7",
          8454 => x"74",
          8455 => x"38",
          8456 => x"73",
          8457 => x"81",
          8458 => x"81",
          8459 => x"39",
          8460 => x"81",
          8461 => x"74",
          8462 => x"81",
          8463 => x"91",
          8464 => x"80",
          8465 => x"18",
          8466 => x"54",
          8467 => x"70",
          8468 => x"34",
          8469 => x"eb",
          8470 => x"34",
          8471 => x"98",
          8472 => x"3d",
          8473 => x"3d",
          8474 => x"8d",
          8475 => x"54",
          8476 => x"55",
          8477 => x"82",
          8478 => x"53",
          8479 => x"08",
          8480 => x"91",
          8481 => x"72",
          8482 => x"8c",
          8483 => x"73",
          8484 => x"38",
          8485 => x"70",
          8486 => x"81",
          8487 => x"57",
          8488 => x"73",
          8489 => x"08",
          8490 => x"94",
          8491 => x"75",
          8492 => x"9b",
          8493 => x"11",
          8494 => x"2b",
          8495 => x"73",
          8496 => x"38",
          8497 => x"16",
          8498 => x"88",
          8499 => x"98",
          8500 => x"78",
          8501 => x"55",
          8502 => x"f8",
          8503 => x"98",
          8504 => x"96",
          8505 => x"70",
          8506 => x"94",
          8507 => x"71",
          8508 => x"08",
          8509 => x"53",
          8510 => x"15",
          8511 => x"a7",
          8512 => x"74",
          8513 => x"d3",
          8514 => x"98",
          8515 => x"e0",
          8516 => x"2e",
          8517 => x"82",
          8518 => x"ff",
          8519 => x"38",
          8520 => x"08",
          8521 => x"73",
          8522 => x"73",
          8523 => x"9f",
          8524 => x"27",
          8525 => x"75",
          8526 => x"16",
          8527 => x"17",
          8528 => x"33",
          8529 => x"70",
          8530 => x"55",
          8531 => x"80",
          8532 => x"73",
          8533 => x"ff",
          8534 => x"82",
          8535 => x"54",
          8536 => x"08",
          8537 => x"e0",
          8538 => x"a8",
          8539 => x"74",
          8540 => x"8b",
          8541 => x"98",
          8542 => x"ff",
          8543 => x"81",
          8544 => x"38",
          8545 => x"9c",
          8546 => x"a7",
          8547 => x"16",
          8548 => x"39",
          8549 => x"16",
          8550 => x"75",
          8551 => x"53",
          8552 => x"ab",
          8553 => x"79",
          8554 => x"a9",
          8555 => x"98",
          8556 => x"82",
          8557 => x"34",
          8558 => x"c4",
          8559 => x"91",
          8560 => x"53",
          8561 => x"89",
          8562 => x"98",
          8563 => x"94",
          8564 => x"8c",
          8565 => x"27",
          8566 => x"8c",
          8567 => x"15",
          8568 => x"07",
          8569 => x"16",
          8570 => x"ff",
          8571 => x"80",
          8572 => x"77",
          8573 => x"2e",
          8574 => x"9c",
          8575 => x"53",
          8576 => x"98",
          8577 => x"0d",
          8578 => x"0d",
          8579 => x"54",
          8580 => x"81",
          8581 => x"53",
          8582 => x"05",
          8583 => x"84",
          8584 => x"d9",
          8585 => x"98",
          8586 => x"e0",
          8587 => x"eb",
          8588 => x"0c",
          8589 => x"51",
          8590 => x"82",
          8591 => x"55",
          8592 => x"08",
          8593 => x"ab",
          8594 => x"98",
          8595 => x"80",
          8596 => x"38",
          8597 => x"70",
          8598 => x"81",
          8599 => x"57",
          8600 => x"ae",
          8601 => x"08",
          8602 => x"c1",
          8603 => x"e0",
          8604 => x"17",
          8605 => x"86",
          8606 => x"17",
          8607 => x"75",
          8608 => x"ea",
          8609 => x"98",
          8610 => x"84",
          8611 => x"06",
          8612 => x"55",
          8613 => x"80",
          8614 => x"80",
          8615 => x"54",
          8616 => x"98",
          8617 => x"0d",
          8618 => x"0d",
          8619 => x"fc",
          8620 => x"52",
          8621 => x"3f",
          8622 => x"08",
          8623 => x"e0",
          8624 => x"0c",
          8625 => x"04",
          8626 => x"77",
          8627 => x"fc",
          8628 => x"53",
          8629 => x"9a",
          8630 => x"98",
          8631 => x"e0",
          8632 => x"e1",
          8633 => x"38",
          8634 => x"08",
          8635 => x"ff",
          8636 => x"82",
          8637 => x"53",
          8638 => x"82",
          8639 => x"52",
          8640 => x"df",
          8641 => x"98",
          8642 => x"e0",
          8643 => x"2e",
          8644 => x"85",
          8645 => x"87",
          8646 => x"98",
          8647 => x"74",
          8648 => x"ce",
          8649 => x"52",
          8650 => x"bd",
          8651 => x"e0",
          8652 => x"32",
          8653 => x"72",
          8654 => x"70",
          8655 => x"08",
          8656 => x"54",
          8657 => x"e0",
          8658 => x"3d",
          8659 => x"3d",
          8660 => x"80",
          8661 => x"70",
          8662 => x"52",
          8663 => x"3f",
          8664 => x"08",
          8665 => x"98",
          8666 => x"65",
          8667 => x"d2",
          8668 => x"e0",
          8669 => x"82",
          8670 => x"a0",
          8671 => x"cb",
          8672 => x"98",
          8673 => x"73",
          8674 => x"38",
          8675 => x"39",
          8676 => x"88",
          8677 => x"75",
          8678 => x"3f",
          8679 => x"98",
          8680 => x"0d",
          8681 => x"0d",
          8682 => x"5c",
          8683 => x"3d",
          8684 => x"93",
          8685 => x"c5",
          8686 => x"98",
          8687 => x"e0",
          8688 => x"82",
          8689 => x"0c",
          8690 => x"11",
          8691 => x"94",
          8692 => x"56",
          8693 => x"74",
          8694 => x"75",
          8695 => x"e6",
          8696 => x"81",
          8697 => x"5b",
          8698 => x"82",
          8699 => x"75",
          8700 => x"73",
          8701 => x"81",
          8702 => x"38",
          8703 => x"57",
          8704 => x"3d",
          8705 => x"ff",
          8706 => x"82",
          8707 => x"ff",
          8708 => x"82",
          8709 => x"81",
          8710 => x"82",
          8711 => x"30",
          8712 => x"98",
          8713 => x"25",
          8714 => x"19",
          8715 => x"5a",
          8716 => x"08",
          8717 => x"38",
          8718 => x"a8",
          8719 => x"e0",
          8720 => x"58",
          8721 => x"77",
          8722 => x"7d",
          8723 => x"ad",
          8724 => x"e0",
          8725 => x"82",
          8726 => x"80",
          8727 => x"70",
          8728 => x"ff",
          8729 => x"56",
          8730 => x"2e",
          8731 => x"9e",
          8732 => x"51",
          8733 => x"3f",
          8734 => x"08",
          8735 => x"06",
          8736 => x"80",
          8737 => x"19",
          8738 => x"54",
          8739 => x"14",
          8740 => x"88",
          8741 => x"98",
          8742 => x"06",
          8743 => x"80",
          8744 => x"19",
          8745 => x"54",
          8746 => x"06",
          8747 => x"79",
          8748 => x"78",
          8749 => x"79",
          8750 => x"84",
          8751 => x"07",
          8752 => x"84",
          8753 => x"82",
          8754 => x"92",
          8755 => x"f9",
          8756 => x"8a",
          8757 => x"53",
          8758 => x"e3",
          8759 => x"e0",
          8760 => x"82",
          8761 => x"81",
          8762 => x"17",
          8763 => x"81",
          8764 => x"17",
          8765 => x"2a",
          8766 => x"51",
          8767 => x"55",
          8768 => x"81",
          8769 => x"17",
          8770 => x"8c",
          8771 => x"81",
          8772 => x"9c",
          8773 => x"98",
          8774 => x"17",
          8775 => x"51",
          8776 => x"3f",
          8777 => x"08",
          8778 => x"0c",
          8779 => x"39",
          8780 => x"52",
          8781 => x"ad",
          8782 => x"e0",
          8783 => x"2e",
          8784 => x"83",
          8785 => x"82",
          8786 => x"81",
          8787 => x"06",
          8788 => x"56",
          8789 => x"a1",
          8790 => x"82",
          8791 => x"9c",
          8792 => x"95",
          8793 => x"08",
          8794 => x"98",
          8795 => x"51",
          8796 => x"3f",
          8797 => x"08",
          8798 => x"08",
          8799 => x"90",
          8800 => x"c0",
          8801 => x"90",
          8802 => x"80",
          8803 => x"75",
          8804 => x"75",
          8805 => x"e0",
          8806 => x"3d",
          8807 => x"3d",
          8808 => x"a2",
          8809 => x"05",
          8810 => x"51",
          8811 => x"82",
          8812 => x"55",
          8813 => x"08",
          8814 => x"78",
          8815 => x"08",
          8816 => x"70",
          8817 => x"cf",
          8818 => x"98",
          8819 => x"e0",
          8820 => x"df",
          8821 => x"ff",
          8822 => x"85",
          8823 => x"06",
          8824 => x"86",
          8825 => x"cb",
          8826 => x"2b",
          8827 => x"24",
          8828 => x"02",
          8829 => x"33",
          8830 => x"58",
          8831 => x"76",
          8832 => x"6c",
          8833 => x"ff",
          8834 => x"82",
          8835 => x"74",
          8836 => x"81",
          8837 => x"56",
          8838 => x"80",
          8839 => x"54",
          8840 => x"08",
          8841 => x"2e",
          8842 => x"73",
          8843 => x"98",
          8844 => x"52",
          8845 => x"52",
          8846 => x"b2",
          8847 => x"98",
          8848 => x"e0",
          8849 => x"eb",
          8850 => x"98",
          8851 => x"51",
          8852 => x"3f",
          8853 => x"08",
          8854 => x"98",
          8855 => x"87",
          8856 => x"39",
          8857 => x"08",
          8858 => x"38",
          8859 => x"08",
          8860 => x"77",
          8861 => x"3f",
          8862 => x"08",
          8863 => x"08",
          8864 => x"e0",
          8865 => x"80",
          8866 => x"55",
          8867 => x"95",
          8868 => x"2e",
          8869 => x"53",
          8870 => x"51",
          8871 => x"3f",
          8872 => x"08",
          8873 => x"38",
          8874 => x"a8",
          8875 => x"e0",
          8876 => x"74",
          8877 => x"0c",
          8878 => x"04",
          8879 => x"82",
          8880 => x"ff",
          8881 => x"9b",
          8882 => x"b1",
          8883 => x"98",
          8884 => x"e0",
          8885 => x"b7",
          8886 => x"6a",
          8887 => x"70",
          8888 => x"b3",
          8889 => x"98",
          8890 => x"e0",
          8891 => x"38",
          8892 => x"9b",
          8893 => x"98",
          8894 => x"09",
          8895 => x"8f",
          8896 => x"df",
          8897 => x"85",
          8898 => x"51",
          8899 => x"74",
          8900 => x"78",
          8901 => x"8a",
          8902 => x"57",
          8903 => x"3f",
          8904 => x"08",
          8905 => x"82",
          8906 => x"83",
          8907 => x"82",
          8908 => x"81",
          8909 => x"06",
          8910 => x"54",
          8911 => x"08",
          8912 => x"81",
          8913 => x"81",
          8914 => x"39",
          8915 => x"38",
          8916 => x"08",
          8917 => x"ff",
          8918 => x"82",
          8919 => x"54",
          8920 => x"08",
          8921 => x"8b",
          8922 => x"b8",
          8923 => x"a4",
          8924 => x"54",
          8925 => x"15",
          8926 => x"90",
          8927 => x"15",
          8928 => x"b2",
          8929 => x"ce",
          8930 => x"a3",
          8931 => x"53",
          8932 => x"53",
          8933 => x"ee",
          8934 => x"78",
          8935 => x"80",
          8936 => x"ff",
          8937 => x"78",
          8938 => x"80",
          8939 => x"7f",
          8940 => x"d8",
          8941 => x"ff",
          8942 => x"78",
          8943 => x"83",
          8944 => x"51",
          8945 => x"3f",
          8946 => x"08",
          8947 => x"98",
          8948 => x"82",
          8949 => x"52",
          8950 => x"51",
          8951 => x"3f",
          8952 => x"52",
          8953 => x"b7",
          8954 => x"54",
          8955 => x"15",
          8956 => x"81",
          8957 => x"34",
          8958 => x"a6",
          8959 => x"e0",
          8960 => x"8b",
          8961 => x"75",
          8962 => x"ff",
          8963 => x"73",
          8964 => x"0c",
          8965 => x"04",
          8966 => x"ab",
          8967 => x"51",
          8968 => x"82",
          8969 => x"fe",
          8970 => x"ab",
          8971 => x"cd",
          8972 => x"98",
          8973 => x"e0",
          8974 => x"d8",
          8975 => x"ab",
          8976 => x"9e",
          8977 => x"58",
          8978 => x"82",
          8979 => x"55",
          8980 => x"08",
          8981 => x"02",
          8982 => x"33",
          8983 => x"54",
          8984 => x"82",
          8985 => x"53",
          8986 => x"52",
          8987 => x"80",
          8988 => x"a2",
          8989 => x"53",
          8990 => x"3d",
          8991 => x"ff",
          8992 => x"ac",
          8993 => x"73",
          8994 => x"3f",
          8995 => x"08",
          8996 => x"98",
          8997 => x"63",
          8998 => x"2e",
          8999 => x"88",
          9000 => x"3d",
          9001 => x"38",
          9002 => x"e8",
          9003 => x"98",
          9004 => x"09",
          9005 => x"bb",
          9006 => x"ff",
          9007 => x"82",
          9008 => x"55",
          9009 => x"08",
          9010 => x"68",
          9011 => x"aa",
          9012 => x"05",
          9013 => x"51",
          9014 => x"3f",
          9015 => x"33",
          9016 => x"8b",
          9017 => x"84",
          9018 => x"06",
          9019 => x"73",
          9020 => x"a0",
          9021 => x"8b",
          9022 => x"54",
          9023 => x"15",
          9024 => x"33",
          9025 => x"70",
          9026 => x"55",
          9027 => x"2e",
          9028 => x"6f",
          9029 => x"e1",
          9030 => x"78",
          9031 => x"ad",
          9032 => x"98",
          9033 => x"51",
          9034 => x"3f",
          9035 => x"e0",
          9036 => x"2e",
          9037 => x"82",
          9038 => x"52",
          9039 => x"a3",
          9040 => x"e0",
          9041 => x"80",
          9042 => x"58",
          9043 => x"98",
          9044 => x"38",
          9045 => x"54",
          9046 => x"09",
          9047 => x"38",
          9048 => x"52",
          9049 => x"b4",
          9050 => x"54",
          9051 => x"15",
          9052 => x"82",
          9053 => x"9c",
          9054 => x"c1",
          9055 => x"e0",
          9056 => x"82",
          9057 => x"8c",
          9058 => x"ff",
          9059 => x"82",
          9060 => x"55",
          9061 => x"98",
          9062 => x"0d",
          9063 => x"0d",
          9064 => x"05",
          9065 => x"05",
          9066 => x"33",
          9067 => x"53",
          9068 => x"05",
          9069 => x"51",
          9070 => x"82",
          9071 => x"55",
          9072 => x"08",
          9073 => x"78",
          9074 => x"96",
          9075 => x"51",
          9076 => x"82",
          9077 => x"55",
          9078 => x"08",
          9079 => x"80",
          9080 => x"81",
          9081 => x"86",
          9082 => x"38",
          9083 => x"61",
          9084 => x"12",
          9085 => x"7a",
          9086 => x"51",
          9087 => x"74",
          9088 => x"78",
          9089 => x"83",
          9090 => x"51",
          9091 => x"3f",
          9092 => x"08",
          9093 => x"e0",
          9094 => x"3d",
          9095 => x"3d",
          9096 => x"82",
          9097 => x"cc",
          9098 => x"3d",
          9099 => x"3f",
          9100 => x"08",
          9101 => x"98",
          9102 => x"38",
          9103 => x"52",
          9104 => x"05",
          9105 => x"3f",
          9106 => x"08",
          9107 => x"98",
          9108 => x"02",
          9109 => x"33",
          9110 => x"54",
          9111 => x"a6",
          9112 => x"22",
          9113 => x"71",
          9114 => x"53",
          9115 => x"51",
          9116 => x"3f",
          9117 => x"0b",
          9118 => x"76",
          9119 => x"a6",
          9120 => x"98",
          9121 => x"82",
          9122 => x"94",
          9123 => x"e9",
          9124 => x"6c",
          9125 => x"53",
          9126 => x"05",
          9127 => x"51",
          9128 => x"82",
          9129 => x"82",
          9130 => x"30",
          9131 => x"98",
          9132 => x"25",
          9133 => x"79",
          9134 => x"86",
          9135 => x"75",
          9136 => x"73",
          9137 => x"fa",
          9138 => x"80",
          9139 => x"8d",
          9140 => x"54",
          9141 => x"3f",
          9142 => x"08",
          9143 => x"98",
          9144 => x"38",
          9145 => x"51",
          9146 => x"3f",
          9147 => x"08",
          9148 => x"98",
          9149 => x"82",
          9150 => x"82",
          9151 => x"65",
          9152 => x"78",
          9153 => x"7b",
          9154 => x"55",
          9155 => x"34",
          9156 => x"8a",
          9157 => x"38",
          9158 => x"1a",
          9159 => x"34",
          9160 => x"9e",
          9161 => x"70",
          9162 => x"51",
          9163 => x"a0",
          9164 => x"8e",
          9165 => x"2e",
          9166 => x"86",
          9167 => x"34",
          9168 => x"30",
          9169 => x"80",
          9170 => x"7a",
          9171 => x"c1",
          9172 => x"2e",
          9173 => x"a4",
          9174 => x"51",
          9175 => x"3f",
          9176 => x"08",
          9177 => x"98",
          9178 => x"7b",
          9179 => x"55",
          9180 => x"73",
          9181 => x"38",
          9182 => x"73",
          9183 => x"38",
          9184 => x"15",
          9185 => x"ff",
          9186 => x"82",
          9187 => x"7b",
          9188 => x"e0",
          9189 => x"3d",
          9190 => x"3d",
          9191 => x"9c",
          9192 => x"05",
          9193 => x"51",
          9194 => x"82",
          9195 => x"82",
          9196 => x"56",
          9197 => x"98",
          9198 => x"38",
          9199 => x"52",
          9200 => x"52",
          9201 => x"ef",
          9202 => x"70",
          9203 => x"56",
          9204 => x"81",
          9205 => x"57",
          9206 => x"ff",
          9207 => x"82",
          9208 => x"83",
          9209 => x"80",
          9210 => x"e0",
          9211 => x"96",
          9212 => x"b5",
          9213 => x"98",
          9214 => x"90",
          9215 => x"98",
          9216 => x"ff",
          9217 => x"80",
          9218 => x"74",
          9219 => x"b8",
          9220 => x"ee",
          9221 => x"98",
          9222 => x"81",
          9223 => x"88",
          9224 => x"26",
          9225 => x"39",
          9226 => x"86",
          9227 => x"81",
          9228 => x"ff",
          9229 => x"38",
          9230 => x"54",
          9231 => x"81",
          9232 => x"81",
          9233 => x"77",
          9234 => x"59",
          9235 => x"6d",
          9236 => x"55",
          9237 => x"26",
          9238 => x"8a",
          9239 => x"86",
          9240 => x"e5",
          9241 => x"38",
          9242 => x"99",
          9243 => x"05",
          9244 => x"70",
          9245 => x"73",
          9246 => x"81",
          9247 => x"ff",
          9248 => x"ed",
          9249 => x"80",
          9250 => x"90",
          9251 => x"55",
          9252 => x"3f",
          9253 => x"08",
          9254 => x"98",
          9255 => x"38",
          9256 => x"51",
          9257 => x"3f",
          9258 => x"08",
          9259 => x"98",
          9260 => x"75",
          9261 => x"66",
          9262 => x"34",
          9263 => x"82",
          9264 => x"84",
          9265 => x"06",
          9266 => x"80",
          9267 => x"2e",
          9268 => x"81",
          9269 => x"ff",
          9270 => x"82",
          9271 => x"54",
          9272 => x"08",
          9273 => x"53",
          9274 => x"08",
          9275 => x"ff",
          9276 => x"66",
          9277 => x"8b",
          9278 => x"53",
          9279 => x"51",
          9280 => x"3f",
          9281 => x"0b",
          9282 => x"78",
          9283 => x"96",
          9284 => x"98",
          9285 => x"55",
          9286 => x"98",
          9287 => x"0d",
          9288 => x"0d",
          9289 => x"88",
          9290 => x"05",
          9291 => x"fc",
          9292 => x"54",
          9293 => x"d2",
          9294 => x"e0",
          9295 => x"82",
          9296 => x"82",
          9297 => x"1a",
          9298 => x"82",
          9299 => x"80",
          9300 => x"8c",
          9301 => x"78",
          9302 => x"1a",
          9303 => x"2a",
          9304 => x"51",
          9305 => x"90",
          9306 => x"82",
          9307 => x"58",
          9308 => x"81",
          9309 => x"39",
          9310 => x"22",
          9311 => x"70",
          9312 => x"56",
          9313 => x"a2",
          9314 => x"14",
          9315 => x"30",
          9316 => x"9f",
          9317 => x"98",
          9318 => x"19",
          9319 => x"5a",
          9320 => x"81",
          9321 => x"38",
          9322 => x"77",
          9323 => x"82",
          9324 => x"56",
          9325 => x"74",
          9326 => x"ff",
          9327 => x"81",
          9328 => x"55",
          9329 => x"75",
          9330 => x"82",
          9331 => x"98",
          9332 => x"ff",
          9333 => x"e0",
          9334 => x"2e",
          9335 => x"82",
          9336 => x"8e",
          9337 => x"56",
          9338 => x"09",
          9339 => x"38",
          9340 => x"59",
          9341 => x"77",
          9342 => x"06",
          9343 => x"87",
          9344 => x"39",
          9345 => x"ba",
          9346 => x"55",
          9347 => x"2e",
          9348 => x"15",
          9349 => x"2e",
          9350 => x"83",
          9351 => x"75",
          9352 => x"7e",
          9353 => x"d0",
          9354 => x"98",
          9355 => x"e0",
          9356 => x"ce",
          9357 => x"16",
          9358 => x"56",
          9359 => x"38",
          9360 => x"19",
          9361 => x"90",
          9362 => x"7d",
          9363 => x"38",
          9364 => x"0c",
          9365 => x"0c",
          9366 => x"80",
          9367 => x"73",
          9368 => x"9c",
          9369 => x"05",
          9370 => x"57",
          9371 => x"26",
          9372 => x"7b",
          9373 => x"0c",
          9374 => x"81",
          9375 => x"84",
          9376 => x"54",
          9377 => x"98",
          9378 => x"0d",
          9379 => x"0d",
          9380 => x"88",
          9381 => x"05",
          9382 => x"54",
          9383 => x"c4",
          9384 => x"56",
          9385 => x"e0",
          9386 => x"8d",
          9387 => x"e0",
          9388 => x"29",
          9389 => x"05",
          9390 => x"55",
          9391 => x"84",
          9392 => x"34",
          9393 => x"08",
          9394 => x"08",
          9395 => x"8c",
          9396 => x"e0",
          9397 => x"47",
          9398 => x"52",
          9399 => x"8e",
          9400 => x"e0",
          9401 => x"ff",
          9402 => x"06",
          9403 => x"56",
          9404 => x"38",
          9405 => x"70",
          9406 => x"55",
          9407 => x"8c",
          9408 => x"3d",
          9409 => x"83",
          9410 => x"ff",
          9411 => x"82",
          9412 => x"99",
          9413 => x"74",
          9414 => x"38",
          9415 => x"80",
          9416 => x"ff",
          9417 => x"55",
          9418 => x"83",
          9419 => x"78",
          9420 => x"38",
          9421 => x"26",
          9422 => x"81",
          9423 => x"8b",
          9424 => x"79",
          9425 => x"80",
          9426 => x"93",
          9427 => x"39",
          9428 => x"6f",
          9429 => x"89",
          9430 => x"49",
          9431 => x"83",
          9432 => x"61",
          9433 => x"25",
          9434 => x"55",
          9435 => x"8b",
          9436 => x"80",
          9437 => x"38",
          9438 => x"53",
          9439 => x"51",
          9440 => x"3f",
          9441 => x"e0",
          9442 => x"c1",
          9443 => x"1b",
          9444 => x"f1",
          9445 => x"98",
          9446 => x"ff",
          9447 => x"56",
          9448 => x"d5",
          9449 => x"06",
          9450 => x"64",
          9451 => x"83",
          9452 => x"56",
          9453 => x"2e",
          9454 => x"83",
          9455 => x"ff",
          9456 => x"82",
          9457 => x"83",
          9458 => x"5f",
          9459 => x"3f",
          9460 => x"08",
          9461 => x"9a",
          9462 => x"53",
          9463 => x"51",
          9464 => x"3f",
          9465 => x"e0",
          9466 => x"e1",
          9467 => x"2a",
          9468 => x"82",
          9469 => x"41",
          9470 => x"83",
          9471 => x"67",
          9472 => x"7e",
          9473 => x"c5",
          9474 => x"31",
          9475 => x"80",
          9476 => x"8a",
          9477 => x"56",
          9478 => x"26",
          9479 => x"62",
          9480 => x"81",
          9481 => x"74",
          9482 => x"38",
          9483 => x"55",
          9484 => x"83",
          9485 => x"81",
          9486 => x"80",
          9487 => x"38",
          9488 => x"55",
          9489 => x"5e",
          9490 => x"8a",
          9491 => x"5a",
          9492 => x"09",
          9493 => x"e1",
          9494 => x"38",
          9495 => x"57",
          9496 => x"d3",
          9497 => x"5a",
          9498 => x"9d",
          9499 => x"26",
          9500 => x"d3",
          9501 => x"10",
          9502 => x"22",
          9503 => x"74",
          9504 => x"38",
          9505 => x"ee",
          9506 => x"67",
          9507 => x"c4",
          9508 => x"98",
          9509 => x"84",
          9510 => x"89",
          9511 => x"a0",
          9512 => x"82",
          9513 => x"fc",
          9514 => x"56",
          9515 => x"f0",
          9516 => x"80",
          9517 => x"88",
          9518 => x"38",
          9519 => x"57",
          9520 => x"d3",
          9521 => x"5a",
          9522 => x"9d",
          9523 => x"26",
          9524 => x"d3",
          9525 => x"10",
          9526 => x"22",
          9527 => x"74",
          9528 => x"38",
          9529 => x"ee",
          9530 => x"67",
          9531 => x"e4",
          9532 => x"98",
          9533 => x"05",
          9534 => x"98",
          9535 => x"26",
          9536 => x"0b",
          9537 => x"08",
          9538 => x"98",
          9539 => x"11",
          9540 => x"05",
          9541 => x"83",
          9542 => x"2a",
          9543 => x"a0",
          9544 => x"7d",
          9545 => x"6a",
          9546 => x"05",
          9547 => x"72",
          9548 => x"5c",
          9549 => x"59",
          9550 => x"2e",
          9551 => x"89",
          9552 => x"61",
          9553 => x"84",
          9554 => x"5d",
          9555 => x"18",
          9556 => x"69",
          9557 => x"74",
          9558 => x"e4",
          9559 => x"31",
          9560 => x"53",
          9561 => x"52",
          9562 => x"e8",
          9563 => x"98",
          9564 => x"83",
          9565 => x"06",
          9566 => x"e0",
          9567 => x"ff",
          9568 => x"dd",
          9569 => x"b8",
          9570 => x"2a",
          9571 => x"be",
          9572 => x"39",
          9573 => x"09",
          9574 => x"c5",
          9575 => x"f5",
          9576 => x"98",
          9577 => x"38",
          9578 => x"79",
          9579 => x"80",
          9580 => x"38",
          9581 => x"96",
          9582 => x"06",
          9583 => x"2e",
          9584 => x"5e",
          9585 => x"82",
          9586 => x"9f",
          9587 => x"38",
          9588 => x"38",
          9589 => x"81",
          9590 => x"fc",
          9591 => x"e0",
          9592 => x"7d",
          9593 => x"81",
          9594 => x"7d",
          9595 => x"78",
          9596 => x"74",
          9597 => x"8e",
          9598 => x"d1",
          9599 => x"53",
          9600 => x"51",
          9601 => x"3f",
          9602 => x"d1",
          9603 => x"51",
          9604 => x"3f",
          9605 => x"8b",
          9606 => x"8e",
          9607 => x"8d",
          9608 => x"83",
          9609 => x"52",
          9610 => x"ff",
          9611 => x"81",
          9612 => x"34",
          9613 => x"70",
          9614 => x"2a",
          9615 => x"54",
          9616 => x"1b",
          9617 => x"ff",
          9618 => x"74",
          9619 => x"26",
          9620 => x"83",
          9621 => x"52",
          9622 => x"ff",
          9623 => x"8a",
          9624 => x"a0",
          9625 => x"8d",
          9626 => x"0b",
          9627 => x"bf",
          9628 => x"51",
          9629 => x"3f",
          9630 => x"9a",
          9631 => x"8d",
          9632 => x"52",
          9633 => x"ff",
          9634 => x"7d",
          9635 => x"81",
          9636 => x"38",
          9637 => x"0a",
          9638 => x"1b",
          9639 => x"c5",
          9640 => x"a4",
          9641 => x"8d",
          9642 => x"52",
          9643 => x"ff",
          9644 => x"81",
          9645 => x"51",
          9646 => x"3f",
          9647 => x"1b",
          9648 => x"83",
          9649 => x"0b",
          9650 => x"34",
          9651 => x"c2",
          9652 => x"53",
          9653 => x"52",
          9654 => x"51",
          9655 => x"88",
          9656 => x"a7",
          9657 => x"8c",
          9658 => x"83",
          9659 => x"52",
          9660 => x"ff",
          9661 => x"ff",
          9662 => x"1c",
          9663 => x"a6",
          9664 => x"53",
          9665 => x"52",
          9666 => x"ff",
          9667 => x"82",
          9668 => x"83",
          9669 => x"52",
          9670 => x"ab",
          9671 => x"7e",
          9672 => x"7f",
          9673 => x"ce",
          9674 => x"82",
          9675 => x"84",
          9676 => x"83",
          9677 => x"06",
          9678 => x"75",
          9679 => x"53",
          9680 => x"51",
          9681 => x"3f",
          9682 => x"80",
          9683 => x"ff",
          9684 => x"84",
          9685 => x"d2",
          9686 => x"ff",
          9687 => x"86",
          9688 => x"f2",
          9689 => x"1b",
          9690 => x"f9",
          9691 => x"52",
          9692 => x"51",
          9693 => x"3f",
          9694 => x"ec",
          9695 => x"8b",
          9696 => x"d4",
          9697 => x"51",
          9698 => x"3f",
          9699 => x"1f",
          9700 => x"7f",
          9701 => x"de",
          9702 => x"75",
          9703 => x"52",
          9704 => x"87",
          9705 => x"53",
          9706 => x"51",
          9707 => x"3f",
          9708 => x"58",
          9709 => x"09",
          9710 => x"38",
          9711 => x"51",
          9712 => x"3f",
          9713 => x"1b",
          9714 => x"99",
          9715 => x"52",
          9716 => x"91",
          9717 => x"ff",
          9718 => x"81",
          9719 => x"f8",
          9720 => x"7a",
          9721 => x"fd",
          9722 => x"61",
          9723 => x"26",
          9724 => x"57",
          9725 => x"53",
          9726 => x"51",
          9727 => x"3f",
          9728 => x"08",
          9729 => x"84",
          9730 => x"e0",
          9731 => x"7a",
          9732 => x"a3",
          9733 => x"75",
          9734 => x"56",
          9735 => x"81",
          9736 => x"80",
          9737 => x"38",
          9738 => x"83",
          9739 => x"65",
          9740 => x"74",
          9741 => x"38",
          9742 => x"54",
          9743 => x"52",
          9744 => x"86",
          9745 => x"e0",
          9746 => x"f8",
          9747 => x"75",
          9748 => x"56",
          9749 => x"8c",
          9750 => x"2e",
          9751 => x"57",
          9752 => x"ff",
          9753 => x"84",
          9754 => x"2e",
          9755 => x"57",
          9756 => x"b2",
          9757 => x"80",
          9758 => x"7f",
          9759 => x"8c",
          9760 => x"82",
          9761 => x"81",
          9762 => x"90",
          9763 => x"76",
          9764 => x"34",
          9765 => x"e0",
          9766 => x"7a",
          9767 => x"ff",
          9768 => x"81",
          9769 => x"83",
          9770 => x"58",
          9771 => x"38",
          9772 => x"77",
          9773 => x"ff",
          9774 => x"82",
          9775 => x"78",
          9776 => x"83",
          9777 => x"1b",
          9778 => x"34",
          9779 => x"16",
          9780 => x"82",
          9781 => x"83",
          9782 => x"84",
          9783 => x"1f",
          9784 => x"c1",
          9785 => x"fe",
          9786 => x"fe",
          9787 => x"34",
          9788 => x"08",
          9789 => x"07",
          9790 => x"16",
          9791 => x"98",
          9792 => x"34",
          9793 => x"c6",
          9794 => x"88",
          9795 => x"52",
          9796 => x"51",
          9797 => x"3f",
          9798 => x"53",
          9799 => x"51",
          9800 => x"3f",
          9801 => x"e0",
          9802 => x"38",
          9803 => x"52",
          9804 => x"86",
          9805 => x"56",
          9806 => x"08",
          9807 => x"39",
          9808 => x"39",
          9809 => x"39",
          9810 => x"08",
          9811 => x"e0",
          9812 => x"3d",
          9813 => x"3d",
          9814 => x"5b",
          9815 => x"60",
          9816 => x"57",
          9817 => x"25",
          9818 => x"3d",
          9819 => x"55",
          9820 => x"15",
          9821 => x"c8",
          9822 => x"81",
          9823 => x"06",
          9824 => x"3d",
          9825 => x"8d",
          9826 => x"74",
          9827 => x"05",
          9828 => x"17",
          9829 => x"2e",
          9830 => x"c9",
          9831 => x"34",
          9832 => x"83",
          9833 => x"74",
          9834 => x"0c",
          9835 => x"04",
          9836 => x"7b",
          9837 => x"b3",
          9838 => x"57",
          9839 => x"09",
          9840 => x"38",
          9841 => x"51",
          9842 => x"17",
          9843 => x"76",
          9844 => x"88",
          9845 => x"17",
          9846 => x"59",
          9847 => x"81",
          9848 => x"76",
          9849 => x"8b",
          9850 => x"54",
          9851 => x"17",
          9852 => x"51",
          9853 => x"79",
          9854 => x"30",
          9855 => x"9f",
          9856 => x"53",
          9857 => x"75",
          9858 => x"81",
          9859 => x"0c",
          9860 => x"04",
          9861 => x"79",
          9862 => x"56",
          9863 => x"24",
          9864 => x"3d",
          9865 => x"74",
          9866 => x"52",
          9867 => x"c9",
          9868 => x"e0",
          9869 => x"38",
          9870 => x"78",
          9871 => x"06",
          9872 => x"16",
          9873 => x"39",
          9874 => x"82",
          9875 => x"89",
          9876 => x"fd",
          9877 => x"54",
          9878 => x"80",
          9879 => x"ff",
          9880 => x"76",
          9881 => x"3d",
          9882 => x"3d",
          9883 => x"e3",
          9884 => x"53",
          9885 => x"53",
          9886 => x"3f",
          9887 => x"51",
          9888 => x"72",
          9889 => x"3f",
          9890 => x"04",
          9891 => x"75",
          9892 => x"9a",
          9893 => x"53",
          9894 => x"80",
          9895 => x"38",
          9896 => x"ff",
          9897 => x"c3",
          9898 => x"ff",
          9899 => x"73",
          9900 => x"09",
          9901 => x"38",
          9902 => x"af",
          9903 => x"ec",
          9904 => x"71",
          9905 => x"81",
          9906 => x"ff",
          9907 => x"51",
          9908 => x"26",
          9909 => x"10",
          9910 => x"05",
          9911 => x"51",
          9912 => x"80",
          9913 => x"ff",
          9914 => x"71",
          9915 => x"0c",
          9916 => x"04",
          9917 => x"02",
          9918 => x"02",
          9919 => x"05",
          9920 => x"80",
          9921 => x"ff",
          9922 => x"70",
          9923 => x"71",
          9924 => x"09",
          9925 => x"38",
          9926 => x"26",
          9927 => x"10",
          9928 => x"05",
          9929 => x"51",
          9930 => x"98",
          9931 => x"0d",
          9932 => x"0d",
          9933 => x"83",
          9934 => x"81",
          9935 => x"83",
          9936 => x"82",
          9937 => x"52",
          9938 => x"27",
          9939 => x"d9",
          9940 => x"70",
          9941 => x"22",
          9942 => x"80",
          9943 => x"26",
          9944 => x"55",
          9945 => x"38",
          9946 => x"05",
          9947 => x"88",
          9948 => x"ff",
          9949 => x"54",
          9950 => x"71",
          9951 => x"d7",
          9952 => x"26",
          9953 => x"73",
          9954 => x"b9",
          9955 => x"70",
          9956 => x"75",
          9957 => x"11",
          9958 => x"51",
          9959 => x"39",
          9960 => x"81",
          9961 => x"31",
          9962 => x"39",
          9963 => x"9f",
          9964 => x"51",
          9965 => x"12",
          9966 => x"e6",
          9967 => x"39",
          9968 => x"8b",
          9969 => x"12",
          9970 => x"c7",
          9971 => x"70",
          9972 => x"06",
          9973 => x"73",
          9974 => x"72",
          9975 => x"fe",
          9976 => x"51",
          9977 => x"98",
          9978 => x"0d",
          9979 => x"ff",
          9980 => x"ff",
          9981 => x"00",
          9982 => x"ff",
          9983 => x"31",
          9984 => x"30",
          9985 => x"30",
          9986 => x"30",
          9987 => x"30",
          9988 => x"30",
          9989 => x"30",
          9990 => x"30",
          9991 => x"30",
          9992 => x"30",
          9993 => x"30",
          9994 => x"30",
          9995 => x"30",
          9996 => x"30",
          9997 => x"30",
          9998 => x"30",
          9999 => x"30",
         10000 => x"30",
         10001 => x"30",
         10002 => x"30",
         10003 => x"47",
         10004 => x"47",
         10005 => x"47",
         10006 => x"47",
         10007 => x"47",
         10008 => x"4d",
         10009 => x"4e",
         10010 => x"4f",
         10011 => x"51",
         10012 => x"4e",
         10013 => x"4c",
         10014 => x"50",
         10015 => x"51",
         10016 => x"50",
         10017 => x"51",
         10018 => x"50",
         10019 => x"4f",
         10020 => x"4c",
         10021 => x"4f",
         10022 => x"4f",
         10023 => x"50",
         10024 => x"4c",
         10025 => x"4c",
         10026 => x"50",
         10027 => x"51",
         10028 => x"51",
         10029 => x"51",
         10030 => x"9b",
         10031 => x"9b",
         10032 => x"9b",
         10033 => x"9b",
         10034 => x"9b",
         10035 => x"9b",
         10036 => x"9b",
         10037 => x"9b",
         10038 => x"9b",
         10039 => x"0e",
         10040 => x"17",
         10041 => x"17",
         10042 => x"0e",
         10043 => x"17",
         10044 => x"17",
         10045 => x"17",
         10046 => x"17",
         10047 => x"17",
         10048 => x"17",
         10049 => x"17",
         10050 => x"0e",
         10051 => x"17",
         10052 => x"0e",
         10053 => x"0e",
         10054 => x"17",
         10055 => x"17",
         10056 => x"17",
         10057 => x"17",
         10058 => x"17",
         10059 => x"17",
         10060 => x"17",
         10061 => x"17",
         10062 => x"17",
         10063 => x"17",
         10064 => x"17",
         10065 => x"17",
         10066 => x"17",
         10067 => x"17",
         10068 => x"17",
         10069 => x"17",
         10070 => x"17",
         10071 => x"17",
         10072 => x"17",
         10073 => x"17",
         10074 => x"17",
         10075 => x"17",
         10076 => x"17",
         10077 => x"17",
         10078 => x"17",
         10079 => x"17",
         10080 => x"17",
         10081 => x"17",
         10082 => x"17",
         10083 => x"17",
         10084 => x"17",
         10085 => x"17",
         10086 => x"17",
         10087 => x"17",
         10088 => x"17",
         10089 => x"17",
         10090 => x"0f",
         10091 => x"17",
         10092 => x"17",
         10093 => x"17",
         10094 => x"17",
         10095 => x"11",
         10096 => x"17",
         10097 => x"17",
         10098 => x"17",
         10099 => x"17",
         10100 => x"17",
         10101 => x"17",
         10102 => x"17",
         10103 => x"17",
         10104 => x"17",
         10105 => x"17",
         10106 => x"0f",
         10107 => x"10",
         10108 => x"0e",
         10109 => x"0e",
         10110 => x"0e",
         10111 => x"17",
         10112 => x"10",
         10113 => x"17",
         10114 => x"17",
         10115 => x"0e",
         10116 => x"17",
         10117 => x"17",
         10118 => x"11",
         10119 => x"11",
         10120 => x"17",
         10121 => x"17",
         10122 => x"0f",
         10123 => x"17",
         10124 => x"11",
         10125 => x"17",
         10126 => x"17",
         10127 => x"11",
         10128 => x"6e",
         10129 => x"00",
         10130 => x"6f",
         10131 => x"00",
         10132 => x"6e",
         10133 => x"00",
         10134 => x"6f",
         10135 => x"00",
         10136 => x"78",
         10137 => x"00",
         10138 => x"6c",
         10139 => x"00",
         10140 => x"6f",
         10141 => x"00",
         10142 => x"69",
         10143 => x"00",
         10144 => x"75",
         10145 => x"00",
         10146 => x"62",
         10147 => x"68",
         10148 => x"77",
         10149 => x"64",
         10150 => x"65",
         10151 => x"64",
         10152 => x"65",
         10153 => x"6c",
         10154 => x"00",
         10155 => x"70",
         10156 => x"73",
         10157 => x"74",
         10158 => x"73",
         10159 => x"00",
         10160 => x"66",
         10161 => x"00",
         10162 => x"61",
         10163 => x"00",
         10164 => x"61",
         10165 => x"00",
         10166 => x"6c",
         10167 => x"00",
         10168 => x"00",
         10169 => x"73",
         10170 => x"72",
         10171 => x"00",
         10172 => x"74",
         10173 => x"61",
         10174 => x"72",
         10175 => x"2e",
         10176 => x"73",
         10177 => x"6f",
         10178 => x"65",
         10179 => x"2e",
         10180 => x"20",
         10181 => x"65",
         10182 => x"75",
         10183 => x"00",
         10184 => x"20",
         10185 => x"68",
         10186 => x"75",
         10187 => x"00",
         10188 => x"76",
         10189 => x"64",
         10190 => x"6c",
         10191 => x"6d",
         10192 => x"00",
         10193 => x"63",
         10194 => x"20",
         10195 => x"69",
         10196 => x"00",
         10197 => x"6c",
         10198 => x"6c",
         10199 => x"64",
         10200 => x"78",
         10201 => x"73",
         10202 => x"00",
         10203 => x"6c",
         10204 => x"61",
         10205 => x"65",
         10206 => x"76",
         10207 => x"64",
         10208 => x"00",
         10209 => x"20",
         10210 => x"77",
         10211 => x"65",
         10212 => x"6f",
         10213 => x"74",
         10214 => x"00",
         10215 => x"69",
         10216 => x"6e",
         10217 => x"65",
         10218 => x"73",
         10219 => x"76",
         10220 => x"64",
         10221 => x"00",
         10222 => x"73",
         10223 => x"6f",
         10224 => x"6e",
         10225 => x"65",
         10226 => x"00",
         10227 => x"20",
         10228 => x"70",
         10229 => x"62",
         10230 => x"66",
         10231 => x"73",
         10232 => x"65",
         10233 => x"6f",
         10234 => x"20",
         10235 => x"64",
         10236 => x"2e",
         10237 => x"72",
         10238 => x"20",
         10239 => x"72",
         10240 => x"2e",
         10241 => x"6d",
         10242 => x"74",
         10243 => x"70",
         10244 => x"74",
         10245 => x"20",
         10246 => x"63",
         10247 => x"65",
         10248 => x"00",
         10249 => x"6c",
         10250 => x"73",
         10251 => x"63",
         10252 => x"2e",
         10253 => x"73",
         10254 => x"69",
         10255 => x"6e",
         10256 => x"65",
         10257 => x"79",
         10258 => x"00",
         10259 => x"6f",
         10260 => x"6e",
         10261 => x"70",
         10262 => x"66",
         10263 => x"73",
         10264 => x"00",
         10265 => x"72",
         10266 => x"74",
         10267 => x"20",
         10268 => x"6f",
         10269 => x"63",
         10270 => x"00",
         10271 => x"63",
         10272 => x"73",
         10273 => x"00",
         10274 => x"6b",
         10275 => x"6e",
         10276 => x"72",
         10277 => x"00",
         10278 => x"6c",
         10279 => x"79",
         10280 => x"20",
         10281 => x"61",
         10282 => x"6c",
         10283 => x"79",
         10284 => x"2f",
         10285 => x"2e",
         10286 => x"00",
         10287 => x"61",
         10288 => x"00",
         10289 => x"38",
         10290 => x"00",
         10291 => x"20",
         10292 => x"34",
         10293 => x"00",
         10294 => x"20",
         10295 => x"20",
         10296 => x"00",
         10297 => x"32",
         10298 => x"00",
         10299 => x"00",
         10300 => x"00",
         10301 => x"00",
         10302 => x"53",
         10303 => x"20",
         10304 => x"28",
         10305 => x"2f",
         10306 => x"32",
         10307 => x"00",
         10308 => x"2e",
         10309 => x"00",
         10310 => x"50",
         10311 => x"72",
         10312 => x"25",
         10313 => x"29",
         10314 => x"20",
         10315 => x"2a",
         10316 => x"00",
         10317 => x"55",
         10318 => x"74",
         10319 => x"75",
         10320 => x"48",
         10321 => x"6c",
         10322 => x"00",
         10323 => x"6d",
         10324 => x"69",
         10325 => x"72",
         10326 => x"74",
         10327 => x"32",
         10328 => x"74",
         10329 => x"75",
         10330 => x"00",
         10331 => x"43",
         10332 => x"52",
         10333 => x"6e",
         10334 => x"72",
         10335 => x"00",
         10336 => x"43",
         10337 => x"57",
         10338 => x"6e",
         10339 => x"72",
         10340 => x"00",
         10341 => x"52",
         10342 => x"52",
         10343 => x"6e",
         10344 => x"72",
         10345 => x"00",
         10346 => x"52",
         10347 => x"54",
         10348 => x"6e",
         10349 => x"72",
         10350 => x"00",
         10351 => x"52",
         10352 => x"52",
         10353 => x"6e",
         10354 => x"72",
         10355 => x"00",
         10356 => x"52",
         10357 => x"54",
         10358 => x"6e",
         10359 => x"72",
         10360 => x"00",
         10361 => x"74",
         10362 => x"67",
         10363 => x"20",
         10364 => x"65",
         10365 => x"2e",
         10366 => x"61",
         10367 => x"6e",
         10368 => x"69",
         10369 => x"2e",
         10370 => x"00",
         10371 => x"74",
         10372 => x"65",
         10373 => x"61",
         10374 => x"00",
         10375 => x"53",
         10376 => x"75",
         10377 => x"74",
         10378 => x"00",
         10379 => x"69",
         10380 => x"20",
         10381 => x"69",
         10382 => x"69",
         10383 => x"73",
         10384 => x"64",
         10385 => x"72",
         10386 => x"2c",
         10387 => x"65",
         10388 => x"20",
         10389 => x"74",
         10390 => x"6e",
         10391 => x"6c",
         10392 => x"00",
         10393 => x"00",
         10394 => x"65",
         10395 => x"6e",
         10396 => x"2e",
         10397 => x"00",
         10398 => x"70",
         10399 => x"67",
         10400 => x"00",
         10401 => x"6d",
         10402 => x"69",
         10403 => x"2e",
         10404 => x"00",
         10405 => x"38",
         10406 => x"25",
         10407 => x"29",
         10408 => x"30",
         10409 => x"28",
         10410 => x"78",
         10411 => x"00",
         10412 => x"6d",
         10413 => x"65",
         10414 => x"79",
         10415 => x"6f",
         10416 => x"65",
         10417 => x"00",
         10418 => x"38",
         10419 => x"25",
         10420 => x"2d",
         10421 => x"3f",
         10422 => x"38",
         10423 => x"25",
         10424 => x"2d",
         10425 => x"38",
         10426 => x"25",
         10427 => x"58",
         10428 => x"00",
         10429 => x"65",
         10430 => x"69",
         10431 => x"63",
         10432 => x"20",
         10433 => x"30",
         10434 => x"20",
         10435 => x"0a",
         10436 => x"6c",
         10437 => x"67",
         10438 => x"64",
         10439 => x"20",
         10440 => x"6c",
         10441 => x"2e",
         10442 => x"00",
         10443 => x"6c",
         10444 => x"65",
         10445 => x"6e",
         10446 => x"63",
         10447 => x"20",
         10448 => x"29",
         10449 => x"00",
         10450 => x"73",
         10451 => x"74",
         10452 => x"20",
         10453 => x"6c",
         10454 => x"74",
         10455 => x"2e",
         10456 => x"00",
         10457 => x"6c",
         10458 => x"65",
         10459 => x"74",
         10460 => x"2e",
         10461 => x"00",
         10462 => x"55",
         10463 => x"6e",
         10464 => x"3a",
         10465 => x"5c",
         10466 => x"25",
         10467 => x"00",
         10468 => x"3a",
         10469 => x"5c",
         10470 => x"00",
         10471 => x"3a",
         10472 => x"00",
         10473 => x"64",
         10474 => x"6d",
         10475 => x"64",
         10476 => x"00",
         10477 => x"6d",
         10478 => x"20",
         10479 => x"61",
         10480 => x"65",
         10481 => x"63",
         10482 => x"6f",
         10483 => x"72",
         10484 => x"73",
         10485 => x"6f",
         10486 => x"6e",
         10487 => x"00",
         10488 => x"6e",
         10489 => x"67",
         10490 => x"00",
         10491 => x"61",
         10492 => x"6e",
         10493 => x"6e",
         10494 => x"72",
         10495 => x"73",
         10496 => x"00",
         10497 => x"2f",
         10498 => x"25",
         10499 => x"64",
         10500 => x"3a",
         10501 => x"25",
         10502 => x"0a",
         10503 => x"43",
         10504 => x"6e",
         10505 => x"75",
         10506 => x"69",
         10507 => x"00",
         10508 => x"66",
         10509 => x"20",
         10510 => x"20",
         10511 => x"66",
         10512 => x"00",
         10513 => x"44",
         10514 => x"63",
         10515 => x"69",
         10516 => x"65",
         10517 => x"74",
         10518 => x"00",
         10519 => x"20",
         10520 => x"20",
         10521 => x"41",
         10522 => x"28",
         10523 => x"58",
         10524 => x"38",
         10525 => x"0a",
         10526 => x"20",
         10527 => x"52",
         10528 => x"20",
         10529 => x"28",
         10530 => x"58",
         10531 => x"38",
         10532 => x"0a",
         10533 => x"20",
         10534 => x"53",
         10535 => x"52",
         10536 => x"28",
         10537 => x"58",
         10538 => x"38",
         10539 => x"0a",
         10540 => x"20",
         10541 => x"41",
         10542 => x"20",
         10543 => x"28",
         10544 => x"58",
         10545 => x"38",
         10546 => x"0a",
         10547 => x"20",
         10548 => x"4d",
         10549 => x"20",
         10550 => x"28",
         10551 => x"58",
         10552 => x"38",
         10553 => x"0a",
         10554 => x"20",
         10555 => x"20",
         10556 => x"44",
         10557 => x"28",
         10558 => x"69",
         10559 => x"20",
         10560 => x"32",
         10561 => x"0a",
         10562 => x"20",
         10563 => x"4d",
         10564 => x"20",
         10565 => x"28",
         10566 => x"65",
         10567 => x"20",
         10568 => x"32",
         10569 => x"0a",
         10570 => x"20",
         10571 => x"54",
         10572 => x"54",
         10573 => x"28",
         10574 => x"6e",
         10575 => x"73",
         10576 => x"32",
         10577 => x"0a",
         10578 => x"20",
         10579 => x"53",
         10580 => x"4e",
         10581 => x"55",
         10582 => x"00",
         10583 => x"20",
         10584 => x"20",
         10585 => x"00",
         10586 => x"20",
         10587 => x"43",
         10588 => x"00",
         10589 => x"20",
         10590 => x"32",
         10591 => x"20",
         10592 => x"49",
         10593 => x"64",
         10594 => x"73",
         10595 => x"00",
         10596 => x"20",
         10597 => x"55",
         10598 => x"73",
         10599 => x"56",
         10600 => x"6f",
         10601 => x"64",
         10602 => x"73",
         10603 => x"20",
         10604 => x"58",
         10605 => x"00",
         10606 => x"20",
         10607 => x"55",
         10608 => x"6d",
         10609 => x"20",
         10610 => x"72",
         10611 => x"64",
         10612 => x"73",
         10613 => x"20",
         10614 => x"58",
         10615 => x"00",
         10616 => x"20",
         10617 => x"61",
         10618 => x"53",
         10619 => x"74",
         10620 => x"64",
         10621 => x"73",
         10622 => x"20",
         10623 => x"20",
         10624 => x"58",
         10625 => x"00",
         10626 => x"73",
         10627 => x"00",
         10628 => x"20",
         10629 => x"55",
         10630 => x"20",
         10631 => x"20",
         10632 => x"20",
         10633 => x"20",
         10634 => x"20",
         10635 => x"20",
         10636 => x"58",
         10637 => x"00",
         10638 => x"20",
         10639 => x"73",
         10640 => x"20",
         10641 => x"63",
         10642 => x"72",
         10643 => x"20",
         10644 => x"20",
         10645 => x"20",
         10646 => x"25",
         10647 => x"4d",
         10648 => x"00",
         10649 => x"20",
         10650 => x"52",
         10651 => x"43",
         10652 => x"6b",
         10653 => x"65",
         10654 => x"20",
         10655 => x"20",
         10656 => x"20",
         10657 => x"25",
         10658 => x"4d",
         10659 => x"00",
         10660 => x"20",
         10661 => x"73",
         10662 => x"6e",
         10663 => x"44",
         10664 => x"20",
         10665 => x"63",
         10666 => x"72",
         10667 => x"20",
         10668 => x"25",
         10669 => x"4d",
         10670 => x"00",
         10671 => x"61",
         10672 => x"00",
         10673 => x"64",
         10674 => x"00",
         10675 => x"65",
         10676 => x"00",
         10677 => x"4f",
         10678 => x"4f",
         10679 => x"00",
         10680 => x"6b",
         10681 => x"6e",
         10682 => x"a8",
         10683 => x"00",
         10684 => x"00",
         10685 => x"a8",
         10686 => x"00",
         10687 => x"00",
         10688 => x"a8",
         10689 => x"00",
         10690 => x"00",
         10691 => x"a8",
         10692 => x"00",
         10693 => x"00",
         10694 => x"a8",
         10695 => x"00",
         10696 => x"00",
         10697 => x"a8",
         10698 => x"00",
         10699 => x"00",
         10700 => x"a8",
         10701 => x"00",
         10702 => x"00",
         10703 => x"a8",
         10704 => x"00",
         10705 => x"00",
         10706 => x"a8",
         10707 => x"00",
         10708 => x"00",
         10709 => x"a8",
         10710 => x"00",
         10711 => x"00",
         10712 => x"a8",
         10713 => x"00",
         10714 => x"00",
         10715 => x"a8",
         10716 => x"00",
         10717 => x"00",
         10718 => x"a8",
         10719 => x"00",
         10720 => x"00",
         10721 => x"a8",
         10722 => x"00",
         10723 => x"00",
         10724 => x"a8",
         10725 => x"00",
         10726 => x"00",
         10727 => x"a8",
         10728 => x"00",
         10729 => x"00",
         10730 => x"a8",
         10731 => x"00",
         10732 => x"00",
         10733 => x"a8",
         10734 => x"00",
         10735 => x"00",
         10736 => x"a7",
         10737 => x"00",
         10738 => x"00",
         10739 => x"a7",
         10740 => x"00",
         10741 => x"00",
         10742 => x"a7",
         10743 => x"00",
         10744 => x"00",
         10745 => x"a7",
         10746 => x"00",
         10747 => x"00",
         10748 => x"44",
         10749 => x"43",
         10750 => x"42",
         10751 => x"41",
         10752 => x"36",
         10753 => x"35",
         10754 => x"34",
         10755 => x"46",
         10756 => x"33",
         10757 => x"32",
         10758 => x"31",
         10759 => x"00",
         10760 => x"00",
         10761 => x"00",
         10762 => x"00",
         10763 => x"00",
         10764 => x"00",
         10765 => x"00",
         10766 => x"00",
         10767 => x"00",
         10768 => x"00",
         10769 => x"00",
         10770 => x"73",
         10771 => x"79",
         10772 => x"73",
         10773 => x"00",
         10774 => x"00",
         10775 => x"34",
         10776 => x"20",
         10777 => x"00",
         10778 => x"69",
         10779 => x"20",
         10780 => x"72",
         10781 => x"74",
         10782 => x"65",
         10783 => x"73",
         10784 => x"79",
         10785 => x"6c",
         10786 => x"6f",
         10787 => x"46",
         10788 => x"00",
         10789 => x"6e",
         10790 => x"20",
         10791 => x"6e",
         10792 => x"65",
         10793 => x"20",
         10794 => x"74",
         10795 => x"20",
         10796 => x"65",
         10797 => x"69",
         10798 => x"6c",
         10799 => x"2e",
         10800 => x"00",
         10801 => x"3a",
         10802 => x"7c",
         10803 => x"00",
         10804 => x"3b",
         10805 => x"00",
         10806 => x"54",
         10807 => x"54",
         10808 => x"00",
         10809 => x"90",
         10810 => x"4f",
         10811 => x"30",
         10812 => x"20",
         10813 => x"45",
         10814 => x"20",
         10815 => x"33",
         10816 => x"20",
         10817 => x"20",
         10818 => x"45",
         10819 => x"20",
         10820 => x"20",
         10821 => x"20",
         10822 => x"a8",
         10823 => x"00",
         10824 => x"00",
         10825 => x"00",
         10826 => x"05",
         10827 => x"10",
         10828 => x"18",
         10829 => x"00",
         10830 => x"45",
         10831 => x"8f",
         10832 => x"45",
         10833 => x"8e",
         10834 => x"92",
         10835 => x"55",
         10836 => x"9a",
         10837 => x"9e",
         10838 => x"4f",
         10839 => x"a6",
         10840 => x"aa",
         10841 => x"ae",
         10842 => x"b2",
         10843 => x"b6",
         10844 => x"ba",
         10845 => x"be",
         10846 => x"c2",
         10847 => x"c6",
         10848 => x"ca",
         10849 => x"ce",
         10850 => x"d2",
         10851 => x"d6",
         10852 => x"da",
         10853 => x"de",
         10854 => x"e2",
         10855 => x"e6",
         10856 => x"ea",
         10857 => x"ee",
         10858 => x"f2",
         10859 => x"f6",
         10860 => x"fa",
         10861 => x"fe",
         10862 => x"2c",
         10863 => x"5d",
         10864 => x"2a",
         10865 => x"3f",
         10866 => x"00",
         10867 => x"00",
         10868 => x"00",
         10869 => x"02",
         10870 => x"00",
         10871 => x"00",
         10872 => x"00",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"01",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"23",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"25",
         10900 => x"25",
         10901 => x"25",
         10902 => x"25",
         10903 => x"25",
         10904 => x"25",
         10905 => x"25",
         10906 => x"25",
         10907 => x"25",
         10908 => x"25",
         10909 => x"25",
         10910 => x"25",
         10911 => x"25",
         10912 => x"25",
         10913 => x"25",
         10914 => x"25",
         10915 => x"25",
         10916 => x"25",
         10917 => x"25",
         10918 => x"25",
         10919 => x"25",
         10920 => x"25",
         10921 => x"25",
         10922 => x"25",
         10923 => x"00",
         10924 => x"03",
         10925 => x"03",
         10926 => x"03",
         10927 => x"03",
         10928 => x"03",
         10929 => x"03",
         10930 => x"22",
         10931 => x"00",
         10932 => x"22",
         10933 => x"23",
         10934 => x"22",
         10935 => x"22",
         10936 => x"22",
         10937 => x"00",
         10938 => x"00",
         10939 => x"03",
         10940 => x"03",
         10941 => x"03",
         10942 => x"00",
         10943 => x"01",
         10944 => x"01",
         10945 => x"01",
         10946 => x"01",
         10947 => x"01",
         10948 => x"01",
         10949 => x"02",
         10950 => x"01",
         10951 => x"01",
         10952 => x"01",
         10953 => x"01",
         10954 => x"01",
         10955 => x"01",
         10956 => x"01",
         10957 => x"01",
         10958 => x"01",
         10959 => x"01",
         10960 => x"01",
         10961 => x"01",
         10962 => x"02",
         10963 => x"01",
         10964 => x"02",
         10965 => x"01",
         10966 => x"01",
         10967 => x"01",
         10968 => x"01",
         10969 => x"01",
         10970 => x"01",
         10971 => x"01",
         10972 => x"01",
         10973 => x"01",
         10974 => x"01",
         10975 => x"01",
         10976 => x"01",
         10977 => x"01",
         10978 => x"01",
         10979 => x"01",
         10980 => x"01",
         10981 => x"01",
         10982 => x"01",
         10983 => x"01",
         10984 => x"01",
         10985 => x"01",
         10986 => x"01",
         10987 => x"01",
         10988 => x"01",
         10989 => x"00",
         10990 => x"01",
         10991 => x"01",
         10992 => x"01",
         10993 => x"01",
         10994 => x"01",
         10995 => x"01",
         10996 => x"00",
         10997 => x"02",
         10998 => x"02",
         10999 => x"02",
         11000 => x"02",
         11001 => x"02",
         11002 => x"02",
         11003 => x"01",
         11004 => x"02",
         11005 => x"01",
         11006 => x"01",
         11007 => x"01",
         11008 => x"02",
         11009 => x"02",
         11010 => x"02",
         11011 => x"01",
         11012 => x"02",
         11013 => x"02",
         11014 => x"01",
         11015 => x"2c",
         11016 => x"02",
         11017 => x"01",
         11018 => x"02",
         11019 => x"02",
         11020 => x"01",
         11021 => x"02",
         11022 => x"02",
         11023 => x"02",
         11024 => x"2c",
         11025 => x"02",
         11026 => x"02",
         11027 => x"01",
         11028 => x"02",
         11029 => x"02",
         11030 => x"02",
         11031 => x"01",
         11032 => x"02",
         11033 => x"02",
         11034 => x"02",
         11035 => x"03",
         11036 => x"03",
         11037 => x"03",
         11038 => x"00",
         11039 => x"03",
         11040 => x"03",
         11041 => x"03",
         11042 => x"00",
         11043 => x"03",
         11044 => x"03",
         11045 => x"00",
         11046 => x"03",
         11047 => x"03",
         11048 => x"03",
         11049 => x"03",
         11050 => x"03",
         11051 => x"03",
         11052 => x"03",
         11053 => x"03",
         11054 => x"04",
         11055 => x"04",
         11056 => x"04",
         11057 => x"04",
         11058 => x"04",
         11059 => x"04",
         11060 => x"04",
         11061 => x"01",
         11062 => x"04",
         11063 => x"00",
         11064 => x"00",
         11065 => x"1e",
         11066 => x"1e",
         11067 => x"1f",
         11068 => x"1f",
         11069 => x"1f",
         11070 => x"1f",
         11071 => x"1f",
         11072 => x"1f",
         11073 => x"1f",
         11074 => x"1f",
         11075 => x"1f",
         11076 => x"1f",
         11077 => x"06",
         11078 => x"00",
         11079 => x"1f",
         11080 => x"1f",
         11081 => x"1f",
         11082 => x"1f",
         11083 => x"1f",
         11084 => x"1f",
         11085 => x"1f",
         11086 => x"06",
         11087 => x"06",
         11088 => x"06",
         11089 => x"00",
         11090 => x"1f",
         11091 => x"1f",
         11092 => x"00",
         11093 => x"1f",
         11094 => x"1f",
         11095 => x"1f",
         11096 => x"1f",
         11097 => x"00",
         11098 => x"21",
         11099 => x"21",
         11100 => x"02",
         11101 => x"00",
         11102 => x"24",
         11103 => x"2c",
         11104 => x"2c",
         11105 => x"2c",
         11106 => x"2c",
         11107 => x"2c",
         11108 => x"2d",
         11109 => x"ff",
         11110 => x"00",
         11111 => x"00",
         11112 => x"9e",
         11113 => x"01",
         11114 => x"00",
         11115 => x"00",
         11116 => x"9e",
         11117 => x"01",
         11118 => x"00",
         11119 => x"00",
         11120 => x"9e",
         11121 => x"03",
         11122 => x"00",
         11123 => x"00",
         11124 => x"9e",
         11125 => x"03",
         11126 => x"00",
         11127 => x"00",
         11128 => x"9e",
         11129 => x"03",
         11130 => x"00",
         11131 => x"00",
         11132 => x"9e",
         11133 => x"04",
         11134 => x"00",
         11135 => x"00",
         11136 => x"9e",
         11137 => x"04",
         11138 => x"00",
         11139 => x"00",
         11140 => x"9e",
         11141 => x"04",
         11142 => x"00",
         11143 => x"00",
         11144 => x"9e",
         11145 => x"04",
         11146 => x"00",
         11147 => x"00",
         11148 => x"9e",
         11149 => x"04",
         11150 => x"00",
         11151 => x"00",
         11152 => x"9e",
         11153 => x"04",
         11154 => x"00",
         11155 => x"00",
         11156 => x"9e",
         11157 => x"04",
         11158 => x"00",
         11159 => x"00",
         11160 => x"9e",
         11161 => x"05",
         11162 => x"00",
         11163 => x"00",
         11164 => x"9e",
         11165 => x"05",
         11166 => x"00",
         11167 => x"00",
         11168 => x"9e",
         11169 => x"05",
         11170 => x"00",
         11171 => x"00",
         11172 => x"9e",
         11173 => x"05",
         11174 => x"00",
         11175 => x"00",
         11176 => x"9e",
         11177 => x"07",
         11178 => x"00",
         11179 => x"00",
         11180 => x"9e",
         11181 => x"07",
         11182 => x"00",
         11183 => x"00",
         11184 => x"9e",
         11185 => x"08",
         11186 => x"00",
         11187 => x"00",
         11188 => x"9e",
         11189 => x"08",
         11190 => x"00",
         11191 => x"00",
         11192 => x"9e",
         11193 => x"08",
         11194 => x"00",
         11195 => x"00",
         11196 => x"9e",
         11197 => x"09",
         11198 => x"00",
         11199 => x"00",
         11200 => x"9e",
         11201 => x"09",
         11202 => x"00",
         11203 => x"00",
         11204 => x"9e",
         11205 => x"09",
         11206 => x"00",
         11207 => x"00",
         11208 => x"9e",
         11209 => x"09",
         11210 => x"00",
         11211 => x"00",
         11212 => x"00",
         11213 => x"00",
         11214 => x"7f",
         11215 => x"00",
         11216 => x"7f",
         11217 => x"00",
         11218 => x"7f",
         11219 => x"00",
         11220 => x"00",
         11221 => x"00",
         11222 => x"ff",
         11223 => x"00",
         11224 => x"00",
         11225 => x"78",
         11226 => x"00",
         11227 => x"e1",
         11228 => x"e1",
         11229 => x"e1",
         11230 => x"00",
         11231 => x"01",
         11232 => x"01",
         11233 => x"10",
         11234 => x"00",
         11235 => x"00",
         11236 => x"00",
         11237 => x"00",
         11238 => x"00",
         11239 => x"00",
         11240 => x"00",
         11241 => x"00",
         11242 => x"00",
         11243 => x"00",
         11244 => x"00",
         11245 => x"00",
         11246 => x"00",
         11247 => x"00",
         11248 => x"00",
         11249 => x"00",
         11250 => x"00",
         11251 => x"00",
         11252 => x"00",
         11253 => x"00",
         11254 => x"00",
         11255 => x"00",
         11256 => x"00",
         11257 => x"00",
         11258 => x"00",
         11259 => x"a8",
         11260 => x"00",
         11261 => x"a8",
         11262 => x"00",
         11263 => x"a8",
         11264 => x"00",
         11265 => x"00",
         11266 => x"00",
         11267 => x"00",
         11268 => x"00",
         11269 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0d",
             2 => x"93",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"2d",
            11 => x"0c",
            12 => x"00",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"b9",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"04",
           266 => x"8c",
           267 => x"0b",
           268 => x"04",
           269 => x"8c",
           270 => x"0b",
           271 => x"04",
           272 => x"8c",
           273 => x"0b",
           274 => x"04",
           275 => x"8c",
           276 => x"0b",
           277 => x"04",
           278 => x"8d",
           279 => x"0b",
           280 => x"04",
           281 => x"8d",
           282 => x"0b",
           283 => x"04",
           284 => x"8d",
           285 => x"0b",
           286 => x"04",
           287 => x"8d",
           288 => x"0b",
           289 => x"04",
           290 => x"8e",
           291 => x"0b",
           292 => x"04",
           293 => x"8e",
           294 => x"0b",
           295 => x"04",
           296 => x"8e",
           297 => x"0b",
           298 => x"04",
           299 => x"8e",
           300 => x"0b",
           301 => x"04",
           302 => x"8f",
           303 => x"0b",
           304 => x"04",
           305 => x"8f",
           306 => x"0b",
           307 => x"04",
           308 => x"8f",
           309 => x"0b",
           310 => x"04",
           311 => x"8f",
           312 => x"0b",
           313 => x"04",
           314 => x"90",
           315 => x"0b",
           316 => x"04",
           317 => x"90",
           318 => x"0b",
           319 => x"04",
           320 => x"90",
           321 => x"0b",
           322 => x"04",
           323 => x"91",
           324 => x"0b",
           325 => x"04",
           326 => x"91",
           327 => x"0b",
           328 => x"04",
           329 => x"91",
           330 => x"0b",
           331 => x"04",
           332 => x"91",
           333 => x"0b",
           334 => x"04",
           335 => x"92",
           336 => x"0b",
           337 => x"04",
           338 => x"92",
           339 => x"0b",
           340 => x"04",
           341 => x"92",
           342 => x"0b",
           343 => x"04",
           344 => x"92",
           345 => x"0b",
           346 => x"04",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"00",
           385 => x"82",
           386 => x"81",
           387 => x"82",
           388 => x"80",
           389 => x"04",
           390 => x"0c",
           391 => x"82",
           392 => x"80",
           393 => x"04",
           394 => x"0c",
           395 => x"82",
           396 => x"80",
           397 => x"04",
           398 => x"0c",
           399 => x"82",
           400 => x"80",
           401 => x"04",
           402 => x"0c",
           403 => x"82",
           404 => x"80",
           405 => x"04",
           406 => x"0c",
           407 => x"82",
           408 => x"80",
           409 => x"04",
           410 => x"0c",
           411 => x"2d",
           412 => x"08",
           413 => x"90",
           414 => x"a4",
           415 => x"ce",
           416 => x"a4",
           417 => x"80",
           418 => x"e0",
           419 => x"8c",
           420 => x"a4",
           421 => x"80",
           422 => x"e0",
           423 => x"f4",
           424 => x"a4",
           425 => x"80",
           426 => x"e0",
           427 => x"81",
           428 => x"a4",
           429 => x"80",
           430 => x"e0",
           431 => x"e0",
           432 => x"e0",
           433 => x"c0",
           434 => x"82",
           435 => x"80",
           436 => x"82",
           437 => x"80",
           438 => x"04",
           439 => x"0c",
           440 => x"2d",
           441 => x"08",
           442 => x"90",
           443 => x"a4",
           444 => x"b2",
           445 => x"a4",
           446 => x"80",
           447 => x"e0",
           448 => x"fe",
           449 => x"e0",
           450 => x"c0",
           451 => x"82",
           452 => x"81",
           453 => x"82",
           454 => x"80",
           455 => x"04",
           456 => x"0c",
           457 => x"2d",
           458 => x"08",
           459 => x"90",
           460 => x"a4",
           461 => x"8c",
           462 => x"a4",
           463 => x"80",
           464 => x"e0",
           465 => x"fe",
           466 => x"e0",
           467 => x"c0",
           468 => x"82",
           469 => x"82",
           470 => x"82",
           471 => x"80",
           472 => x"04",
           473 => x"0c",
           474 => x"2d",
           475 => x"08",
           476 => x"90",
           477 => x"a4",
           478 => x"84",
           479 => x"a4",
           480 => x"80",
           481 => x"e0",
           482 => x"8c",
           483 => x"e0",
           484 => x"c0",
           485 => x"82",
           486 => x"82",
           487 => x"82",
           488 => x"80",
           489 => x"04",
           490 => x"0c",
           491 => x"2d",
           492 => x"08",
           493 => x"90",
           494 => x"a4",
           495 => x"bb",
           496 => x"a4",
           497 => x"80",
           498 => x"e0",
           499 => x"93",
           500 => x"e0",
           501 => x"c0",
           502 => x"82",
           503 => x"82",
           504 => x"82",
           505 => x"80",
           506 => x"04",
           507 => x"0c",
           508 => x"2d",
           509 => x"08",
           510 => x"90",
           511 => x"a4",
           512 => x"9c",
           513 => x"a4",
           514 => x"80",
           515 => x"e0",
           516 => x"9c",
           517 => x"e0",
           518 => x"c0",
           519 => x"82",
           520 => x"82",
           521 => x"82",
           522 => x"80",
           523 => x"04",
           524 => x"0c",
           525 => x"2d",
           526 => x"08",
           527 => x"90",
           528 => x"a4",
           529 => x"8b",
           530 => x"a4",
           531 => x"80",
           532 => x"e0",
           533 => x"8f",
           534 => x"e0",
           535 => x"c0",
           536 => x"82",
           537 => x"82",
           538 => x"82",
           539 => x"80",
           540 => x"04",
           541 => x"0c",
           542 => x"2d",
           543 => x"08",
           544 => x"90",
           545 => x"a4",
           546 => x"a0",
           547 => x"a4",
           548 => x"80",
           549 => x"e0",
           550 => x"f5",
           551 => x"e0",
           552 => x"c0",
           553 => x"82",
           554 => x"82",
           555 => x"82",
           556 => x"80",
           557 => x"04",
           558 => x"0c",
           559 => x"2d",
           560 => x"08",
           561 => x"90",
           562 => x"a4",
           563 => x"d5",
           564 => x"a4",
           565 => x"80",
           566 => x"e0",
           567 => x"b5",
           568 => x"e0",
           569 => x"c0",
           570 => x"82",
           571 => x"81",
           572 => x"82",
           573 => x"80",
           574 => x"04",
           575 => x"0c",
           576 => x"2d",
           577 => x"08",
           578 => x"90",
           579 => x"a4",
           580 => x"e4",
           581 => x"a4",
           582 => x"80",
           583 => x"e0",
           584 => x"fd",
           585 => x"e0",
           586 => x"c0",
           587 => x"82",
           588 => x"81",
           589 => x"82",
           590 => x"80",
           591 => x"04",
           592 => x"0c",
           593 => x"2d",
           594 => x"08",
           595 => x"90",
           596 => x"a4",
           597 => x"9f",
           598 => x"a4",
           599 => x"80",
           600 => x"e0",
           601 => x"af",
           602 => x"e0",
           603 => x"c0",
           604 => x"82",
           605 => x"81",
           606 => x"82",
           607 => x"80",
           608 => x"04",
           609 => x"0c",
           610 => x"2d",
           611 => x"08",
           612 => x"90",
           613 => x"10",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"10",
           621 => x"51",
           622 => x"73",
           623 => x"73",
           624 => x"81",
           625 => x"10",
           626 => x"07",
           627 => x"0c",
           628 => x"72",
           629 => x"81",
           630 => x"09",
           631 => x"71",
           632 => x"0a",
           633 => x"72",
           634 => x"51",
           635 => x"82",
           636 => x"82",
           637 => x"8e",
           638 => x"70",
           639 => x"0c",
           640 => x"93",
           641 => x"81",
           642 => x"a7",
           643 => x"e0",
           644 => x"82",
           645 => x"fb",
           646 => x"e0",
           647 => x"05",
           648 => x"a4",
           649 => x"0c",
           650 => x"08",
           651 => x"54",
           652 => x"08",
           653 => x"53",
           654 => x"08",
           655 => x"9a",
           656 => x"98",
           657 => x"e0",
           658 => x"05",
           659 => x"a4",
           660 => x"08",
           661 => x"98",
           662 => x"87",
           663 => x"e0",
           664 => x"82",
           665 => x"02",
           666 => x"0c",
           667 => x"82",
           668 => x"90",
           669 => x"11",
           670 => x"32",
           671 => x"51",
           672 => x"71",
           673 => x"0b",
           674 => x"08",
           675 => x"25",
           676 => x"39",
           677 => x"e0",
           678 => x"05",
           679 => x"39",
           680 => x"08",
           681 => x"ff",
           682 => x"a4",
           683 => x"0c",
           684 => x"e0",
           685 => x"05",
           686 => x"a4",
           687 => x"08",
           688 => x"08",
           689 => x"82",
           690 => x"f8",
           691 => x"2e",
           692 => x"80",
           693 => x"a4",
           694 => x"08",
           695 => x"38",
           696 => x"08",
           697 => x"51",
           698 => x"82",
           699 => x"70",
           700 => x"08",
           701 => x"52",
           702 => x"08",
           703 => x"ff",
           704 => x"06",
           705 => x"0b",
           706 => x"08",
           707 => x"80",
           708 => x"e0",
           709 => x"05",
           710 => x"a4",
           711 => x"08",
           712 => x"73",
           713 => x"a4",
           714 => x"08",
           715 => x"e0",
           716 => x"05",
           717 => x"a4",
           718 => x"08",
           719 => x"e0",
           720 => x"05",
           721 => x"39",
           722 => x"08",
           723 => x"52",
           724 => x"82",
           725 => x"88",
           726 => x"82",
           727 => x"f4",
           728 => x"82",
           729 => x"f4",
           730 => x"e0",
           731 => x"3d",
           732 => x"a4",
           733 => x"e0",
           734 => x"82",
           735 => x"f4",
           736 => x"0b",
           737 => x"08",
           738 => x"82",
           739 => x"88",
           740 => x"e0",
           741 => x"05",
           742 => x"0b",
           743 => x"08",
           744 => x"82",
           745 => x"90",
           746 => x"e0",
           747 => x"05",
           748 => x"a4",
           749 => x"08",
           750 => x"a4",
           751 => x"08",
           752 => x"a4",
           753 => x"70",
           754 => x"81",
           755 => x"e0",
           756 => x"82",
           757 => x"dc",
           758 => x"e0",
           759 => x"05",
           760 => x"a4",
           761 => x"08",
           762 => x"80",
           763 => x"e0",
           764 => x"05",
           765 => x"e0",
           766 => x"8e",
           767 => x"e0",
           768 => x"82",
           769 => x"02",
           770 => x"0c",
           771 => x"82",
           772 => x"90",
           773 => x"e0",
           774 => x"05",
           775 => x"a4",
           776 => x"08",
           777 => x"a4",
           778 => x"08",
           779 => x"a4",
           780 => x"08",
           781 => x"3f",
           782 => x"08",
           783 => x"a4",
           784 => x"0c",
           785 => x"08",
           786 => x"70",
           787 => x"0c",
           788 => x"3d",
           789 => x"a4",
           790 => x"e0",
           791 => x"82",
           792 => x"ed",
           793 => x"0b",
           794 => x"08",
           795 => x"82",
           796 => x"88",
           797 => x"80",
           798 => x"0c",
           799 => x"08",
           800 => x"85",
           801 => x"81",
           802 => x"32",
           803 => x"51",
           804 => x"53",
           805 => x"8d",
           806 => x"82",
           807 => x"e0",
           808 => x"ac",
           809 => x"a4",
           810 => x"08",
           811 => x"53",
           812 => x"a4",
           813 => x"34",
           814 => x"06",
           815 => x"2e",
           816 => x"82",
           817 => x"8c",
           818 => x"05",
           819 => x"08",
           820 => x"82",
           821 => x"e4",
           822 => x"81",
           823 => x"72",
           824 => x"8b",
           825 => x"a4",
           826 => x"33",
           827 => x"27",
           828 => x"82",
           829 => x"f8",
           830 => x"72",
           831 => x"ee",
           832 => x"a4",
           833 => x"33",
           834 => x"2e",
           835 => x"80",
           836 => x"e0",
           837 => x"05",
           838 => x"2b",
           839 => x"51",
           840 => x"b2",
           841 => x"a4",
           842 => x"22",
           843 => x"70",
           844 => x"81",
           845 => x"51",
           846 => x"2e",
           847 => x"e0",
           848 => x"05",
           849 => x"80",
           850 => x"72",
           851 => x"08",
           852 => x"fe",
           853 => x"e0",
           854 => x"05",
           855 => x"2b",
           856 => x"70",
           857 => x"72",
           858 => x"51",
           859 => x"51",
           860 => x"82",
           861 => x"e8",
           862 => x"e0",
           863 => x"05",
           864 => x"e0",
           865 => x"05",
           866 => x"d0",
           867 => x"53",
           868 => x"a4",
           869 => x"34",
           870 => x"08",
           871 => x"70",
           872 => x"98",
           873 => x"53",
           874 => x"8b",
           875 => x"0b",
           876 => x"08",
           877 => x"82",
           878 => x"e4",
           879 => x"83",
           880 => x"06",
           881 => x"72",
           882 => x"82",
           883 => x"e8",
           884 => x"88",
           885 => x"2b",
           886 => x"70",
           887 => x"51",
           888 => x"72",
           889 => x"08",
           890 => x"fd",
           891 => x"e0",
           892 => x"05",
           893 => x"2a",
           894 => x"51",
           895 => x"80",
           896 => x"82",
           897 => x"e8",
           898 => x"98",
           899 => x"2c",
           900 => x"72",
           901 => x"0b",
           902 => x"08",
           903 => x"82",
           904 => x"f8",
           905 => x"11",
           906 => x"08",
           907 => x"53",
           908 => x"08",
           909 => x"80",
           910 => x"94",
           911 => x"a4",
           912 => x"08",
           913 => x"82",
           914 => x"70",
           915 => x"51",
           916 => x"82",
           917 => x"e4",
           918 => x"90",
           919 => x"72",
           920 => x"08",
           921 => x"82",
           922 => x"e4",
           923 => x"a0",
           924 => x"72",
           925 => x"08",
           926 => x"fc",
           927 => x"e0",
           928 => x"05",
           929 => x"80",
           930 => x"72",
           931 => x"08",
           932 => x"fc",
           933 => x"e0",
           934 => x"05",
           935 => x"c0",
           936 => x"72",
           937 => x"08",
           938 => x"fb",
           939 => x"e0",
           940 => x"05",
           941 => x"07",
           942 => x"82",
           943 => x"e4",
           944 => x"0b",
           945 => x"08",
           946 => x"fb",
           947 => x"e0",
           948 => x"05",
           949 => x"07",
           950 => x"82",
           951 => x"e4",
           952 => x"c1",
           953 => x"82",
           954 => x"fc",
           955 => x"e0",
           956 => x"05",
           957 => x"51",
           958 => x"e0",
           959 => x"05",
           960 => x"0b",
           961 => x"08",
           962 => x"8d",
           963 => x"e0",
           964 => x"05",
           965 => x"a4",
           966 => x"08",
           967 => x"e0",
           968 => x"05",
           969 => x"51",
           970 => x"e0",
           971 => x"05",
           972 => x"a4",
           973 => x"22",
           974 => x"53",
           975 => x"a4",
           976 => x"23",
           977 => x"82",
           978 => x"90",
           979 => x"e0",
           980 => x"05",
           981 => x"82",
           982 => x"90",
           983 => x"08",
           984 => x"08",
           985 => x"82",
           986 => x"e4",
           987 => x"83",
           988 => x"06",
           989 => x"53",
           990 => x"ab",
           991 => x"a4",
           992 => x"33",
           993 => x"53",
           994 => x"53",
           995 => x"08",
           996 => x"52",
           997 => x"3f",
           998 => x"08",
           999 => x"e0",
          1000 => x"05",
          1001 => x"82",
          1002 => x"fc",
          1003 => x"9d",
          1004 => x"e0",
          1005 => x"72",
          1006 => x"08",
          1007 => x"82",
          1008 => x"ec",
          1009 => x"82",
          1010 => x"f4",
          1011 => x"71",
          1012 => x"72",
          1013 => x"08",
          1014 => x"8b",
          1015 => x"e0",
          1016 => x"05",
          1017 => x"a4",
          1018 => x"08",
          1019 => x"e0",
          1020 => x"05",
          1021 => x"82",
          1022 => x"fc",
          1023 => x"e0",
          1024 => x"05",
          1025 => x"2a",
          1026 => x"51",
          1027 => x"72",
          1028 => x"38",
          1029 => x"08",
          1030 => x"70",
          1031 => x"72",
          1032 => x"82",
          1033 => x"fc",
          1034 => x"53",
          1035 => x"82",
          1036 => x"53",
          1037 => x"a4",
          1038 => x"23",
          1039 => x"e0",
          1040 => x"05",
          1041 => x"f3",
          1042 => x"98",
          1043 => x"82",
          1044 => x"f4",
          1045 => x"e0",
          1046 => x"05",
          1047 => x"e0",
          1048 => x"05",
          1049 => x"31",
          1050 => x"82",
          1051 => x"ec",
          1052 => x"c1",
          1053 => x"a4",
          1054 => x"22",
          1055 => x"70",
          1056 => x"51",
          1057 => x"2e",
          1058 => x"e0",
          1059 => x"05",
          1060 => x"a4",
          1061 => x"08",
          1062 => x"e0",
          1063 => x"05",
          1064 => x"82",
          1065 => x"dc",
          1066 => x"a2",
          1067 => x"a4",
          1068 => x"08",
          1069 => x"08",
          1070 => x"84",
          1071 => x"a4",
          1072 => x"0c",
          1073 => x"e0",
          1074 => x"05",
          1075 => x"e0",
          1076 => x"05",
          1077 => x"a4",
          1078 => x"0c",
          1079 => x"08",
          1080 => x"80",
          1081 => x"82",
          1082 => x"e4",
          1083 => x"82",
          1084 => x"72",
          1085 => x"08",
          1086 => x"82",
          1087 => x"fc",
          1088 => x"82",
          1089 => x"fc",
          1090 => x"e0",
          1091 => x"05",
          1092 => x"bf",
          1093 => x"72",
          1094 => x"08",
          1095 => x"81",
          1096 => x"0b",
          1097 => x"08",
          1098 => x"a9",
          1099 => x"a4",
          1100 => x"22",
          1101 => x"07",
          1102 => x"82",
          1103 => x"e4",
          1104 => x"f8",
          1105 => x"a4",
          1106 => x"34",
          1107 => x"e0",
          1108 => x"05",
          1109 => x"a4",
          1110 => x"22",
          1111 => x"70",
          1112 => x"51",
          1113 => x"2e",
          1114 => x"e0",
          1115 => x"05",
          1116 => x"a4",
          1117 => x"08",
          1118 => x"e0",
          1119 => x"05",
          1120 => x"82",
          1121 => x"d8",
          1122 => x"a2",
          1123 => x"a4",
          1124 => x"08",
          1125 => x"08",
          1126 => x"84",
          1127 => x"a4",
          1128 => x"0c",
          1129 => x"e0",
          1130 => x"05",
          1131 => x"e0",
          1132 => x"05",
          1133 => x"a4",
          1134 => x"0c",
          1135 => x"08",
          1136 => x"70",
          1137 => x"53",
          1138 => x"a4",
          1139 => x"23",
          1140 => x"0b",
          1141 => x"08",
          1142 => x"82",
          1143 => x"f0",
          1144 => x"e0",
          1145 => x"05",
          1146 => x"a4",
          1147 => x"08",
          1148 => x"54",
          1149 => x"aa",
          1150 => x"e0",
          1151 => x"72",
          1152 => x"e0",
          1153 => x"05",
          1154 => x"a4",
          1155 => x"0c",
          1156 => x"08",
          1157 => x"70",
          1158 => x"89",
          1159 => x"38",
          1160 => x"08",
          1161 => x"53",
          1162 => x"82",
          1163 => x"f8",
          1164 => x"15",
          1165 => x"51",
          1166 => x"e0",
          1167 => x"05",
          1168 => x"82",
          1169 => x"f0",
          1170 => x"72",
          1171 => x"51",
          1172 => x"e0",
          1173 => x"05",
          1174 => x"a4",
          1175 => x"08",
          1176 => x"a4",
          1177 => x"33",
          1178 => x"e0",
          1179 => x"05",
          1180 => x"82",
          1181 => x"f0",
          1182 => x"e0",
          1183 => x"05",
          1184 => x"82",
          1185 => x"fc",
          1186 => x"53",
          1187 => x"82",
          1188 => x"70",
          1189 => x"08",
          1190 => x"53",
          1191 => x"08",
          1192 => x"80",
          1193 => x"fe",
          1194 => x"e0",
          1195 => x"05",
          1196 => x"a8",
          1197 => x"54",
          1198 => x"31",
          1199 => x"82",
          1200 => x"fc",
          1201 => x"e0",
          1202 => x"05",
          1203 => x"06",
          1204 => x"80",
          1205 => x"82",
          1206 => x"ec",
          1207 => x"11",
          1208 => x"82",
          1209 => x"ec",
          1210 => x"e0",
          1211 => x"05",
          1212 => x"2a",
          1213 => x"51",
          1214 => x"80",
          1215 => x"38",
          1216 => x"08",
          1217 => x"70",
          1218 => x"e0",
          1219 => x"05",
          1220 => x"a4",
          1221 => x"08",
          1222 => x"e0",
          1223 => x"05",
          1224 => x"a4",
          1225 => x"22",
          1226 => x"90",
          1227 => x"06",
          1228 => x"e0",
          1229 => x"05",
          1230 => x"53",
          1231 => x"a4",
          1232 => x"23",
          1233 => x"e0",
          1234 => x"05",
          1235 => x"53",
          1236 => x"a4",
          1237 => x"23",
          1238 => x"08",
          1239 => x"82",
          1240 => x"ec",
          1241 => x"e0",
          1242 => x"05",
          1243 => x"2a",
          1244 => x"51",
          1245 => x"80",
          1246 => x"38",
          1247 => x"08",
          1248 => x"70",
          1249 => x"98",
          1250 => x"a4",
          1251 => x"33",
          1252 => x"53",
          1253 => x"97",
          1254 => x"a4",
          1255 => x"22",
          1256 => x"51",
          1257 => x"e0",
          1258 => x"05",
          1259 => x"82",
          1260 => x"e8",
          1261 => x"82",
          1262 => x"fc",
          1263 => x"71",
          1264 => x"72",
          1265 => x"08",
          1266 => x"82",
          1267 => x"e4",
          1268 => x"83",
          1269 => x"06",
          1270 => x"72",
          1271 => x"38",
          1272 => x"08",
          1273 => x"70",
          1274 => x"90",
          1275 => x"2c",
          1276 => x"51",
          1277 => x"53",
          1278 => x"e0",
          1279 => x"05",
          1280 => x"31",
          1281 => x"82",
          1282 => x"ec",
          1283 => x"39",
          1284 => x"08",
          1285 => x"70",
          1286 => x"90",
          1287 => x"2c",
          1288 => x"51",
          1289 => x"53",
          1290 => x"e0",
          1291 => x"05",
          1292 => x"31",
          1293 => x"82",
          1294 => x"ec",
          1295 => x"e0",
          1296 => x"05",
          1297 => x"80",
          1298 => x"72",
          1299 => x"e0",
          1300 => x"05",
          1301 => x"54",
          1302 => x"e0",
          1303 => x"05",
          1304 => x"2b",
          1305 => x"51",
          1306 => x"25",
          1307 => x"e0",
          1308 => x"05",
          1309 => x"51",
          1310 => x"d2",
          1311 => x"a4",
          1312 => x"22",
          1313 => x"70",
          1314 => x"51",
          1315 => x"2e",
          1316 => x"e0",
          1317 => x"05",
          1318 => x"51",
          1319 => x"80",
          1320 => x"e0",
          1321 => x"05",
          1322 => x"2a",
          1323 => x"51",
          1324 => x"80",
          1325 => x"82",
          1326 => x"88",
          1327 => x"ab",
          1328 => x"3f",
          1329 => x"e0",
          1330 => x"05",
          1331 => x"2a",
          1332 => x"51",
          1333 => x"80",
          1334 => x"82",
          1335 => x"88",
          1336 => x"a0",
          1337 => x"3f",
          1338 => x"08",
          1339 => x"70",
          1340 => x"81",
          1341 => x"53",
          1342 => x"b1",
          1343 => x"a4",
          1344 => x"08",
          1345 => x"89",
          1346 => x"e0",
          1347 => x"05",
          1348 => x"90",
          1349 => x"06",
          1350 => x"e0",
          1351 => x"05",
          1352 => x"e0",
          1353 => x"05",
          1354 => x"bc",
          1355 => x"a4",
          1356 => x"22",
          1357 => x"70",
          1358 => x"51",
          1359 => x"2e",
          1360 => x"e0",
          1361 => x"05",
          1362 => x"54",
          1363 => x"e0",
          1364 => x"05",
          1365 => x"2b",
          1366 => x"51",
          1367 => x"25",
          1368 => x"e0",
          1369 => x"05",
          1370 => x"51",
          1371 => x"d2",
          1372 => x"a4",
          1373 => x"22",
          1374 => x"70",
          1375 => x"51",
          1376 => x"2e",
          1377 => x"e0",
          1378 => x"05",
          1379 => x"54",
          1380 => x"e0",
          1381 => x"05",
          1382 => x"2b",
          1383 => x"51",
          1384 => x"25",
          1385 => x"e0",
          1386 => x"05",
          1387 => x"51",
          1388 => x"d2",
          1389 => x"a4",
          1390 => x"22",
          1391 => x"70",
          1392 => x"51",
          1393 => x"38",
          1394 => x"08",
          1395 => x"ff",
          1396 => x"72",
          1397 => x"08",
          1398 => x"73",
          1399 => x"90",
          1400 => x"80",
          1401 => x"38",
          1402 => x"08",
          1403 => x"52",
          1404 => x"f4",
          1405 => x"82",
          1406 => x"f8",
          1407 => x"72",
          1408 => x"09",
          1409 => x"38",
          1410 => x"08",
          1411 => x"52",
          1412 => x"08",
          1413 => x"51",
          1414 => x"81",
          1415 => x"e0",
          1416 => x"05",
          1417 => x"80",
          1418 => x"81",
          1419 => x"38",
          1420 => x"08",
          1421 => x"ff",
          1422 => x"72",
          1423 => x"08",
          1424 => x"72",
          1425 => x"06",
          1426 => x"ff",
          1427 => x"bb",
          1428 => x"a4",
          1429 => x"08",
          1430 => x"a4",
          1431 => x"08",
          1432 => x"82",
          1433 => x"fc",
          1434 => x"05",
          1435 => x"08",
          1436 => x"53",
          1437 => x"ff",
          1438 => x"e0",
          1439 => x"05",
          1440 => x"80",
          1441 => x"81",
          1442 => x"38",
          1443 => x"08",
          1444 => x"ff",
          1445 => x"72",
          1446 => x"08",
          1447 => x"72",
          1448 => x"06",
          1449 => x"ff",
          1450 => x"df",
          1451 => x"a4",
          1452 => x"08",
          1453 => x"a4",
          1454 => x"08",
          1455 => x"53",
          1456 => x"82",
          1457 => x"fc",
          1458 => x"05",
          1459 => x"08",
          1460 => x"ff",
          1461 => x"e0",
          1462 => x"05",
          1463 => x"a8",
          1464 => x"82",
          1465 => x"88",
          1466 => x"82",
          1467 => x"f0",
          1468 => x"05",
          1469 => x"08",
          1470 => x"82",
          1471 => x"f0",
          1472 => x"33",
          1473 => x"e0",
          1474 => x"82",
          1475 => x"e4",
          1476 => x"87",
          1477 => x"06",
          1478 => x"72",
          1479 => x"c3",
          1480 => x"a4",
          1481 => x"22",
          1482 => x"54",
          1483 => x"a4",
          1484 => x"23",
          1485 => x"70",
          1486 => x"53",
          1487 => x"a3",
          1488 => x"a4",
          1489 => x"08",
          1490 => x"85",
          1491 => x"39",
          1492 => x"08",
          1493 => x"52",
          1494 => x"08",
          1495 => x"51",
          1496 => x"80",
          1497 => x"a4",
          1498 => x"23",
          1499 => x"82",
          1500 => x"f8",
          1501 => x"72",
          1502 => x"81",
          1503 => x"81",
          1504 => x"a4",
          1505 => x"23",
          1506 => x"e0",
          1507 => x"05",
          1508 => x"82",
          1509 => x"e8",
          1510 => x"0b",
          1511 => x"08",
          1512 => x"ea",
          1513 => x"e0",
          1514 => x"05",
          1515 => x"e0",
          1516 => x"05",
          1517 => x"b0",
          1518 => x"39",
          1519 => x"08",
          1520 => x"8c",
          1521 => x"82",
          1522 => x"e0",
          1523 => x"53",
          1524 => x"08",
          1525 => x"82",
          1526 => x"95",
          1527 => x"e0",
          1528 => x"82",
          1529 => x"02",
          1530 => x"0c",
          1531 => x"82",
          1532 => x"53",
          1533 => x"08",
          1534 => x"52",
          1535 => x"08",
          1536 => x"51",
          1537 => x"82",
          1538 => x"70",
          1539 => x"0c",
          1540 => x"0d",
          1541 => x"0c",
          1542 => x"a4",
          1543 => x"e0",
          1544 => x"3d",
          1545 => x"82",
          1546 => x"f8",
          1547 => x"fb",
          1548 => x"11",
          1549 => x"2a",
          1550 => x"70",
          1551 => x"51",
          1552 => x"72",
          1553 => x"38",
          1554 => x"e0",
          1555 => x"05",
          1556 => x"39",
          1557 => x"08",
          1558 => x"53",
          1559 => x"e0",
          1560 => x"05",
          1561 => x"82",
          1562 => x"88",
          1563 => x"72",
          1564 => x"08",
          1565 => x"72",
          1566 => x"53",
          1567 => x"b0",
          1568 => x"fc",
          1569 => x"fc",
          1570 => x"e0",
          1571 => x"05",
          1572 => x"11",
          1573 => x"72",
          1574 => x"98",
          1575 => x"80",
          1576 => x"38",
          1577 => x"e0",
          1578 => x"05",
          1579 => x"39",
          1580 => x"08",
          1581 => x"08",
          1582 => x"51",
          1583 => x"53",
          1584 => x"e0",
          1585 => x"72",
          1586 => x"38",
          1587 => x"e0",
          1588 => x"05",
          1589 => x"a4",
          1590 => x"08",
          1591 => x"a4",
          1592 => x"0c",
          1593 => x"a4",
          1594 => x"08",
          1595 => x"0c",
          1596 => x"82",
          1597 => x"04",
          1598 => x"08",
          1599 => x"a4",
          1600 => x"0d",
          1601 => x"e0",
          1602 => x"05",
          1603 => x"a4",
          1604 => x"08",
          1605 => x"70",
          1606 => x"81",
          1607 => x"06",
          1608 => x"51",
          1609 => x"2e",
          1610 => x"0b",
          1611 => x"08",
          1612 => x"80",
          1613 => x"e0",
          1614 => x"05",
          1615 => x"33",
          1616 => x"08",
          1617 => x"81",
          1618 => x"a4",
          1619 => x"0c",
          1620 => x"e0",
          1621 => x"05",
          1622 => x"ff",
          1623 => x"80",
          1624 => x"82",
          1625 => x"8c",
          1626 => x"e0",
          1627 => x"05",
          1628 => x"e0",
          1629 => x"05",
          1630 => x"11",
          1631 => x"72",
          1632 => x"98",
          1633 => x"80",
          1634 => x"38",
          1635 => x"e0",
          1636 => x"05",
          1637 => x"39",
          1638 => x"08",
          1639 => x"70",
          1640 => x"08",
          1641 => x"53",
          1642 => x"08",
          1643 => x"82",
          1644 => x"87",
          1645 => x"e0",
          1646 => x"82",
          1647 => x"02",
          1648 => x"0c",
          1649 => x"82",
          1650 => x"52",
          1651 => x"08",
          1652 => x"51",
          1653 => x"e0",
          1654 => x"82",
          1655 => x"53",
          1656 => x"82",
          1657 => x"04",
          1658 => x"08",
          1659 => x"a4",
          1660 => x"0d",
          1661 => x"08",
          1662 => x"85",
          1663 => x"81",
          1664 => x"32",
          1665 => x"51",
          1666 => x"53",
          1667 => x"8d",
          1668 => x"82",
          1669 => x"fc",
          1670 => x"cb",
          1671 => x"a4",
          1672 => x"08",
          1673 => x"70",
          1674 => x"81",
          1675 => x"51",
          1676 => x"2e",
          1677 => x"82",
          1678 => x"8c",
          1679 => x"e0",
          1680 => x"05",
          1681 => x"8c",
          1682 => x"14",
          1683 => x"38",
          1684 => x"08",
          1685 => x"70",
          1686 => x"e0",
          1687 => x"05",
          1688 => x"54",
          1689 => x"34",
          1690 => x"05",
          1691 => x"e0",
          1692 => x"05",
          1693 => x"08",
          1694 => x"12",
          1695 => x"a4",
          1696 => x"08",
          1697 => x"a4",
          1698 => x"0c",
          1699 => x"d7",
          1700 => x"a4",
          1701 => x"08",
          1702 => x"08",
          1703 => x"53",
          1704 => x"08",
          1705 => x"70",
          1706 => x"53",
          1707 => x"51",
          1708 => x"2d",
          1709 => x"08",
          1710 => x"38",
          1711 => x"08",
          1712 => x"8c",
          1713 => x"05",
          1714 => x"82",
          1715 => x"88",
          1716 => x"82",
          1717 => x"fc",
          1718 => x"53",
          1719 => x"0b",
          1720 => x"08",
          1721 => x"82",
          1722 => x"fc",
          1723 => x"e0",
          1724 => x"3d",
          1725 => x"a4",
          1726 => x"e0",
          1727 => x"82",
          1728 => x"f9",
          1729 => x"e0",
          1730 => x"05",
          1731 => x"33",
          1732 => x"70",
          1733 => x"51",
          1734 => x"80",
          1735 => x"ff",
          1736 => x"a4",
          1737 => x"0c",
          1738 => x"82",
          1739 => x"88",
          1740 => x"11",
          1741 => x"2a",
          1742 => x"51",
          1743 => x"71",
          1744 => x"c5",
          1745 => x"a4",
          1746 => x"08",
          1747 => x"08",
          1748 => x"53",
          1749 => x"33",
          1750 => x"06",
          1751 => x"85",
          1752 => x"e0",
          1753 => x"05",
          1754 => x"08",
          1755 => x"12",
          1756 => x"a4",
          1757 => x"08",
          1758 => x"70",
          1759 => x"08",
          1760 => x"51",
          1761 => x"b6",
          1762 => x"a4",
          1763 => x"08",
          1764 => x"70",
          1765 => x"81",
          1766 => x"51",
          1767 => x"2e",
          1768 => x"82",
          1769 => x"88",
          1770 => x"08",
          1771 => x"e0",
          1772 => x"05",
          1773 => x"82",
          1774 => x"fc",
          1775 => x"38",
          1776 => x"08",
          1777 => x"82",
          1778 => x"88",
          1779 => x"53",
          1780 => x"70",
          1781 => x"52",
          1782 => x"34",
          1783 => x"e0",
          1784 => x"05",
          1785 => x"39",
          1786 => x"08",
          1787 => x"70",
          1788 => x"71",
          1789 => x"a1",
          1790 => x"a4",
          1791 => x"08",
          1792 => x"08",
          1793 => x"52",
          1794 => x"51",
          1795 => x"82",
          1796 => x"70",
          1797 => x"08",
          1798 => x"52",
          1799 => x"08",
          1800 => x"80",
          1801 => x"38",
          1802 => x"08",
          1803 => x"82",
          1804 => x"f4",
          1805 => x"e0",
          1806 => x"05",
          1807 => x"33",
          1808 => x"08",
          1809 => x"52",
          1810 => x"08",
          1811 => x"ff",
          1812 => x"06",
          1813 => x"e0",
          1814 => x"05",
          1815 => x"52",
          1816 => x"a4",
          1817 => x"34",
          1818 => x"e0",
          1819 => x"05",
          1820 => x"52",
          1821 => x"a4",
          1822 => x"34",
          1823 => x"08",
          1824 => x"52",
          1825 => x"08",
          1826 => x"85",
          1827 => x"0b",
          1828 => x"08",
          1829 => x"a6",
          1830 => x"a4",
          1831 => x"08",
          1832 => x"81",
          1833 => x"0c",
          1834 => x"08",
          1835 => x"70",
          1836 => x"70",
          1837 => x"08",
          1838 => x"51",
          1839 => x"e0",
          1840 => x"05",
          1841 => x"98",
          1842 => x"0d",
          1843 => x"0c",
          1844 => x"a4",
          1845 => x"e0",
          1846 => x"3d",
          1847 => x"a4",
          1848 => x"08",
          1849 => x"08",
          1850 => x"82",
          1851 => x"8c",
          1852 => x"e0",
          1853 => x"05",
          1854 => x"a4",
          1855 => x"08",
          1856 => x"a2",
          1857 => x"a4",
          1858 => x"08",
          1859 => x"08",
          1860 => x"26",
          1861 => x"82",
          1862 => x"f8",
          1863 => x"e0",
          1864 => x"05",
          1865 => x"82",
          1866 => x"fc",
          1867 => x"27",
          1868 => x"82",
          1869 => x"fc",
          1870 => x"e0",
          1871 => x"05",
          1872 => x"e0",
          1873 => x"05",
          1874 => x"a4",
          1875 => x"08",
          1876 => x"08",
          1877 => x"05",
          1878 => x"08",
          1879 => x"82",
          1880 => x"90",
          1881 => x"05",
          1882 => x"08",
          1883 => x"82",
          1884 => x"90",
          1885 => x"05",
          1886 => x"08",
          1887 => x"82",
          1888 => x"90",
          1889 => x"2e",
          1890 => x"82",
          1891 => x"fc",
          1892 => x"05",
          1893 => x"08",
          1894 => x"82",
          1895 => x"f8",
          1896 => x"05",
          1897 => x"08",
          1898 => x"82",
          1899 => x"fc",
          1900 => x"e0",
          1901 => x"05",
          1902 => x"71",
          1903 => x"ff",
          1904 => x"e0",
          1905 => x"05",
          1906 => x"82",
          1907 => x"90",
          1908 => x"e0",
          1909 => x"05",
          1910 => x"82",
          1911 => x"90",
          1912 => x"e0",
          1913 => x"05",
          1914 => x"ba",
          1915 => x"a4",
          1916 => x"08",
          1917 => x"82",
          1918 => x"f8",
          1919 => x"05",
          1920 => x"08",
          1921 => x"82",
          1922 => x"fc",
          1923 => x"52",
          1924 => x"82",
          1925 => x"fc",
          1926 => x"05",
          1927 => x"08",
          1928 => x"ff",
          1929 => x"e0",
          1930 => x"05",
          1931 => x"e0",
          1932 => x"85",
          1933 => x"e0",
          1934 => x"82",
          1935 => x"02",
          1936 => x"0c",
          1937 => x"82",
          1938 => x"88",
          1939 => x"e0",
          1940 => x"05",
          1941 => x"a4",
          1942 => x"08",
          1943 => x"82",
          1944 => x"fc",
          1945 => x"05",
          1946 => x"08",
          1947 => x"70",
          1948 => x"51",
          1949 => x"2e",
          1950 => x"39",
          1951 => x"08",
          1952 => x"ff",
          1953 => x"a4",
          1954 => x"0c",
          1955 => x"08",
          1956 => x"82",
          1957 => x"88",
          1958 => x"70",
          1959 => x"0c",
          1960 => x"0d",
          1961 => x"0c",
          1962 => x"a4",
          1963 => x"e0",
          1964 => x"3d",
          1965 => x"a4",
          1966 => x"08",
          1967 => x"08",
          1968 => x"82",
          1969 => x"8c",
          1970 => x"71",
          1971 => x"a4",
          1972 => x"08",
          1973 => x"e0",
          1974 => x"05",
          1975 => x"a4",
          1976 => x"08",
          1977 => x"72",
          1978 => x"a4",
          1979 => x"08",
          1980 => x"e0",
          1981 => x"05",
          1982 => x"ff",
          1983 => x"80",
          1984 => x"ff",
          1985 => x"e0",
          1986 => x"05",
          1987 => x"e0",
          1988 => x"84",
          1989 => x"e0",
          1990 => x"82",
          1991 => x"02",
          1992 => x"0c",
          1993 => x"82",
          1994 => x"88",
          1995 => x"e0",
          1996 => x"05",
          1997 => x"a4",
          1998 => x"08",
          1999 => x"08",
          2000 => x"82",
          2001 => x"90",
          2002 => x"2e",
          2003 => x"82",
          2004 => x"90",
          2005 => x"05",
          2006 => x"08",
          2007 => x"82",
          2008 => x"90",
          2009 => x"05",
          2010 => x"08",
          2011 => x"82",
          2012 => x"90",
          2013 => x"2e",
          2014 => x"e0",
          2015 => x"05",
          2016 => x"33",
          2017 => x"08",
          2018 => x"81",
          2019 => x"a4",
          2020 => x"0c",
          2021 => x"08",
          2022 => x"52",
          2023 => x"34",
          2024 => x"08",
          2025 => x"81",
          2026 => x"a4",
          2027 => x"0c",
          2028 => x"82",
          2029 => x"88",
          2030 => x"82",
          2031 => x"51",
          2032 => x"82",
          2033 => x"04",
          2034 => x"08",
          2035 => x"a4",
          2036 => x"0d",
          2037 => x"08",
          2038 => x"80",
          2039 => x"38",
          2040 => x"08",
          2041 => x"52",
          2042 => x"e0",
          2043 => x"05",
          2044 => x"82",
          2045 => x"8c",
          2046 => x"e0",
          2047 => x"05",
          2048 => x"72",
          2049 => x"53",
          2050 => x"71",
          2051 => x"38",
          2052 => x"82",
          2053 => x"88",
          2054 => x"71",
          2055 => x"a4",
          2056 => x"08",
          2057 => x"e0",
          2058 => x"05",
          2059 => x"ff",
          2060 => x"70",
          2061 => x"0b",
          2062 => x"08",
          2063 => x"81",
          2064 => x"e0",
          2065 => x"05",
          2066 => x"82",
          2067 => x"90",
          2068 => x"e0",
          2069 => x"05",
          2070 => x"84",
          2071 => x"39",
          2072 => x"08",
          2073 => x"80",
          2074 => x"38",
          2075 => x"08",
          2076 => x"70",
          2077 => x"70",
          2078 => x"0b",
          2079 => x"08",
          2080 => x"80",
          2081 => x"e0",
          2082 => x"05",
          2083 => x"82",
          2084 => x"8c",
          2085 => x"e0",
          2086 => x"05",
          2087 => x"52",
          2088 => x"38",
          2089 => x"e0",
          2090 => x"05",
          2091 => x"82",
          2092 => x"88",
          2093 => x"33",
          2094 => x"08",
          2095 => x"70",
          2096 => x"31",
          2097 => x"a4",
          2098 => x"0c",
          2099 => x"52",
          2100 => x"80",
          2101 => x"a4",
          2102 => x"0c",
          2103 => x"08",
          2104 => x"82",
          2105 => x"85",
          2106 => x"e0",
          2107 => x"82",
          2108 => x"02",
          2109 => x"0c",
          2110 => x"82",
          2111 => x"8c",
          2112 => x"82",
          2113 => x"88",
          2114 => x"81",
          2115 => x"e0",
          2116 => x"82",
          2117 => x"f8",
          2118 => x"e0",
          2119 => x"05",
          2120 => x"70",
          2121 => x"80",
          2122 => x"82",
          2123 => x"70",
          2124 => x"08",
          2125 => x"54",
          2126 => x"08",
          2127 => x"8c",
          2128 => x"82",
          2129 => x"f4",
          2130 => x"39",
          2131 => x"08",
          2132 => x"82",
          2133 => x"f8",
          2134 => x"54",
          2135 => x"82",
          2136 => x"f8",
          2137 => x"82",
          2138 => x"88",
          2139 => x"82",
          2140 => x"fc",
          2141 => x"fb",
          2142 => x"e0",
          2143 => x"82",
          2144 => x"f4",
          2145 => x"82",
          2146 => x"f4",
          2147 => x"e0",
          2148 => x"3d",
          2149 => x"a4",
          2150 => x"e0",
          2151 => x"82",
          2152 => x"fd",
          2153 => x"e0",
          2154 => x"05",
          2155 => x"a4",
          2156 => x"0c",
          2157 => x"08",
          2158 => x"8d",
          2159 => x"82",
          2160 => x"fc",
          2161 => x"ec",
          2162 => x"a4",
          2163 => x"08",
          2164 => x"82",
          2165 => x"f8",
          2166 => x"05",
          2167 => x"08",
          2168 => x"70",
          2169 => x"51",
          2170 => x"2e",
          2171 => x"e0",
          2172 => x"05",
          2173 => x"82",
          2174 => x"8c",
          2175 => x"e0",
          2176 => x"05",
          2177 => x"84",
          2178 => x"39",
          2179 => x"08",
          2180 => x"ff",
          2181 => x"a4",
          2182 => x"0c",
          2183 => x"08",
          2184 => x"82",
          2185 => x"88",
          2186 => x"70",
          2187 => x"08",
          2188 => x"51",
          2189 => x"08",
          2190 => x"82",
          2191 => x"85",
          2192 => x"e0",
          2193 => x"82",
          2194 => x"02",
          2195 => x"0c",
          2196 => x"82",
          2197 => x"88",
          2198 => x"e0",
          2199 => x"05",
          2200 => x"a4",
          2201 => x"08",
          2202 => x"d4",
          2203 => x"a4",
          2204 => x"08",
          2205 => x"e0",
          2206 => x"05",
          2207 => x"a4",
          2208 => x"08",
          2209 => x"e0",
          2210 => x"05",
          2211 => x"a4",
          2212 => x"08",
          2213 => x"38",
          2214 => x"08",
          2215 => x"51",
          2216 => x"a4",
          2217 => x"08",
          2218 => x"71",
          2219 => x"a4",
          2220 => x"08",
          2221 => x"e0",
          2222 => x"05",
          2223 => x"39",
          2224 => x"08",
          2225 => x"70",
          2226 => x"0c",
          2227 => x"0d",
          2228 => x"0c",
          2229 => x"a4",
          2230 => x"e0",
          2231 => x"3d",
          2232 => x"a4",
          2233 => x"08",
          2234 => x"a4",
          2235 => x"08",
          2236 => x"82",
          2237 => x"70",
          2238 => x"0c",
          2239 => x"0d",
          2240 => x"0c",
          2241 => x"a4",
          2242 => x"e0",
          2243 => x"3d",
          2244 => x"82",
          2245 => x"fc",
          2246 => x"e0",
          2247 => x"05",
          2248 => x"9b",
          2249 => x"a4",
          2250 => x"08",
          2251 => x"3f",
          2252 => x"08",
          2253 => x"a4",
          2254 => x"0c",
          2255 => x"82",
          2256 => x"fc",
          2257 => x"e0",
          2258 => x"05",
          2259 => x"a4",
          2260 => x"08",
          2261 => x"38",
          2262 => x"08",
          2263 => x"51",
          2264 => x"82",
          2265 => x"82",
          2266 => x"e4",
          2267 => x"31",
          2268 => x"08",
          2269 => x"52",
          2270 => x"e0",
          2271 => x"05",
          2272 => x"a4",
          2273 => x"08",
          2274 => x"a4",
          2275 => x"0c",
          2276 => x"08",
          2277 => x"82",
          2278 => x"f8",
          2279 => x"e0",
          2280 => x"05",
          2281 => x"52",
          2282 => x"a4",
          2283 => x"08",
          2284 => x"80",
          2285 => x"a4",
          2286 => x"0c",
          2287 => x"82",
          2288 => x"fc",
          2289 => x"05",
          2290 => x"e0",
          2291 => x"05",
          2292 => x"81",
          2293 => x"82",
          2294 => x"88",
          2295 => x"82",
          2296 => x"e8",
          2297 => x"82",
          2298 => x"e0",
          2299 => x"05",
          2300 => x"82",
          2301 => x"f8",
          2302 => x"e0",
          2303 => x"05",
          2304 => x"a4",
          2305 => x"08",
          2306 => x"a4",
          2307 => x"0c",
          2308 => x"08",
          2309 => x"82",
          2310 => x"f8",
          2311 => x"82",
          2312 => x"88",
          2313 => x"2b",
          2314 => x"08",
          2315 => x"52",
          2316 => x"e0",
          2317 => x"05",
          2318 => x"a4",
          2319 => x"08",
          2320 => x"ab",
          2321 => x"a4",
          2322 => x"08",
          2323 => x"a4",
          2324 => x"08",
          2325 => x"e0",
          2326 => x"05",
          2327 => x"70",
          2328 => x"e0",
          2329 => x"05",
          2330 => x"a4",
          2331 => x"08",
          2332 => x"e0",
          2333 => x"05",
          2334 => x"e0",
          2335 => x"05",
          2336 => x"a4",
          2337 => x"08",
          2338 => x"08",
          2339 => x"31",
          2340 => x"e0",
          2341 => x"05",
          2342 => x"71",
          2343 => x"e0",
          2344 => x"05",
          2345 => x"a4",
          2346 => x"08",
          2347 => x"e0",
          2348 => x"05",
          2349 => x"a4",
          2350 => x"08",
          2351 => x"08",
          2352 => x"06",
          2353 => x"08",
          2354 => x"71",
          2355 => x"a4",
          2356 => x"0c",
          2357 => x"08",
          2358 => x"ff",
          2359 => x"a4",
          2360 => x"0c",
          2361 => x"51",
          2362 => x"53",
          2363 => x"82",
          2364 => x"88",
          2365 => x"70",
          2366 => x"08",
          2367 => x"07",
          2368 => x"08",
          2369 => x"82",
          2370 => x"88",
          2371 => x"82",
          2372 => x"e8",
          2373 => x"52",
          2374 => x"08",
          2375 => x"82",
          2376 => x"8c",
          2377 => x"e0",
          2378 => x"82",
          2379 => x"02",
          2380 => x"0c",
          2381 => x"82",
          2382 => x"88",
          2383 => x"e0",
          2384 => x"05",
          2385 => x"a4",
          2386 => x"08",
          2387 => x"06",
          2388 => x"38",
          2389 => x"e0",
          2390 => x"05",
          2391 => x"80",
          2392 => x"a4",
          2393 => x"0c",
          2394 => x"08",
          2395 => x"82",
          2396 => x"f8",
          2397 => x"0b",
          2398 => x"08",
          2399 => x"31",
          2400 => x"08",
          2401 => x"71",
          2402 => x"a4",
          2403 => x"0c",
          2404 => x"08",
          2405 => x"82",
          2406 => x"f4",
          2407 => x"e0",
          2408 => x"05",
          2409 => x"80",
          2410 => x"70",
          2411 => x"0b",
          2412 => x"08",
          2413 => x"8a",
          2414 => x"82",
          2415 => x"ec",
          2416 => x"e0",
          2417 => x"05",
          2418 => x"a4",
          2419 => x"0c",
          2420 => x"e0",
          2421 => x"05",
          2422 => x"e0",
          2423 => x"05",
          2424 => x"82",
          2425 => x"fc",
          2426 => x"e0",
          2427 => x"05",
          2428 => x"a4",
          2429 => x"08",
          2430 => x"a4",
          2431 => x"0c",
          2432 => x"08",
          2433 => x"81",
          2434 => x"51",
          2435 => x"84",
          2436 => x"a4",
          2437 => x"0c",
          2438 => x"0b",
          2439 => x"08",
          2440 => x"82",
          2441 => x"e8",
          2442 => x"e0",
          2443 => x"05",
          2444 => x"82",
          2445 => x"f8",
          2446 => x"82",
          2447 => x"fc",
          2448 => x"2a",
          2449 => x"08",
          2450 => x"82",
          2451 => x"f4",
          2452 => x"e0",
          2453 => x"05",
          2454 => x"e0",
          2455 => x"05",
          2456 => x"a4",
          2457 => x"08",
          2458 => x"51",
          2459 => x"82",
          2460 => x"a4",
          2461 => x"0c",
          2462 => x"0b",
          2463 => x"08",
          2464 => x"82",
          2465 => x"e4",
          2466 => x"e0",
          2467 => x"05",
          2468 => x"82",
          2469 => x"f8",
          2470 => x"82",
          2471 => x"fc",
          2472 => x"2a",
          2473 => x"08",
          2474 => x"82",
          2475 => x"f4",
          2476 => x"e0",
          2477 => x"05",
          2478 => x"e0",
          2479 => x"05",
          2480 => x"82",
          2481 => x"fc",
          2482 => x"82",
          2483 => x"fc",
          2484 => x"2a",
          2485 => x"70",
          2486 => x"30",
          2487 => x"82",
          2488 => x"f4",
          2489 => x"70",
          2490 => x"98",
          2491 => x"55",
          2492 => x"52",
          2493 => x"3d",
          2494 => x"a4",
          2495 => x"e0",
          2496 => x"82",
          2497 => x"fe",
          2498 => x"e0",
          2499 => x"05",
          2500 => x"e0",
          2501 => x"05",
          2502 => x"e4",
          2503 => x"98",
          2504 => x"e0",
          2505 => x"05",
          2506 => x"e0",
          2507 => x"05",
          2508 => x"70",
          2509 => x"0c",
          2510 => x"84",
          2511 => x"e0",
          2512 => x"82",
          2513 => x"02",
          2514 => x"0c",
          2515 => x"82",
          2516 => x"8c",
          2517 => x"82",
          2518 => x"88",
          2519 => x"93",
          2520 => x"98",
          2521 => x"e0",
          2522 => x"84",
          2523 => x"e0",
          2524 => x"82",
          2525 => x"02",
          2526 => x"0c",
          2527 => x"a0",
          2528 => x"a4",
          2529 => x"0c",
          2530 => x"08",
          2531 => x"80",
          2532 => x"82",
          2533 => x"8c",
          2534 => x"fb",
          2535 => x"e0",
          2536 => x"82",
          2537 => x"e4",
          2538 => x"8f",
          2539 => x"a4",
          2540 => x"08",
          2541 => x"08",
          2542 => x"82",
          2543 => x"88",
          2544 => x"2e",
          2545 => x"e0",
          2546 => x"05",
          2547 => x"db",
          2548 => x"98",
          2549 => x"a4",
          2550 => x"08",
          2551 => x"e0",
          2552 => x"05",
          2553 => x"39",
          2554 => x"08",
          2555 => x"82",
          2556 => x"fc",
          2557 => x"82",
          2558 => x"e0",
          2559 => x"e0",
          2560 => x"05",
          2561 => x"a4",
          2562 => x"0c",
          2563 => x"08",
          2564 => x"ff",
          2565 => x"82",
          2566 => x"f8",
          2567 => x"94",
          2568 => x"a4",
          2569 => x"08",
          2570 => x"a4",
          2571 => x"0c",
          2572 => x"39",
          2573 => x"08",
          2574 => x"ff",
          2575 => x"82",
          2576 => x"f8",
          2577 => x"09",
          2578 => x"38",
          2579 => x"e0",
          2580 => x"05",
          2581 => x"39",
          2582 => x"08",
          2583 => x"81",
          2584 => x"a4",
          2585 => x"0c",
          2586 => x"08",
          2587 => x"82",
          2588 => x"f8",
          2589 => x"82",
          2590 => x"f4",
          2591 => x"e0",
          2592 => x"05",
          2593 => x"a4",
          2594 => x"08",
          2595 => x"a4",
          2596 => x"08",
          2597 => x"e0",
          2598 => x"05",
          2599 => x"0b",
          2600 => x"08",
          2601 => x"82",
          2602 => x"f8",
          2603 => x"2e",
          2604 => x"82",
          2605 => x"f4",
          2606 => x"82",
          2607 => x"fc",
          2608 => x"05",
          2609 => x"08",
          2610 => x"71",
          2611 => x"07",
          2612 => x"08",
          2613 => x"82",
          2614 => x"88",
          2615 => x"70",
          2616 => x"08",
          2617 => x"07",
          2618 => x"08",
          2619 => x"82",
          2620 => x"8c",
          2621 => x"e0",
          2622 => x"05",
          2623 => x"11",
          2624 => x"08",
          2625 => x"ff",
          2626 => x"2c",
          2627 => x"08",
          2628 => x"82",
          2629 => x"ec",
          2630 => x"06",
          2631 => x"08",
          2632 => x"82",
          2633 => x"8c",
          2634 => x"e0",
          2635 => x"05",
          2636 => x"e0",
          2637 => x"05",
          2638 => x"82",
          2639 => x"f4",
          2640 => x"e0",
          2641 => x"05",
          2642 => x"82",
          2643 => x"f8",
          2644 => x"52",
          2645 => x"51",
          2646 => x"cb",
          2647 => x"a4",
          2648 => x"08",
          2649 => x"a4",
          2650 => x"0c",
          2651 => x"a4",
          2652 => x"08",
          2653 => x"0c",
          2654 => x"82",
          2655 => x"04",
          2656 => x"08",
          2657 => x"a4",
          2658 => x"0d",
          2659 => x"e0",
          2660 => x"05",
          2661 => x"a4",
          2662 => x"08",
          2663 => x"08",
          2664 => x"2c",
          2665 => x"08",
          2666 => x"82",
          2667 => x"8c",
          2668 => x"e0",
          2669 => x"05",
          2670 => x"e0",
          2671 => x"05",
          2672 => x"a4",
          2673 => x"08",
          2674 => x"08",
          2675 => x"32",
          2676 => x"a4",
          2677 => x"08",
          2678 => x"a4",
          2679 => x"0c",
          2680 => x"08",
          2681 => x"82",
          2682 => x"f4",
          2683 => x"70",
          2684 => x"08",
          2685 => x"31",
          2686 => x"08",
          2687 => x"82",
          2688 => x"f8",
          2689 => x"e0",
          2690 => x"05",
          2691 => x"e0",
          2692 => x"05",
          2693 => x"a4",
          2694 => x"08",
          2695 => x"a4",
          2696 => x"08",
          2697 => x"f1",
          2698 => x"e0",
          2699 => x"82",
          2700 => x"f8",
          2701 => x"70",
          2702 => x"08",
          2703 => x"31",
          2704 => x"98",
          2705 => x"53",
          2706 => x"82",
          2707 => x"04",
          2708 => x"08",
          2709 => x"a4",
          2710 => x"0d",
          2711 => x"e0",
          2712 => x"05",
          2713 => x"a4",
          2714 => x"08",
          2715 => x"0c",
          2716 => x"08",
          2717 => x"70",
          2718 => x"72",
          2719 => x"82",
          2720 => x"f8",
          2721 => x"81",
          2722 => x"72",
          2723 => x"81",
          2724 => x"82",
          2725 => x"88",
          2726 => x"08",
          2727 => x"0c",
          2728 => x"82",
          2729 => x"f8",
          2730 => x"72",
          2731 => x"81",
          2732 => x"81",
          2733 => x"a4",
          2734 => x"34",
          2735 => x"08",
          2736 => x"70",
          2737 => x"71",
          2738 => x"51",
          2739 => x"82",
          2740 => x"f8",
          2741 => x"e0",
          2742 => x"05",
          2743 => x"b0",
          2744 => x"06",
          2745 => x"82",
          2746 => x"88",
          2747 => x"08",
          2748 => x"0c",
          2749 => x"53",
          2750 => x"e0",
          2751 => x"05",
          2752 => x"a4",
          2753 => x"33",
          2754 => x"08",
          2755 => x"82",
          2756 => x"e8",
          2757 => x"e2",
          2758 => x"82",
          2759 => x"e8",
          2760 => x"f8",
          2761 => x"80",
          2762 => x"0b",
          2763 => x"08",
          2764 => x"82",
          2765 => x"88",
          2766 => x"08",
          2767 => x"0c",
          2768 => x"53",
          2769 => x"e0",
          2770 => x"05",
          2771 => x"39",
          2772 => x"e0",
          2773 => x"05",
          2774 => x"a4",
          2775 => x"08",
          2776 => x"05",
          2777 => x"08",
          2778 => x"33",
          2779 => x"08",
          2780 => x"80",
          2781 => x"e0",
          2782 => x"05",
          2783 => x"a0",
          2784 => x"81",
          2785 => x"a4",
          2786 => x"0c",
          2787 => x"82",
          2788 => x"f8",
          2789 => x"af",
          2790 => x"38",
          2791 => x"08",
          2792 => x"53",
          2793 => x"83",
          2794 => x"80",
          2795 => x"a4",
          2796 => x"0c",
          2797 => x"88",
          2798 => x"a4",
          2799 => x"34",
          2800 => x"e0",
          2801 => x"05",
          2802 => x"73",
          2803 => x"82",
          2804 => x"f8",
          2805 => x"72",
          2806 => x"38",
          2807 => x"0b",
          2808 => x"08",
          2809 => x"82",
          2810 => x"0b",
          2811 => x"08",
          2812 => x"80",
          2813 => x"a4",
          2814 => x"0c",
          2815 => x"08",
          2816 => x"53",
          2817 => x"81",
          2818 => x"e0",
          2819 => x"05",
          2820 => x"e0",
          2821 => x"38",
          2822 => x"08",
          2823 => x"e0",
          2824 => x"72",
          2825 => x"08",
          2826 => x"82",
          2827 => x"f8",
          2828 => x"11",
          2829 => x"82",
          2830 => x"f8",
          2831 => x"e0",
          2832 => x"05",
          2833 => x"73",
          2834 => x"82",
          2835 => x"f8",
          2836 => x"11",
          2837 => x"82",
          2838 => x"f8",
          2839 => x"e0",
          2840 => x"05",
          2841 => x"89",
          2842 => x"80",
          2843 => x"a4",
          2844 => x"0c",
          2845 => x"82",
          2846 => x"f8",
          2847 => x"e0",
          2848 => x"05",
          2849 => x"72",
          2850 => x"38",
          2851 => x"e0",
          2852 => x"05",
          2853 => x"39",
          2854 => x"08",
          2855 => x"70",
          2856 => x"08",
          2857 => x"29",
          2858 => x"08",
          2859 => x"70",
          2860 => x"a4",
          2861 => x"0c",
          2862 => x"08",
          2863 => x"70",
          2864 => x"71",
          2865 => x"51",
          2866 => x"53",
          2867 => x"e0",
          2868 => x"05",
          2869 => x"39",
          2870 => x"08",
          2871 => x"53",
          2872 => x"90",
          2873 => x"a4",
          2874 => x"08",
          2875 => x"a4",
          2876 => x"0c",
          2877 => x"08",
          2878 => x"82",
          2879 => x"fc",
          2880 => x"0c",
          2881 => x"82",
          2882 => x"ec",
          2883 => x"e0",
          2884 => x"05",
          2885 => x"98",
          2886 => x"0d",
          2887 => x"0c",
          2888 => x"a4",
          2889 => x"e0",
          2890 => x"3d",
          2891 => x"82",
          2892 => x"f0",
          2893 => x"e0",
          2894 => x"05",
          2895 => x"73",
          2896 => x"a4",
          2897 => x"08",
          2898 => x"53",
          2899 => x"72",
          2900 => x"08",
          2901 => x"72",
          2902 => x"53",
          2903 => x"09",
          2904 => x"38",
          2905 => x"08",
          2906 => x"70",
          2907 => x"71",
          2908 => x"39",
          2909 => x"08",
          2910 => x"53",
          2911 => x"09",
          2912 => x"38",
          2913 => x"e0",
          2914 => x"05",
          2915 => x"a4",
          2916 => x"08",
          2917 => x"05",
          2918 => x"08",
          2919 => x"33",
          2920 => x"08",
          2921 => x"82",
          2922 => x"f8",
          2923 => x"72",
          2924 => x"81",
          2925 => x"38",
          2926 => x"08",
          2927 => x"70",
          2928 => x"71",
          2929 => x"51",
          2930 => x"82",
          2931 => x"f8",
          2932 => x"e0",
          2933 => x"05",
          2934 => x"a4",
          2935 => x"0c",
          2936 => x"08",
          2937 => x"80",
          2938 => x"38",
          2939 => x"08",
          2940 => x"80",
          2941 => x"38",
          2942 => x"90",
          2943 => x"a4",
          2944 => x"34",
          2945 => x"08",
          2946 => x"70",
          2947 => x"71",
          2948 => x"51",
          2949 => x"82",
          2950 => x"f8",
          2951 => x"a4",
          2952 => x"82",
          2953 => x"f4",
          2954 => x"e0",
          2955 => x"05",
          2956 => x"81",
          2957 => x"70",
          2958 => x"72",
          2959 => x"a4",
          2960 => x"34",
          2961 => x"82",
          2962 => x"f8",
          2963 => x"72",
          2964 => x"38",
          2965 => x"e0",
          2966 => x"05",
          2967 => x"39",
          2968 => x"08",
          2969 => x"53",
          2970 => x"90",
          2971 => x"a4",
          2972 => x"33",
          2973 => x"26",
          2974 => x"39",
          2975 => x"e0",
          2976 => x"05",
          2977 => x"39",
          2978 => x"e0",
          2979 => x"05",
          2980 => x"82",
          2981 => x"f8",
          2982 => x"af",
          2983 => x"38",
          2984 => x"08",
          2985 => x"53",
          2986 => x"83",
          2987 => x"80",
          2988 => x"a4",
          2989 => x"0c",
          2990 => x"8a",
          2991 => x"a4",
          2992 => x"34",
          2993 => x"e0",
          2994 => x"05",
          2995 => x"a4",
          2996 => x"33",
          2997 => x"27",
          2998 => x"82",
          2999 => x"f8",
          3000 => x"80",
          3001 => x"94",
          3002 => x"a4",
          3003 => x"33",
          3004 => x"53",
          3005 => x"a4",
          3006 => x"34",
          3007 => x"08",
          3008 => x"d0",
          3009 => x"72",
          3010 => x"08",
          3011 => x"82",
          3012 => x"f8",
          3013 => x"90",
          3014 => x"38",
          3015 => x"08",
          3016 => x"f9",
          3017 => x"72",
          3018 => x"08",
          3019 => x"82",
          3020 => x"f8",
          3021 => x"72",
          3022 => x"38",
          3023 => x"e0",
          3024 => x"05",
          3025 => x"39",
          3026 => x"08",
          3027 => x"82",
          3028 => x"f4",
          3029 => x"54",
          3030 => x"8d",
          3031 => x"82",
          3032 => x"ec",
          3033 => x"f7",
          3034 => x"a4",
          3035 => x"33",
          3036 => x"a4",
          3037 => x"08",
          3038 => x"a4",
          3039 => x"33",
          3040 => x"e0",
          3041 => x"05",
          3042 => x"a4",
          3043 => x"08",
          3044 => x"05",
          3045 => x"08",
          3046 => x"55",
          3047 => x"82",
          3048 => x"f8",
          3049 => x"a5",
          3050 => x"a4",
          3051 => x"33",
          3052 => x"2e",
          3053 => x"e0",
          3054 => x"05",
          3055 => x"e0",
          3056 => x"05",
          3057 => x"a4",
          3058 => x"08",
          3059 => x"08",
          3060 => x"71",
          3061 => x"0b",
          3062 => x"08",
          3063 => x"82",
          3064 => x"ec",
          3065 => x"e0",
          3066 => x"3d",
          3067 => x"a4",
          3068 => x"3d",
          3069 => x"08",
          3070 => x"59",
          3071 => x"80",
          3072 => x"39",
          3073 => x"0c",
          3074 => x"54",
          3075 => x"74",
          3076 => x"a0",
          3077 => x"06",
          3078 => x"15",
          3079 => x"80",
          3080 => x"29",
          3081 => x"05",
          3082 => x"56",
          3083 => x"82",
          3084 => x"82",
          3085 => x"54",
          3086 => x"08",
          3087 => x"88",
          3088 => x"98",
          3089 => x"84",
          3090 => x"73",
          3091 => x"b4",
          3092 => x"70",
          3093 => x"58",
          3094 => x"27",
          3095 => x"54",
          3096 => x"98",
          3097 => x"0d",
          3098 => x"0b",
          3099 => x"0c",
          3100 => x"0d",
          3101 => x"93",
          3102 => x"38",
          3103 => x"82",
          3104 => x"52",
          3105 => x"82",
          3106 => x"81",
          3107 => x"bd",
          3108 => x"f9",
          3109 => x"80",
          3110 => x"39",
          3111 => x"51",
          3112 => x"82",
          3113 => x"80",
          3114 => x"be",
          3115 => x"dd",
          3116 => x"c4",
          3117 => x"39",
          3118 => x"51",
          3119 => x"82",
          3120 => x"80",
          3121 => x"bf",
          3122 => x"c1",
          3123 => x"9c",
          3124 => x"82",
          3125 => x"b5",
          3126 => x"cc",
          3127 => x"82",
          3128 => x"a9",
          3129 => x"84",
          3130 => x"82",
          3131 => x"9d",
          3132 => x"b4",
          3133 => x"82",
          3134 => x"91",
          3135 => x"e4",
          3136 => x"82",
          3137 => x"85",
          3138 => x"88",
          3139 => x"3f",
          3140 => x"04",
          3141 => x"77",
          3142 => x"74",
          3143 => x"8a",
          3144 => x"75",
          3145 => x"51",
          3146 => x"e8",
          3147 => x"e3",
          3148 => x"e0",
          3149 => x"75",
          3150 => x"3f",
          3151 => x"08",
          3152 => x"75",
          3153 => x"98",
          3154 => x"c2",
          3155 => x"0d",
          3156 => x"0d",
          3157 => x"05",
          3158 => x"33",
          3159 => x"68",
          3160 => x"7a",
          3161 => x"51",
          3162 => x"78",
          3163 => x"ff",
          3164 => x"81",
          3165 => x"07",
          3166 => x"06",
          3167 => x"56",
          3168 => x"38",
          3169 => x"52",
          3170 => x"52",
          3171 => x"99",
          3172 => x"98",
          3173 => x"e0",
          3174 => x"38",
          3175 => x"08",
          3176 => x"88",
          3177 => x"98",
          3178 => x"3d",
          3179 => x"84",
          3180 => x"52",
          3181 => x"97",
          3182 => x"e0",
          3183 => x"82",
          3184 => x"90",
          3185 => x"74",
          3186 => x"38",
          3187 => x"19",
          3188 => x"39",
          3189 => x"05",
          3190 => x"cd",
          3191 => x"70",
          3192 => x"25",
          3193 => x"9f",
          3194 => x"51",
          3195 => x"74",
          3196 => x"38",
          3197 => x"53",
          3198 => x"88",
          3199 => x"51",
          3200 => x"76",
          3201 => x"e0",
          3202 => x"3d",
          3203 => x"3d",
          3204 => x"84",
          3205 => x"33",
          3206 => x"58",
          3207 => x"52",
          3208 => x"ad",
          3209 => x"98",
          3210 => x"76",
          3211 => x"38",
          3212 => x"9c",
          3213 => x"82",
          3214 => x"61",
          3215 => x"82",
          3216 => x"7f",
          3217 => x"78",
          3218 => x"98",
          3219 => x"39",
          3220 => x"82",
          3221 => x"8a",
          3222 => x"f3",
          3223 => x"61",
          3224 => x"05",
          3225 => x"33",
          3226 => x"68",
          3227 => x"5b",
          3228 => x"77",
          3229 => x"f1",
          3230 => x"98",
          3231 => x"06",
          3232 => x"72",
          3233 => x"38",
          3234 => x"80",
          3235 => x"38",
          3236 => x"53",
          3237 => x"a0",
          3238 => x"82",
          3239 => x"ff",
          3240 => x"82",
          3241 => x"ff",
          3242 => x"80",
          3243 => x"27",
          3244 => x"7b",
          3245 => x"38",
          3246 => x"a7",
          3247 => x"39",
          3248 => x"72",
          3249 => x"38",
          3250 => x"82",
          3251 => x"ff",
          3252 => x"89",
          3253 => x"dc",
          3254 => x"b2",
          3255 => x"55",
          3256 => x"74",
          3257 => x"7a",
          3258 => x"72",
          3259 => x"c1",
          3260 => x"ae",
          3261 => x"39",
          3262 => x"51",
          3263 => x"3f",
          3264 => x"a1",
          3265 => x"53",
          3266 => x"8e",
          3267 => x"52",
          3268 => x"51",
          3269 => x"3f",
          3270 => x"c1",
          3271 => x"ad",
          3272 => x"15",
          3273 => x"fc",
          3274 => x"51",
          3275 => x"fe",
          3276 => x"c1",
          3277 => x"ad",
          3278 => x"55",
          3279 => x"80",
          3280 => x"19",
          3281 => x"53",
          3282 => x"7a",
          3283 => x"81",
          3284 => x"9f",
          3285 => x"38",
          3286 => x"73",
          3287 => x"ff",
          3288 => x"72",
          3289 => x"38",
          3290 => x"26",
          3291 => x"fb",
          3292 => x"73",
          3293 => x"82",
          3294 => x"52",
          3295 => x"e8",
          3296 => x"55",
          3297 => x"82",
          3298 => x"c9",
          3299 => x"19",
          3300 => x"59",
          3301 => x"e0",
          3302 => x"98",
          3303 => x"70",
          3304 => x"57",
          3305 => x"09",
          3306 => x"38",
          3307 => x"c8",
          3308 => x"98",
          3309 => x"70",
          3310 => x"a0",
          3311 => x"72",
          3312 => x"30",
          3313 => x"73",
          3314 => x"51",
          3315 => x"57",
          3316 => x"73",
          3317 => x"76",
          3318 => x"b6",
          3319 => x"53",
          3320 => x"fd",
          3321 => x"53",
          3322 => x"98",
          3323 => x"0d",
          3324 => x"0d",
          3325 => x"33",
          3326 => x"cb",
          3327 => x"c1",
          3328 => x"c1",
          3329 => x"ac",
          3330 => x"de",
          3331 => x"a6",
          3332 => x"c2",
          3333 => x"c2",
          3334 => x"de",
          3335 => x"82",
          3336 => x"ff",
          3337 => x"74",
          3338 => x"38",
          3339 => x"86",
          3340 => x"fe",
          3341 => x"c0",
          3342 => x"53",
          3343 => x"81",
          3344 => x"3f",
          3345 => x"51",
          3346 => x"80",
          3347 => x"3f",
          3348 => x"70",
          3349 => x"52",
          3350 => x"92",
          3351 => x"99",
          3352 => x"c2",
          3353 => x"b6",
          3354 => x"99",
          3355 => x"82",
          3356 => x"06",
          3357 => x"80",
          3358 => x"81",
          3359 => x"3f",
          3360 => x"51",
          3361 => x"80",
          3362 => x"3f",
          3363 => x"70",
          3364 => x"52",
          3365 => x"92",
          3366 => x"98",
          3367 => x"c2",
          3368 => x"fa",
          3369 => x"98",
          3370 => x"84",
          3371 => x"06",
          3372 => x"80",
          3373 => x"81",
          3374 => x"3f",
          3375 => x"51",
          3376 => x"80",
          3377 => x"3f",
          3378 => x"70",
          3379 => x"52",
          3380 => x"92",
          3381 => x"98",
          3382 => x"c3",
          3383 => x"be",
          3384 => x"98",
          3385 => x"86",
          3386 => x"06",
          3387 => x"80",
          3388 => x"81",
          3389 => x"3f",
          3390 => x"51",
          3391 => x"80",
          3392 => x"3f",
          3393 => x"70",
          3394 => x"52",
          3395 => x"92",
          3396 => x"97",
          3397 => x"c3",
          3398 => x"82",
          3399 => x"97",
          3400 => x"88",
          3401 => x"06",
          3402 => x"80",
          3403 => x"81",
          3404 => x"3f",
          3405 => x"51",
          3406 => x"80",
          3407 => x"3f",
          3408 => x"84",
          3409 => x"fb",
          3410 => x"02",
          3411 => x"05",
          3412 => x"56",
          3413 => x"75",
          3414 => x"3f",
          3415 => x"db",
          3416 => x"73",
          3417 => x"53",
          3418 => x"52",
          3419 => x"51",
          3420 => x"3f",
          3421 => x"08",
          3422 => x"e0",
          3423 => x"80",
          3424 => x"31",
          3425 => x"73",
          3426 => x"db",
          3427 => x"0b",
          3428 => x"33",
          3429 => x"2e",
          3430 => x"af",
          3431 => x"a8",
          3432 => x"75",
          3433 => x"af",
          3434 => x"98",
          3435 => x"8b",
          3436 => x"98",
          3437 => x"e1",
          3438 => x"82",
          3439 => x"81",
          3440 => x"82",
          3441 => x"82",
          3442 => x"0b",
          3443 => x"9c",
          3444 => x"82",
          3445 => x"06",
          3446 => x"c4",
          3447 => x"52",
          3448 => x"f0",
          3449 => x"82",
          3450 => x"87",
          3451 => x"cd",
          3452 => x"70",
          3453 => x"7e",
          3454 => x"0c",
          3455 => x"7d",
          3456 => x"8a",
          3457 => x"98",
          3458 => x"06",
          3459 => x"2e",
          3460 => x"a3",
          3461 => x"59",
          3462 => x"c4",
          3463 => x"51",
          3464 => x"7d",
          3465 => x"82",
          3466 => x"81",
          3467 => x"82",
          3468 => x"7e",
          3469 => x"82",
          3470 => x"8d",
          3471 => x"70",
          3472 => x"c4",
          3473 => x"a7",
          3474 => x"3d",
          3475 => x"80",
          3476 => x"51",
          3477 => x"b5",
          3478 => x"05",
          3479 => x"3f",
          3480 => x"08",
          3481 => x"90",
          3482 => x"78",
          3483 => x"87",
          3484 => x"80",
          3485 => x"38",
          3486 => x"81",
          3487 => x"bd",
          3488 => x"78",
          3489 => x"ba",
          3490 => x"2e",
          3491 => x"8a",
          3492 => x"80",
          3493 => x"99",
          3494 => x"c0",
          3495 => x"38",
          3496 => x"82",
          3497 => x"c5",
          3498 => x"f9",
          3499 => x"38",
          3500 => x"24",
          3501 => x"80",
          3502 => x"8d",
          3503 => x"f8",
          3504 => x"38",
          3505 => x"78",
          3506 => x"8a",
          3507 => x"81",
          3508 => x"38",
          3509 => x"2e",
          3510 => x"8a",
          3511 => x"81",
          3512 => x"83",
          3513 => x"39",
          3514 => x"80",
          3515 => x"84",
          3516 => x"ad",
          3517 => x"98",
          3518 => x"fe",
          3519 => x"3d",
          3520 => x"53",
          3521 => x"51",
          3522 => x"82",
          3523 => x"80",
          3524 => x"38",
          3525 => x"f8",
          3526 => x"84",
          3527 => x"81",
          3528 => x"98",
          3529 => x"82",
          3530 => x"43",
          3531 => x"51",
          3532 => x"3f",
          3533 => x"5a",
          3534 => x"81",
          3535 => x"59",
          3536 => x"84",
          3537 => x"7a",
          3538 => x"38",
          3539 => x"b5",
          3540 => x"11",
          3541 => x"05",
          3542 => x"3f",
          3543 => x"08",
          3544 => x"de",
          3545 => x"fe",
          3546 => x"ff",
          3547 => x"eb",
          3548 => x"e0",
          3549 => x"2e",
          3550 => x"b5",
          3551 => x"11",
          3552 => x"05",
          3553 => x"3f",
          3554 => x"08",
          3555 => x"b2",
          3556 => x"f8",
          3557 => x"f6",
          3558 => x"79",
          3559 => x"89",
          3560 => x"79",
          3561 => x"5b",
          3562 => x"62",
          3563 => x"eb",
          3564 => x"ff",
          3565 => x"ff",
          3566 => x"ea",
          3567 => x"e0",
          3568 => x"2e",
          3569 => x"b5",
          3570 => x"11",
          3571 => x"05",
          3572 => x"3f",
          3573 => x"08",
          3574 => x"e6",
          3575 => x"fe",
          3576 => x"ff",
          3577 => x"ea",
          3578 => x"e0",
          3579 => x"2e",
          3580 => x"82",
          3581 => x"ff",
          3582 => x"64",
          3583 => x"27",
          3584 => x"70",
          3585 => x"5e",
          3586 => x"7c",
          3587 => x"78",
          3588 => x"79",
          3589 => x"52",
          3590 => x"51",
          3591 => x"3f",
          3592 => x"81",
          3593 => x"d5",
          3594 => x"c3",
          3595 => x"92",
          3596 => x"ff",
          3597 => x"ff",
          3598 => x"e9",
          3599 => x"e0",
          3600 => x"df",
          3601 => x"fc",
          3602 => x"80",
          3603 => x"82",
          3604 => x"45",
          3605 => x"82",
          3606 => x"59",
          3607 => x"88",
          3608 => x"bc",
          3609 => x"39",
          3610 => x"33",
          3611 => x"2e",
          3612 => x"de",
          3613 => x"ab",
          3614 => x"ff",
          3615 => x"80",
          3616 => x"82",
          3617 => x"45",
          3618 => x"de",
          3619 => x"78",
          3620 => x"38",
          3621 => x"08",
          3622 => x"82",
          3623 => x"fc",
          3624 => x"b5",
          3625 => x"11",
          3626 => x"05",
          3627 => x"3f",
          3628 => x"08",
          3629 => x"82",
          3630 => x"59",
          3631 => x"89",
          3632 => x"b8",
          3633 => x"cc",
          3634 => x"fd",
          3635 => x"80",
          3636 => x"82",
          3637 => x"44",
          3638 => x"de",
          3639 => x"78",
          3640 => x"38",
          3641 => x"08",
          3642 => x"82",
          3643 => x"59",
          3644 => x"88",
          3645 => x"d0",
          3646 => x"39",
          3647 => x"33",
          3648 => x"2e",
          3649 => x"de",
          3650 => x"88",
          3651 => x"e4",
          3652 => x"44",
          3653 => x"f8",
          3654 => x"84",
          3655 => x"81",
          3656 => x"98",
          3657 => x"a7",
          3658 => x"5c",
          3659 => x"2e",
          3660 => x"5c",
          3661 => x"70",
          3662 => x"07",
          3663 => x"7f",
          3664 => x"5a",
          3665 => x"2e",
          3666 => x"a0",
          3667 => x"88",
          3668 => x"b0",
          3669 => x"c1",
          3670 => x"64",
          3671 => x"63",
          3672 => x"f1",
          3673 => x"c5",
          3674 => x"b6",
          3675 => x"ff",
          3676 => x"ff",
          3677 => x"e7",
          3678 => x"e0",
          3679 => x"2e",
          3680 => x"b5",
          3681 => x"11",
          3682 => x"05",
          3683 => x"3f",
          3684 => x"08",
          3685 => x"38",
          3686 => x"80",
          3687 => x"79",
          3688 => x"05",
          3689 => x"fe",
          3690 => x"ff",
          3691 => x"e6",
          3692 => x"e0",
          3693 => x"38",
          3694 => x"64",
          3695 => x"52",
          3696 => x"51",
          3697 => x"3f",
          3698 => x"08",
          3699 => x"52",
          3700 => x"a1",
          3701 => x"46",
          3702 => x"78",
          3703 => x"e2",
          3704 => x"27",
          3705 => x"3d",
          3706 => x"53",
          3707 => x"51",
          3708 => x"82",
          3709 => x"80",
          3710 => x"64",
          3711 => x"cf",
          3712 => x"34",
          3713 => x"45",
          3714 => x"82",
          3715 => x"ff",
          3716 => x"ff",
          3717 => x"3d",
          3718 => x"53",
          3719 => x"51",
          3720 => x"82",
          3721 => x"80",
          3722 => x"38",
          3723 => x"f0",
          3724 => x"84",
          3725 => x"98",
          3726 => x"98",
          3727 => x"a6",
          3728 => x"02",
          3729 => x"22",
          3730 => x"05",
          3731 => x"42",
          3732 => x"f0",
          3733 => x"84",
          3734 => x"f4",
          3735 => x"98",
          3736 => x"f7",
          3737 => x"70",
          3738 => x"82",
          3739 => x"ff",
          3740 => x"82",
          3741 => x"53",
          3742 => x"79",
          3743 => x"e3",
          3744 => x"79",
          3745 => x"ae",
          3746 => x"38",
          3747 => x"87",
          3748 => x"05",
          3749 => x"b5",
          3750 => x"11",
          3751 => x"05",
          3752 => x"3f",
          3753 => x"08",
          3754 => x"38",
          3755 => x"80",
          3756 => x"79",
          3757 => x"5b",
          3758 => x"ff",
          3759 => x"c5",
          3760 => x"ba",
          3761 => x"9e",
          3762 => x"fe",
          3763 => x"ff",
          3764 => x"de",
          3765 => x"e0",
          3766 => x"2e",
          3767 => x"b5",
          3768 => x"11",
          3769 => x"05",
          3770 => x"3f",
          3771 => x"08",
          3772 => x"38",
          3773 => x"0c",
          3774 => x"05",
          3775 => x"fe",
          3776 => x"ff",
          3777 => x"de",
          3778 => x"e0",
          3779 => x"38",
          3780 => x"61",
          3781 => x"52",
          3782 => x"51",
          3783 => x"3f",
          3784 => x"08",
          3785 => x"52",
          3786 => x"9e",
          3787 => x"46",
          3788 => x"78",
          3789 => x"8a",
          3790 => x"27",
          3791 => x"3d",
          3792 => x"53",
          3793 => x"51",
          3794 => x"82",
          3795 => x"80",
          3796 => x"61",
          3797 => x"59",
          3798 => x"42",
          3799 => x"82",
          3800 => x"ff",
          3801 => x"ff",
          3802 => x"3d",
          3803 => x"53",
          3804 => x"51",
          3805 => x"82",
          3806 => x"80",
          3807 => x"38",
          3808 => x"c5",
          3809 => x"9d",
          3810 => x"59",
          3811 => x"3d",
          3812 => x"53",
          3813 => x"51",
          3814 => x"82",
          3815 => x"80",
          3816 => x"38",
          3817 => x"c6",
          3818 => x"9c",
          3819 => x"59",
          3820 => x"e0",
          3821 => x"2e",
          3822 => x"82",
          3823 => x"52",
          3824 => x"51",
          3825 => x"3f",
          3826 => x"82",
          3827 => x"ff",
          3828 => x"ff",
          3829 => x"f4",
          3830 => x"c6",
          3831 => x"b8",
          3832 => x"59",
          3833 => x"92",
          3834 => x"d6",
          3835 => x"33",
          3836 => x"2e",
          3837 => x"80",
          3838 => x"51",
          3839 => x"82",
          3840 => x"5d",
          3841 => x"08",
          3842 => x"92",
          3843 => x"98",
          3844 => x"3d",
          3845 => x"51",
          3846 => x"82",
          3847 => x"60",
          3848 => x"5c",
          3849 => x"81",
          3850 => x"e0",
          3851 => x"c4",
          3852 => x"e0",
          3853 => x"26",
          3854 => x"81",
          3855 => x"2e",
          3856 => x"82",
          3857 => x"7a",
          3858 => x"38",
          3859 => x"7a",
          3860 => x"38",
          3861 => x"82",
          3862 => x"7b",
          3863 => x"fc",
          3864 => x"82",
          3865 => x"b5",
          3866 => x"05",
          3867 => x"86",
          3868 => x"7b",
          3869 => x"ff",
          3870 => x"c4",
          3871 => x"39",
          3872 => x"c6",
          3873 => x"53",
          3874 => x"52",
          3875 => x"b0",
          3876 => x"9d",
          3877 => x"39",
          3878 => x"53",
          3879 => x"52",
          3880 => x"b0",
          3881 => x"9d",
          3882 => x"de",
          3883 => x"e0",
          3884 => x"56",
          3885 => x"54",
          3886 => x"53",
          3887 => x"52",
          3888 => x"b0",
          3889 => x"c6",
          3890 => x"98",
          3891 => x"98",
          3892 => x"30",
          3893 => x"80",
          3894 => x"5b",
          3895 => x"7a",
          3896 => x"38",
          3897 => x"7a",
          3898 => x"80",
          3899 => x"81",
          3900 => x"ff",
          3901 => x"7a",
          3902 => x"7f",
          3903 => x"81",
          3904 => x"78",
          3905 => x"ff",
          3906 => x"06",
          3907 => x"c7",
          3908 => x"b6",
          3909 => x"51",
          3910 => x"f2",
          3911 => x"c7",
          3912 => x"b5",
          3913 => x"9a",
          3914 => x"0d",
          3915 => x"e0",
          3916 => x"c0",
          3917 => x"08",
          3918 => x"84",
          3919 => x"51",
          3920 => x"82",
          3921 => x"90",
          3922 => x"55",
          3923 => x"80",
          3924 => x"cb",
          3925 => x"82",
          3926 => x"07",
          3927 => x"c0",
          3928 => x"08",
          3929 => x"84",
          3930 => x"51",
          3931 => x"82",
          3932 => x"90",
          3933 => x"55",
          3934 => x"80",
          3935 => x"ca",
          3936 => x"82",
          3937 => x"07",
          3938 => x"80",
          3939 => x"c0",
          3940 => x"8c",
          3941 => x"87",
          3942 => x"0c",
          3943 => x"5a",
          3944 => x"5b",
          3945 => x"05",
          3946 => x"80",
          3947 => x"f8",
          3948 => x"70",
          3949 => x"70",
          3950 => x"fb",
          3951 => x"8a",
          3952 => x"ee",
          3953 => x"e0",
          3954 => x"cd",
          3955 => x"ec",
          3956 => x"c5",
          3957 => x"b1",
          3958 => x"3f",
          3959 => x"91",
          3960 => x"3f",
          3961 => x"3d",
          3962 => x"08",
          3963 => x"73",
          3964 => x"74",
          3965 => x"38",
          3966 => x"70",
          3967 => x"81",
          3968 => x"81",
          3969 => x"39",
          3970 => x"70",
          3971 => x"81",
          3972 => x"81",
          3973 => x"54",
          3974 => x"81",
          3975 => x"06",
          3976 => x"39",
          3977 => x"80",
          3978 => x"54",
          3979 => x"83",
          3980 => x"70",
          3981 => x"38",
          3982 => x"98",
          3983 => x"52",
          3984 => x"52",
          3985 => x"2e",
          3986 => x"54",
          3987 => x"84",
          3988 => x"38",
          3989 => x"52",
          3990 => x"2e",
          3991 => x"83",
          3992 => x"70",
          3993 => x"30",
          3994 => x"76",
          3995 => x"51",
          3996 => x"88",
          3997 => x"70",
          3998 => x"34",
          3999 => x"72",
          4000 => x"e0",
          4001 => x"3d",
          4002 => x"3d",
          4003 => x"72",
          4004 => x"91",
          4005 => x"fc",
          4006 => x"51",
          4007 => x"82",
          4008 => x"85",
          4009 => x"83",
          4010 => x"72",
          4011 => x"0c",
          4012 => x"04",
          4013 => x"76",
          4014 => x"ff",
          4015 => x"81",
          4016 => x"26",
          4017 => x"83",
          4018 => x"05",
          4019 => x"70",
          4020 => x"8a",
          4021 => x"33",
          4022 => x"70",
          4023 => x"fe",
          4024 => x"33",
          4025 => x"70",
          4026 => x"f2",
          4027 => x"33",
          4028 => x"70",
          4029 => x"e6",
          4030 => x"22",
          4031 => x"74",
          4032 => x"80",
          4033 => x"13",
          4034 => x"52",
          4035 => x"26",
          4036 => x"81",
          4037 => x"98",
          4038 => x"22",
          4039 => x"bc",
          4040 => x"33",
          4041 => x"b8",
          4042 => x"33",
          4043 => x"b4",
          4044 => x"33",
          4045 => x"b0",
          4046 => x"33",
          4047 => x"ac",
          4048 => x"33",
          4049 => x"a8",
          4050 => x"c0",
          4051 => x"73",
          4052 => x"a0",
          4053 => x"87",
          4054 => x"0c",
          4055 => x"82",
          4056 => x"86",
          4057 => x"f3",
          4058 => x"5b",
          4059 => x"9c",
          4060 => x"0c",
          4061 => x"bc",
          4062 => x"7b",
          4063 => x"98",
          4064 => x"79",
          4065 => x"87",
          4066 => x"08",
          4067 => x"1c",
          4068 => x"98",
          4069 => x"79",
          4070 => x"87",
          4071 => x"08",
          4072 => x"1c",
          4073 => x"98",
          4074 => x"79",
          4075 => x"87",
          4076 => x"08",
          4077 => x"1c",
          4078 => x"98",
          4079 => x"79",
          4080 => x"80",
          4081 => x"83",
          4082 => x"59",
          4083 => x"ff",
          4084 => x"1b",
          4085 => x"1b",
          4086 => x"1b",
          4087 => x"1b",
          4088 => x"1b",
          4089 => x"83",
          4090 => x"52",
          4091 => x"51",
          4092 => x"3f",
          4093 => x"04",
          4094 => x"02",
          4095 => x"53",
          4096 => x"81",
          4097 => x"06",
          4098 => x"52",
          4099 => x"70",
          4100 => x"25",
          4101 => x"51",
          4102 => x"2e",
          4103 => x"97",
          4104 => x"84",
          4105 => x"e0",
          4106 => x"2b",
          4107 => x"51",
          4108 => x"2e",
          4109 => x"9e",
          4110 => x"72",
          4111 => x"81",
          4112 => x"72",
          4113 => x"32",
          4114 => x"80",
          4115 => x"51",
          4116 => x"ff",
          4117 => x"82",
          4118 => x"85",
          4119 => x"fd",
          4120 => x"53",
          4121 => x"88",
          4122 => x"51",
          4123 => x"82",
          4124 => x"98",
          4125 => x"2c",
          4126 => x"16",
          4127 => x"73",
          4128 => x"38",
          4129 => x"98",
          4130 => x"0d",
          4131 => x"0d",
          4132 => x"33",
          4133 => x"33",
          4134 => x"06",
          4135 => x"87",
          4136 => x"51",
          4137 => x"86",
          4138 => x"94",
          4139 => x"08",
          4140 => x"70",
          4141 => x"54",
          4142 => x"2e",
          4143 => x"91",
          4144 => x"06",
          4145 => x"d7",
          4146 => x"32",
          4147 => x"51",
          4148 => x"2e",
          4149 => x"93",
          4150 => x"06",
          4151 => x"ff",
          4152 => x"81",
          4153 => x"87",
          4154 => x"52",
          4155 => x"86",
          4156 => x"94",
          4157 => x"72",
          4158 => x"e0",
          4159 => x"3d",
          4160 => x"3d",
          4161 => x"05",
          4162 => x"70",
          4163 => x"52",
          4164 => x"de",
          4165 => x"3d",
          4166 => x"3d",
          4167 => x"05",
          4168 => x"8a",
          4169 => x"06",
          4170 => x"52",
          4171 => x"3f",
          4172 => x"33",
          4173 => x"06",
          4174 => x"c0",
          4175 => x"76",
          4176 => x"38",
          4177 => x"94",
          4178 => x"70",
          4179 => x"81",
          4180 => x"54",
          4181 => x"8c",
          4182 => x"2a",
          4183 => x"51",
          4184 => x"38",
          4185 => x"70",
          4186 => x"53",
          4187 => x"8d",
          4188 => x"2a",
          4189 => x"51",
          4190 => x"be",
          4191 => x"ff",
          4192 => x"c0",
          4193 => x"72",
          4194 => x"38",
          4195 => x"90",
          4196 => x"0c",
          4197 => x"e0",
          4198 => x"3d",
          4199 => x"3d",
          4200 => x"80",
          4201 => x"81",
          4202 => x"53",
          4203 => x"2e",
          4204 => x"71",
          4205 => x"81",
          4206 => x"b0",
          4207 => x"ff",
          4208 => x"55",
          4209 => x"94",
          4210 => x"80",
          4211 => x"87",
          4212 => x"51",
          4213 => x"96",
          4214 => x"06",
          4215 => x"70",
          4216 => x"38",
          4217 => x"70",
          4218 => x"51",
          4219 => x"72",
          4220 => x"81",
          4221 => x"70",
          4222 => x"38",
          4223 => x"70",
          4224 => x"51",
          4225 => x"38",
          4226 => x"06",
          4227 => x"94",
          4228 => x"80",
          4229 => x"87",
          4230 => x"52",
          4231 => x"81",
          4232 => x"70",
          4233 => x"53",
          4234 => x"ff",
          4235 => x"82",
          4236 => x"89",
          4237 => x"fe",
          4238 => x"de",
          4239 => x"81",
          4240 => x"52",
          4241 => x"84",
          4242 => x"2e",
          4243 => x"c0",
          4244 => x"70",
          4245 => x"2a",
          4246 => x"51",
          4247 => x"80",
          4248 => x"71",
          4249 => x"51",
          4250 => x"80",
          4251 => x"2e",
          4252 => x"c0",
          4253 => x"71",
          4254 => x"ff",
          4255 => x"98",
          4256 => x"3d",
          4257 => x"af",
          4258 => x"98",
          4259 => x"06",
          4260 => x"0c",
          4261 => x"0d",
          4262 => x"33",
          4263 => x"06",
          4264 => x"c0",
          4265 => x"70",
          4266 => x"38",
          4267 => x"94",
          4268 => x"70",
          4269 => x"81",
          4270 => x"51",
          4271 => x"80",
          4272 => x"72",
          4273 => x"51",
          4274 => x"80",
          4275 => x"2e",
          4276 => x"c0",
          4277 => x"71",
          4278 => x"2b",
          4279 => x"51",
          4280 => x"82",
          4281 => x"84",
          4282 => x"ff",
          4283 => x"c0",
          4284 => x"70",
          4285 => x"06",
          4286 => x"80",
          4287 => x"38",
          4288 => x"a4",
          4289 => x"b4",
          4290 => x"9e",
          4291 => x"de",
          4292 => x"c0",
          4293 => x"82",
          4294 => x"87",
          4295 => x"08",
          4296 => x"0c",
          4297 => x"9c",
          4298 => x"c4",
          4299 => x"9e",
          4300 => x"de",
          4301 => x"c0",
          4302 => x"82",
          4303 => x"87",
          4304 => x"08",
          4305 => x"0c",
          4306 => x"b4",
          4307 => x"d4",
          4308 => x"9e",
          4309 => x"de",
          4310 => x"c0",
          4311 => x"82",
          4312 => x"87",
          4313 => x"08",
          4314 => x"0c",
          4315 => x"c4",
          4316 => x"e4",
          4317 => x"9e",
          4318 => x"70",
          4319 => x"23",
          4320 => x"84",
          4321 => x"ec",
          4322 => x"9e",
          4323 => x"de",
          4324 => x"c0",
          4325 => x"82",
          4326 => x"81",
          4327 => x"f8",
          4328 => x"87",
          4329 => x"08",
          4330 => x"0a",
          4331 => x"52",
          4332 => x"83",
          4333 => x"71",
          4334 => x"34",
          4335 => x"c0",
          4336 => x"70",
          4337 => x"06",
          4338 => x"70",
          4339 => x"38",
          4340 => x"82",
          4341 => x"80",
          4342 => x"9e",
          4343 => x"90",
          4344 => x"51",
          4345 => x"80",
          4346 => x"81",
          4347 => x"de",
          4348 => x"0b",
          4349 => x"90",
          4350 => x"80",
          4351 => x"52",
          4352 => x"2e",
          4353 => x"52",
          4354 => x"fc",
          4355 => x"87",
          4356 => x"08",
          4357 => x"80",
          4358 => x"52",
          4359 => x"83",
          4360 => x"71",
          4361 => x"34",
          4362 => x"c0",
          4363 => x"70",
          4364 => x"06",
          4365 => x"70",
          4366 => x"38",
          4367 => x"82",
          4368 => x"80",
          4369 => x"9e",
          4370 => x"84",
          4371 => x"51",
          4372 => x"80",
          4373 => x"81",
          4374 => x"de",
          4375 => x"0b",
          4376 => x"90",
          4377 => x"80",
          4378 => x"52",
          4379 => x"2e",
          4380 => x"52",
          4381 => x"80",
          4382 => x"87",
          4383 => x"08",
          4384 => x"80",
          4385 => x"52",
          4386 => x"83",
          4387 => x"71",
          4388 => x"34",
          4389 => x"c0",
          4390 => x"70",
          4391 => x"06",
          4392 => x"70",
          4393 => x"38",
          4394 => x"82",
          4395 => x"80",
          4396 => x"9e",
          4397 => x"a0",
          4398 => x"52",
          4399 => x"2e",
          4400 => x"52",
          4401 => x"83",
          4402 => x"9e",
          4403 => x"98",
          4404 => x"8a",
          4405 => x"51",
          4406 => x"84",
          4407 => x"87",
          4408 => x"08",
          4409 => x"06",
          4410 => x"70",
          4411 => x"38",
          4412 => x"82",
          4413 => x"87",
          4414 => x"08",
          4415 => x"06",
          4416 => x"51",
          4417 => x"82",
          4418 => x"80",
          4419 => x"9e",
          4420 => x"88",
          4421 => x"52",
          4422 => x"83",
          4423 => x"71",
          4424 => x"34",
          4425 => x"90",
          4426 => x"06",
          4427 => x"82",
          4428 => x"83",
          4429 => x"fb",
          4430 => x"c8",
          4431 => x"89",
          4432 => x"de",
          4433 => x"73",
          4434 => x"38",
          4435 => x"51",
          4436 => x"3f",
          4437 => x"51",
          4438 => x"3f",
          4439 => x"33",
          4440 => x"2e",
          4441 => x"de",
          4442 => x"de",
          4443 => x"54",
          4444 => x"dc",
          4445 => x"96",
          4446 => x"ff",
          4447 => x"80",
          4448 => x"82",
          4449 => x"82",
          4450 => x"11",
          4451 => x"c8",
          4452 => x"88",
          4453 => x"de",
          4454 => x"73",
          4455 => x"38",
          4456 => x"08",
          4457 => x"08",
          4458 => x"82",
          4459 => x"ff",
          4460 => x"82",
          4461 => x"54",
          4462 => x"94",
          4463 => x"bc",
          4464 => x"c0",
          4465 => x"52",
          4466 => x"51",
          4467 => x"3f",
          4468 => x"33",
          4469 => x"2e",
          4470 => x"de",
          4471 => x"de",
          4472 => x"54",
          4473 => x"cc",
          4474 => x"a2",
          4475 => x"83",
          4476 => x"80",
          4477 => x"82",
          4478 => x"52",
          4479 => x"51",
          4480 => x"3f",
          4481 => x"33",
          4482 => x"2e",
          4483 => x"df",
          4484 => x"82",
          4485 => x"ff",
          4486 => x"82",
          4487 => x"54",
          4488 => x"8e",
          4489 => x"86",
          4490 => x"ca",
          4491 => x"87",
          4492 => x"de",
          4493 => x"73",
          4494 => x"38",
          4495 => x"51",
          4496 => x"3f",
          4497 => x"33",
          4498 => x"2e",
          4499 => x"ca",
          4500 => x"a3",
          4501 => x"df",
          4502 => x"73",
          4503 => x"38",
          4504 => x"51",
          4505 => x"3f",
          4506 => x"33",
          4507 => x"2e",
          4508 => x"ca",
          4509 => x"a3",
          4510 => x"df",
          4511 => x"73",
          4512 => x"38",
          4513 => x"51",
          4514 => x"3f",
          4515 => x"51",
          4516 => x"3f",
          4517 => x"08",
          4518 => x"90",
          4519 => x"ee",
          4520 => x"e0",
          4521 => x"cb",
          4522 => x"86",
          4523 => x"de",
          4524 => x"82",
          4525 => x"ff",
          4526 => x"82",
          4527 => x"ff",
          4528 => x"82",
          4529 => x"52",
          4530 => x"51",
          4531 => x"3f",
          4532 => x"08",
          4533 => x"c0",
          4534 => x"ff",
          4535 => x"82",
          4536 => x"bd",
          4537 => x"76",
          4538 => x"54",
          4539 => x"08",
          4540 => x"b8",
          4541 => x"96",
          4542 => x"ff",
          4543 => x"80",
          4544 => x"82",
          4545 => x"56",
          4546 => x"52",
          4547 => x"b7",
          4548 => x"e0",
          4549 => x"84",
          4550 => x"71",
          4551 => x"82",
          4552 => x"52",
          4553 => x"51",
          4554 => x"3f",
          4555 => x"33",
          4556 => x"2e",
          4557 => x"de",
          4558 => x"bd",
          4559 => x"75",
          4560 => x"91",
          4561 => x"98",
          4562 => x"c0",
          4563 => x"31",
          4564 => x"e0",
          4565 => x"82",
          4566 => x"ff",
          4567 => x"8a",
          4568 => x"d7",
          4569 => x"0d",
          4570 => x"0d",
          4571 => x"33",
          4572 => x"71",
          4573 => x"38",
          4574 => x"82",
          4575 => x"52",
          4576 => x"82",
          4577 => x"9d",
          4578 => x"c4",
          4579 => x"82",
          4580 => x"91",
          4581 => x"d4",
          4582 => x"82",
          4583 => x"85",
          4584 => x"e0",
          4585 => x"e6",
          4586 => x"0d",
          4587 => x"80",
          4588 => x"0b",
          4589 => x"84",
          4590 => x"df",
          4591 => x"c0",
          4592 => x"04",
          4593 => x"76",
          4594 => x"98",
          4595 => x"2b",
          4596 => x"72",
          4597 => x"82",
          4598 => x"51",
          4599 => x"80",
          4600 => x"ec",
          4601 => x"53",
          4602 => x"9c",
          4603 => x"e8",
          4604 => x"02",
          4605 => x"05",
          4606 => x"52",
          4607 => x"72",
          4608 => x"06",
          4609 => x"53",
          4610 => x"98",
          4611 => x"0d",
          4612 => x"0d",
          4613 => x"05",
          4614 => x"71",
          4615 => x"54",
          4616 => x"b1",
          4617 => x"fc",
          4618 => x"51",
          4619 => x"3f",
          4620 => x"08",
          4621 => x"ff",
          4622 => x"82",
          4623 => x"52",
          4624 => x"a3",
          4625 => x"33",
          4626 => x"72",
          4627 => x"81",
          4628 => x"cc",
          4629 => x"ff",
          4630 => x"74",
          4631 => x"3d",
          4632 => x"3d",
          4633 => x"84",
          4634 => x"33",
          4635 => x"bb",
          4636 => x"df",
          4637 => x"84",
          4638 => x"90",
          4639 => x"51",
          4640 => x"58",
          4641 => x"2e",
          4642 => x"51",
          4643 => x"82",
          4644 => x"70",
          4645 => x"df",
          4646 => x"19",
          4647 => x"56",
          4648 => x"3f",
          4649 => x"08",
          4650 => x"df",
          4651 => x"84",
          4652 => x"90",
          4653 => x"51",
          4654 => x"80",
          4655 => x"75",
          4656 => x"74",
          4657 => x"d3",
          4658 => x"e8",
          4659 => x"55",
          4660 => x"e8",
          4661 => x"ff",
          4662 => x"75",
          4663 => x"80",
          4664 => x"e8",
          4665 => x"2e",
          4666 => x"df",
          4667 => x"75",
          4668 => x"38",
          4669 => x"33",
          4670 => x"38",
          4671 => x"05",
          4672 => x"78",
          4673 => x"80",
          4674 => x"82",
          4675 => x"52",
          4676 => x"a2",
          4677 => x"df",
          4678 => x"80",
          4679 => x"8c",
          4680 => x"fd",
          4681 => x"df",
          4682 => x"54",
          4683 => x"71",
          4684 => x"38",
          4685 => x"d3",
          4686 => x"0c",
          4687 => x"14",
          4688 => x"80",
          4689 => x"80",
          4690 => x"e8",
          4691 => x"e4",
          4692 => x"80",
          4693 => x"71",
          4694 => x"cd",
          4695 => x"e4",
          4696 => x"a7",
          4697 => x"82",
          4698 => x"85",
          4699 => x"dc",
          4700 => x"57",
          4701 => x"df",
          4702 => x"80",
          4703 => x"82",
          4704 => x"80",
          4705 => x"df",
          4706 => x"80",
          4707 => x"3d",
          4708 => x"81",
          4709 => x"82",
          4710 => x"80",
          4711 => x"75",
          4712 => x"97",
          4713 => x"98",
          4714 => x"0b",
          4715 => x"08",
          4716 => x"82",
          4717 => x"ff",
          4718 => x"55",
          4719 => x"34",
          4720 => x"52",
          4721 => x"d0",
          4722 => x"ff",
          4723 => x"74",
          4724 => x"81",
          4725 => x"38",
          4726 => x"04",
          4727 => x"aa",
          4728 => x"3d",
          4729 => x"81",
          4730 => x"80",
          4731 => x"e4",
          4732 => x"f4",
          4733 => x"e0",
          4734 => x"95",
          4735 => x"82",
          4736 => x"54",
          4737 => x"52",
          4738 => x"52",
          4739 => x"c7",
          4740 => x"98",
          4741 => x"a5",
          4742 => x"ff",
          4743 => x"82",
          4744 => x"81",
          4745 => x"80",
          4746 => x"98",
          4747 => x"38",
          4748 => x"08",
          4749 => x"17",
          4750 => x"74",
          4751 => x"70",
          4752 => x"07",
          4753 => x"55",
          4754 => x"2e",
          4755 => x"ff",
          4756 => x"df",
          4757 => x"11",
          4758 => x"80",
          4759 => x"82",
          4760 => x"80",
          4761 => x"82",
          4762 => x"fe",
          4763 => x"78",
          4764 => x"81",
          4765 => x"75",
          4766 => x"ff",
          4767 => x"79",
          4768 => x"b7",
          4769 => x"08",
          4770 => x"98",
          4771 => x"80",
          4772 => x"e0",
          4773 => x"3d",
          4774 => x"3d",
          4775 => x"71",
          4776 => x"33",
          4777 => x"58",
          4778 => x"09",
          4779 => x"38",
          4780 => x"05",
          4781 => x"27",
          4782 => x"17",
          4783 => x"71",
          4784 => x"55",
          4785 => x"09",
          4786 => x"38",
          4787 => x"ea",
          4788 => x"73",
          4789 => x"df",
          4790 => x"08",
          4791 => x"a6",
          4792 => x"e0",
          4793 => x"79",
          4794 => x"51",
          4795 => x"3f",
          4796 => x"08",
          4797 => x"84",
          4798 => x"74",
          4799 => x"38",
          4800 => x"88",
          4801 => x"fc",
          4802 => x"39",
          4803 => x"8c",
          4804 => x"53",
          4805 => x"c4",
          4806 => x"e0",
          4807 => x"2e",
          4808 => x"1b",
          4809 => x"77",
          4810 => x"3f",
          4811 => x"08",
          4812 => x"55",
          4813 => x"74",
          4814 => x"81",
          4815 => x"ff",
          4816 => x"82",
          4817 => x"8b",
          4818 => x"73",
          4819 => x"0c",
          4820 => x"04",
          4821 => x"b0",
          4822 => x"3d",
          4823 => x"08",
          4824 => x"80",
          4825 => x"34",
          4826 => x"33",
          4827 => x"08",
          4828 => x"81",
          4829 => x"82",
          4830 => x"55",
          4831 => x"38",
          4832 => x"80",
          4833 => x"38",
          4834 => x"06",
          4835 => x"80",
          4836 => x"38",
          4837 => x"89",
          4838 => x"98",
          4839 => x"e4",
          4840 => x"98",
          4841 => x"81",
          4842 => x"53",
          4843 => x"e0",
          4844 => x"80",
          4845 => x"82",
          4846 => x"80",
          4847 => x"82",
          4848 => x"ff",
          4849 => x"80",
          4850 => x"e0",
          4851 => x"82",
          4852 => x"53",
          4853 => x"90",
          4854 => x"54",
          4855 => x"3f",
          4856 => x"08",
          4857 => x"98",
          4858 => x"09",
          4859 => x"d0",
          4860 => x"98",
          4861 => x"a4",
          4862 => x"e0",
          4863 => x"80",
          4864 => x"98",
          4865 => x"38",
          4866 => x"08",
          4867 => x"17",
          4868 => x"74",
          4869 => x"74",
          4870 => x"52",
          4871 => x"c2",
          4872 => x"70",
          4873 => x"5c",
          4874 => x"27",
          4875 => x"5b",
          4876 => x"09",
          4877 => x"97",
          4878 => x"75",
          4879 => x"34",
          4880 => x"82",
          4881 => x"80",
          4882 => x"f9",
          4883 => x"3d",
          4884 => x"e7",
          4885 => x"e0",
          4886 => x"2b",
          4887 => x"51",
          4888 => x"2e",
          4889 => x"81",
          4890 => x"f7",
          4891 => x"98",
          4892 => x"2c",
          4893 => x"33",
          4894 => x"70",
          4895 => x"98",
          4896 => x"84",
          4897 => x"e8",
          4898 => x"15",
          4899 => x"51",
          4900 => x"59",
          4901 => x"58",
          4902 => x"78",
          4903 => x"38",
          4904 => x"b4",
          4905 => x"80",
          4906 => x"ff",
          4907 => x"98",
          4908 => x"80",
          4909 => x"ce",
          4910 => x"74",
          4911 => x"f6",
          4912 => x"e0",
          4913 => x"ff",
          4914 => x"80",
          4915 => x"74",
          4916 => x"34",
          4917 => x"39",
          4918 => x"0a",
          4919 => x"0a",
          4920 => x"2c",
          4921 => x"06",
          4922 => x"73",
          4923 => x"38",
          4924 => x"52",
          4925 => x"cc",
          4926 => x"98",
          4927 => x"06",
          4928 => x"38",
          4929 => x"56",
          4930 => x"80",
          4931 => x"1c",
          4932 => x"f7",
          4933 => x"98",
          4934 => x"2c",
          4935 => x"33",
          4936 => x"70",
          4937 => x"10",
          4938 => x"2b",
          4939 => x"11",
          4940 => x"51",
          4941 => x"51",
          4942 => x"2e",
          4943 => x"fe",
          4944 => x"cd",
          4945 => x"7d",
          4946 => x"82",
          4947 => x"80",
          4948 => x"d0",
          4949 => x"75",
          4950 => x"34",
          4951 => x"d0",
          4952 => x"3d",
          4953 => x"0c",
          4954 => x"95",
          4955 => x"38",
          4956 => x"82",
          4957 => x"54",
          4958 => x"82",
          4959 => x"54",
          4960 => x"fd",
          4961 => x"f7",
          4962 => x"73",
          4963 => x"38",
          4964 => x"70",
          4965 => x"55",
          4966 => x"9e",
          4967 => x"54",
          4968 => x"15",
          4969 => x"80",
          4970 => x"ff",
          4971 => x"98",
          4972 => x"dc",
          4973 => x"55",
          4974 => x"f7",
          4975 => x"11",
          4976 => x"82",
          4977 => x"73",
          4978 => x"3d",
          4979 => x"82",
          4980 => x"54",
          4981 => x"89",
          4982 => x"54",
          4983 => x"d8",
          4984 => x"dc",
          4985 => x"80",
          4986 => x"ff",
          4987 => x"98",
          4988 => x"d8",
          4989 => x"56",
          4990 => x"25",
          4991 => x"fb",
          4992 => x"74",
          4993 => x"52",
          4994 => x"dc",
          4995 => x"80",
          4996 => x"80",
          4997 => x"98",
          4998 => x"d8",
          4999 => x"55",
          5000 => x"da",
          5001 => x"dc",
          5002 => x"2b",
          5003 => x"82",
          5004 => x"5a",
          5005 => x"74",
          5006 => x"92",
          5007 => x"fc",
          5008 => x"51",
          5009 => x"3f",
          5010 => x"0a",
          5011 => x"0a",
          5012 => x"2c",
          5013 => x"33",
          5014 => x"73",
          5015 => x"38",
          5016 => x"83",
          5017 => x"0b",
          5018 => x"82",
          5019 => x"80",
          5020 => x"b8",
          5021 => x"3f",
          5022 => x"82",
          5023 => x"70",
          5024 => x"55",
          5025 => x"2e",
          5026 => x"82",
          5027 => x"ff",
          5028 => x"82",
          5029 => x"ff",
          5030 => x"82",
          5031 => x"82",
          5032 => x"52",
          5033 => x"96",
          5034 => x"f7",
          5035 => x"98",
          5036 => x"2c",
          5037 => x"33",
          5038 => x"57",
          5039 => x"ad",
          5040 => x"54",
          5041 => x"74",
          5042 => x"fc",
          5043 => x"33",
          5044 => x"94",
          5045 => x"80",
          5046 => x"80",
          5047 => x"98",
          5048 => x"d8",
          5049 => x"55",
          5050 => x"d5",
          5051 => x"fc",
          5052 => x"51",
          5053 => x"3f",
          5054 => x"33",
          5055 => x"70",
          5056 => x"f7",
          5057 => x"51",
          5058 => x"74",
          5059 => x"38",
          5060 => x"08",
          5061 => x"ff",
          5062 => x"74",
          5063 => x"29",
          5064 => x"05",
          5065 => x"82",
          5066 => x"58",
          5067 => x"75",
          5068 => x"fa",
          5069 => x"f7",
          5070 => x"05",
          5071 => x"34",
          5072 => x"08",
          5073 => x"ff",
          5074 => x"82",
          5075 => x"79",
          5076 => x"3f",
          5077 => x"08",
          5078 => x"54",
          5079 => x"82",
          5080 => x"54",
          5081 => x"8f",
          5082 => x"73",
          5083 => x"f1",
          5084 => x"39",
          5085 => x"80",
          5086 => x"dc",
          5087 => x"82",
          5088 => x"79",
          5089 => x"0c",
          5090 => x"04",
          5091 => x"33",
          5092 => x"2e",
          5093 => x"82",
          5094 => x"52",
          5095 => x"94",
          5096 => x"f7",
          5097 => x"05",
          5098 => x"f7",
          5099 => x"81",
          5100 => x"dd",
          5101 => x"dc",
          5102 => x"d8",
          5103 => x"73",
          5104 => x"8a",
          5105 => x"54",
          5106 => x"d8",
          5107 => x"2b",
          5108 => x"75",
          5109 => x"56",
          5110 => x"74",
          5111 => x"74",
          5112 => x"14",
          5113 => x"82",
          5114 => x"52",
          5115 => x"ff",
          5116 => x"74",
          5117 => x"29",
          5118 => x"05",
          5119 => x"82",
          5120 => x"58",
          5121 => x"75",
          5122 => x"82",
          5123 => x"52",
          5124 => x"93",
          5125 => x"f7",
          5126 => x"98",
          5127 => x"2c",
          5128 => x"33",
          5129 => x"57",
          5130 => x"f8",
          5131 => x"fb",
          5132 => x"88",
          5133 => x"b0",
          5134 => x"80",
          5135 => x"80",
          5136 => x"98",
          5137 => x"d8",
          5138 => x"55",
          5139 => x"de",
          5140 => x"39",
          5141 => x"33",
          5142 => x"06",
          5143 => x"33",
          5144 => x"74",
          5145 => x"e6",
          5146 => x"fc",
          5147 => x"14",
          5148 => x"f7",
          5149 => x"1a",
          5150 => x"54",
          5151 => x"3f",
          5152 => x"33",
          5153 => x"06",
          5154 => x"33",
          5155 => x"75",
          5156 => x"38",
          5157 => x"82",
          5158 => x"80",
          5159 => x"b8",
          5160 => x"3f",
          5161 => x"f7",
          5162 => x"0b",
          5163 => x"34",
          5164 => x"7a",
          5165 => x"df",
          5166 => x"74",
          5167 => x"38",
          5168 => x"9a",
          5169 => x"e0",
          5170 => x"f7",
          5171 => x"e0",
          5172 => x"ff",
          5173 => x"53",
          5174 => x"51",
          5175 => x"3f",
          5176 => x"c0",
          5177 => x"29",
          5178 => x"05",
          5179 => x"56",
          5180 => x"2e",
          5181 => x"51",
          5182 => x"3f",
          5183 => x"08",
          5184 => x"34",
          5185 => x"08",
          5186 => x"81",
          5187 => x"52",
          5188 => x"9c",
          5189 => x"1b",
          5190 => x"39",
          5191 => x"74",
          5192 => x"aa",
          5193 => x"ff",
          5194 => x"99",
          5195 => x"2e",
          5196 => x"ae",
          5197 => x"90",
          5198 => x"80",
          5199 => x"74",
          5200 => x"f7",
          5201 => x"98",
          5202 => x"d8",
          5203 => x"98",
          5204 => x"06",
          5205 => x"74",
          5206 => x"ff",
          5207 => x"80",
          5208 => x"84",
          5209 => x"94",
          5210 => x"56",
          5211 => x"2e",
          5212 => x"51",
          5213 => x"3f",
          5214 => x"08",
          5215 => x"34",
          5216 => x"08",
          5217 => x"81",
          5218 => x"52",
          5219 => x"9b",
          5220 => x"1b",
          5221 => x"ff",
          5222 => x"39",
          5223 => x"d8",
          5224 => x"34",
          5225 => x"53",
          5226 => x"33",
          5227 => x"ec",
          5228 => x"9a",
          5229 => x"dc",
          5230 => x"ff",
          5231 => x"d8",
          5232 => x"54",
          5233 => x"f5",
          5234 => x"fb",
          5235 => x"81",
          5236 => x"82",
          5237 => x"74",
          5238 => x"52",
          5239 => x"88",
          5240 => x"39",
          5241 => x"33",
          5242 => x"2e",
          5243 => x"82",
          5244 => x"52",
          5245 => x"8f",
          5246 => x"f7",
          5247 => x"05",
          5248 => x"f7",
          5249 => x"c6",
          5250 => x"0d",
          5251 => x"0b",
          5252 => x"0c",
          5253 => x"82",
          5254 => x"82",
          5255 => x"80",
          5256 => x"f4",
          5257 => x"9f",
          5258 => x"88",
          5259 => x"58",
          5260 => x"81",
          5261 => x"15",
          5262 => x"88",
          5263 => x"84",
          5264 => x"85",
          5265 => x"e0",
          5266 => x"77",
          5267 => x"76",
          5268 => x"82",
          5269 => x"82",
          5270 => x"ff",
          5271 => x"80",
          5272 => x"ff",
          5273 => x"88",
          5274 => x"55",
          5275 => x"17",
          5276 => x"17",
          5277 => x"84",
          5278 => x"29",
          5279 => x"08",
          5280 => x"51",
          5281 => x"82",
          5282 => x"83",
          5283 => x"3d",
          5284 => x"3d",
          5285 => x"81",
          5286 => x"27",
          5287 => x"12",
          5288 => x"11",
          5289 => x"ff",
          5290 => x"51",
          5291 => x"98",
          5292 => x"0d",
          5293 => x"0d",
          5294 => x"22",
          5295 => x"aa",
          5296 => x"05",
          5297 => x"08",
          5298 => x"71",
          5299 => x"2b",
          5300 => x"33",
          5301 => x"71",
          5302 => x"02",
          5303 => x"05",
          5304 => x"ff",
          5305 => x"70",
          5306 => x"51",
          5307 => x"5b",
          5308 => x"54",
          5309 => x"34",
          5310 => x"34",
          5311 => x"08",
          5312 => x"2a",
          5313 => x"82",
          5314 => x"83",
          5315 => x"e0",
          5316 => x"17",
          5317 => x"12",
          5318 => x"2b",
          5319 => x"2b",
          5320 => x"06",
          5321 => x"52",
          5322 => x"83",
          5323 => x"70",
          5324 => x"54",
          5325 => x"12",
          5326 => x"ff",
          5327 => x"83",
          5328 => x"e0",
          5329 => x"56",
          5330 => x"72",
          5331 => x"89",
          5332 => x"fb",
          5333 => x"e0",
          5334 => x"84",
          5335 => x"22",
          5336 => x"72",
          5337 => x"33",
          5338 => x"71",
          5339 => x"83",
          5340 => x"5b",
          5341 => x"52",
          5342 => x"12",
          5343 => x"33",
          5344 => x"07",
          5345 => x"54",
          5346 => x"70",
          5347 => x"73",
          5348 => x"82",
          5349 => x"70",
          5350 => x"33",
          5351 => x"71",
          5352 => x"83",
          5353 => x"59",
          5354 => x"05",
          5355 => x"87",
          5356 => x"88",
          5357 => x"88",
          5358 => x"56",
          5359 => x"13",
          5360 => x"13",
          5361 => x"88",
          5362 => x"33",
          5363 => x"71",
          5364 => x"70",
          5365 => x"06",
          5366 => x"53",
          5367 => x"53",
          5368 => x"70",
          5369 => x"87",
          5370 => x"fa",
          5371 => x"a2",
          5372 => x"e0",
          5373 => x"83",
          5374 => x"70",
          5375 => x"33",
          5376 => x"07",
          5377 => x"15",
          5378 => x"12",
          5379 => x"2b",
          5380 => x"07",
          5381 => x"55",
          5382 => x"57",
          5383 => x"80",
          5384 => x"38",
          5385 => x"ab",
          5386 => x"88",
          5387 => x"70",
          5388 => x"33",
          5389 => x"71",
          5390 => x"74",
          5391 => x"81",
          5392 => x"88",
          5393 => x"83",
          5394 => x"f8",
          5395 => x"54",
          5396 => x"58",
          5397 => x"74",
          5398 => x"52",
          5399 => x"34",
          5400 => x"34",
          5401 => x"08",
          5402 => x"33",
          5403 => x"71",
          5404 => x"83",
          5405 => x"59",
          5406 => x"05",
          5407 => x"12",
          5408 => x"2b",
          5409 => x"ff",
          5410 => x"88",
          5411 => x"52",
          5412 => x"74",
          5413 => x"15",
          5414 => x"0d",
          5415 => x"0d",
          5416 => x"08",
          5417 => x"9e",
          5418 => x"83",
          5419 => x"82",
          5420 => x"12",
          5421 => x"2b",
          5422 => x"07",
          5423 => x"52",
          5424 => x"05",
          5425 => x"13",
          5426 => x"2b",
          5427 => x"05",
          5428 => x"71",
          5429 => x"2a",
          5430 => x"53",
          5431 => x"34",
          5432 => x"34",
          5433 => x"08",
          5434 => x"33",
          5435 => x"71",
          5436 => x"83",
          5437 => x"59",
          5438 => x"05",
          5439 => x"83",
          5440 => x"88",
          5441 => x"88",
          5442 => x"56",
          5443 => x"13",
          5444 => x"13",
          5445 => x"88",
          5446 => x"11",
          5447 => x"33",
          5448 => x"07",
          5449 => x"0c",
          5450 => x"3d",
          5451 => x"3d",
          5452 => x"e0",
          5453 => x"83",
          5454 => x"ff",
          5455 => x"53",
          5456 => x"a7",
          5457 => x"88",
          5458 => x"2b",
          5459 => x"11",
          5460 => x"33",
          5461 => x"71",
          5462 => x"75",
          5463 => x"81",
          5464 => x"98",
          5465 => x"2b",
          5466 => x"40",
          5467 => x"58",
          5468 => x"72",
          5469 => x"38",
          5470 => x"52",
          5471 => x"9d",
          5472 => x"39",
          5473 => x"85",
          5474 => x"8b",
          5475 => x"2b",
          5476 => x"79",
          5477 => x"51",
          5478 => x"76",
          5479 => x"75",
          5480 => x"56",
          5481 => x"34",
          5482 => x"08",
          5483 => x"12",
          5484 => x"33",
          5485 => x"07",
          5486 => x"54",
          5487 => x"53",
          5488 => x"34",
          5489 => x"34",
          5490 => x"08",
          5491 => x"0b",
          5492 => x"80",
          5493 => x"34",
          5494 => x"08",
          5495 => x"14",
          5496 => x"14",
          5497 => x"88",
          5498 => x"33",
          5499 => x"71",
          5500 => x"70",
          5501 => x"07",
          5502 => x"53",
          5503 => x"54",
          5504 => x"72",
          5505 => x"8b",
          5506 => x"ff",
          5507 => x"52",
          5508 => x"08",
          5509 => x"f1",
          5510 => x"2e",
          5511 => x"51",
          5512 => x"83",
          5513 => x"f5",
          5514 => x"7e",
          5515 => x"e2",
          5516 => x"98",
          5517 => x"ff",
          5518 => x"88",
          5519 => x"33",
          5520 => x"71",
          5521 => x"70",
          5522 => x"58",
          5523 => x"ff",
          5524 => x"2e",
          5525 => x"75",
          5526 => x"70",
          5527 => x"33",
          5528 => x"07",
          5529 => x"ff",
          5530 => x"70",
          5531 => x"06",
          5532 => x"52",
          5533 => x"59",
          5534 => x"27",
          5535 => x"80",
          5536 => x"75",
          5537 => x"84",
          5538 => x"16",
          5539 => x"2b",
          5540 => x"75",
          5541 => x"81",
          5542 => x"85",
          5543 => x"59",
          5544 => x"83",
          5545 => x"88",
          5546 => x"33",
          5547 => x"71",
          5548 => x"70",
          5549 => x"06",
          5550 => x"56",
          5551 => x"75",
          5552 => x"81",
          5553 => x"79",
          5554 => x"cc",
          5555 => x"74",
          5556 => x"c4",
          5557 => x"2e",
          5558 => x"89",
          5559 => x"f8",
          5560 => x"ac",
          5561 => x"80",
          5562 => x"75",
          5563 => x"3f",
          5564 => x"08",
          5565 => x"11",
          5566 => x"33",
          5567 => x"71",
          5568 => x"53",
          5569 => x"74",
          5570 => x"70",
          5571 => x"06",
          5572 => x"5c",
          5573 => x"78",
          5574 => x"76",
          5575 => x"57",
          5576 => x"34",
          5577 => x"08",
          5578 => x"71",
          5579 => x"86",
          5580 => x"12",
          5581 => x"2b",
          5582 => x"2a",
          5583 => x"53",
          5584 => x"73",
          5585 => x"75",
          5586 => x"82",
          5587 => x"70",
          5588 => x"33",
          5589 => x"71",
          5590 => x"83",
          5591 => x"5d",
          5592 => x"05",
          5593 => x"15",
          5594 => x"15",
          5595 => x"88",
          5596 => x"71",
          5597 => x"33",
          5598 => x"71",
          5599 => x"70",
          5600 => x"5a",
          5601 => x"54",
          5602 => x"34",
          5603 => x"34",
          5604 => x"08",
          5605 => x"54",
          5606 => x"98",
          5607 => x"0d",
          5608 => x"0d",
          5609 => x"e0",
          5610 => x"38",
          5611 => x"71",
          5612 => x"2e",
          5613 => x"51",
          5614 => x"82",
          5615 => x"53",
          5616 => x"98",
          5617 => x"0d",
          5618 => x"0d",
          5619 => x"5c",
          5620 => x"40",
          5621 => x"08",
          5622 => x"81",
          5623 => x"f4",
          5624 => x"8e",
          5625 => x"ff",
          5626 => x"e0",
          5627 => x"83",
          5628 => x"8b",
          5629 => x"fc",
          5630 => x"54",
          5631 => x"7e",
          5632 => x"3f",
          5633 => x"08",
          5634 => x"06",
          5635 => x"08",
          5636 => x"83",
          5637 => x"ff",
          5638 => x"83",
          5639 => x"70",
          5640 => x"33",
          5641 => x"07",
          5642 => x"70",
          5643 => x"06",
          5644 => x"fc",
          5645 => x"29",
          5646 => x"81",
          5647 => x"88",
          5648 => x"90",
          5649 => x"4e",
          5650 => x"52",
          5651 => x"41",
          5652 => x"5b",
          5653 => x"8f",
          5654 => x"ff",
          5655 => x"31",
          5656 => x"ff",
          5657 => x"82",
          5658 => x"17",
          5659 => x"2b",
          5660 => x"29",
          5661 => x"81",
          5662 => x"98",
          5663 => x"2b",
          5664 => x"45",
          5665 => x"73",
          5666 => x"38",
          5667 => x"70",
          5668 => x"06",
          5669 => x"7b",
          5670 => x"38",
          5671 => x"73",
          5672 => x"81",
          5673 => x"78",
          5674 => x"3f",
          5675 => x"ff",
          5676 => x"e5",
          5677 => x"38",
          5678 => x"89",
          5679 => x"f6",
          5680 => x"a5",
          5681 => x"55",
          5682 => x"80",
          5683 => x"1d",
          5684 => x"83",
          5685 => x"88",
          5686 => x"57",
          5687 => x"3f",
          5688 => x"51",
          5689 => x"82",
          5690 => x"83",
          5691 => x"7e",
          5692 => x"70",
          5693 => x"e0",
          5694 => x"84",
          5695 => x"59",
          5696 => x"3f",
          5697 => x"08",
          5698 => x"75",
          5699 => x"06",
          5700 => x"85",
          5701 => x"54",
          5702 => x"80",
          5703 => x"51",
          5704 => x"82",
          5705 => x"1d",
          5706 => x"83",
          5707 => x"88",
          5708 => x"43",
          5709 => x"3f",
          5710 => x"51",
          5711 => x"82",
          5712 => x"83",
          5713 => x"7e",
          5714 => x"70",
          5715 => x"e0",
          5716 => x"84",
          5717 => x"59",
          5718 => x"3f",
          5719 => x"08",
          5720 => x"60",
          5721 => x"55",
          5722 => x"ff",
          5723 => x"a9",
          5724 => x"52",
          5725 => x"3f",
          5726 => x"08",
          5727 => x"98",
          5728 => x"93",
          5729 => x"73",
          5730 => x"98",
          5731 => x"8b",
          5732 => x"51",
          5733 => x"7a",
          5734 => x"27",
          5735 => x"53",
          5736 => x"51",
          5737 => x"7a",
          5738 => x"82",
          5739 => x"05",
          5740 => x"f6",
          5741 => x"54",
          5742 => x"98",
          5743 => x"0d",
          5744 => x"0d",
          5745 => x"70",
          5746 => x"d5",
          5747 => x"98",
          5748 => x"e0",
          5749 => x"2e",
          5750 => x"53",
          5751 => x"e0",
          5752 => x"ff",
          5753 => x"74",
          5754 => x"0c",
          5755 => x"04",
          5756 => x"02",
          5757 => x"51",
          5758 => x"72",
          5759 => x"82",
          5760 => x"33",
          5761 => x"e0",
          5762 => x"3d",
          5763 => x"3d",
          5764 => x"05",
          5765 => x"05",
          5766 => x"56",
          5767 => x"72",
          5768 => x"e0",
          5769 => x"2b",
          5770 => x"8c",
          5771 => x"88",
          5772 => x"2e",
          5773 => x"88",
          5774 => x"0c",
          5775 => x"8c",
          5776 => x"71",
          5777 => x"87",
          5778 => x"0c",
          5779 => x"08",
          5780 => x"51",
          5781 => x"2e",
          5782 => x"c0",
          5783 => x"51",
          5784 => x"71",
          5785 => x"80",
          5786 => x"92",
          5787 => x"98",
          5788 => x"70",
          5789 => x"38",
          5790 => x"94",
          5791 => x"e0",
          5792 => x"51",
          5793 => x"98",
          5794 => x"0d",
          5795 => x"0d",
          5796 => x"02",
          5797 => x"05",
          5798 => x"58",
          5799 => x"52",
          5800 => x"3f",
          5801 => x"08",
          5802 => x"54",
          5803 => x"be",
          5804 => x"75",
          5805 => x"c0",
          5806 => x"87",
          5807 => x"12",
          5808 => x"84",
          5809 => x"40",
          5810 => x"85",
          5811 => x"98",
          5812 => x"7d",
          5813 => x"0c",
          5814 => x"85",
          5815 => x"06",
          5816 => x"71",
          5817 => x"38",
          5818 => x"71",
          5819 => x"05",
          5820 => x"19",
          5821 => x"a2",
          5822 => x"71",
          5823 => x"38",
          5824 => x"83",
          5825 => x"38",
          5826 => x"8a",
          5827 => x"98",
          5828 => x"71",
          5829 => x"c0",
          5830 => x"52",
          5831 => x"87",
          5832 => x"80",
          5833 => x"81",
          5834 => x"c0",
          5835 => x"53",
          5836 => x"82",
          5837 => x"71",
          5838 => x"1a",
          5839 => x"84",
          5840 => x"19",
          5841 => x"06",
          5842 => x"79",
          5843 => x"38",
          5844 => x"80",
          5845 => x"87",
          5846 => x"26",
          5847 => x"73",
          5848 => x"06",
          5849 => x"2e",
          5850 => x"52",
          5851 => x"82",
          5852 => x"8f",
          5853 => x"f3",
          5854 => x"62",
          5855 => x"05",
          5856 => x"57",
          5857 => x"83",
          5858 => x"52",
          5859 => x"3f",
          5860 => x"08",
          5861 => x"54",
          5862 => x"2e",
          5863 => x"81",
          5864 => x"74",
          5865 => x"c0",
          5866 => x"87",
          5867 => x"12",
          5868 => x"84",
          5869 => x"5f",
          5870 => x"0b",
          5871 => x"8c",
          5872 => x"0c",
          5873 => x"80",
          5874 => x"70",
          5875 => x"81",
          5876 => x"54",
          5877 => x"8c",
          5878 => x"81",
          5879 => x"7c",
          5880 => x"58",
          5881 => x"70",
          5882 => x"52",
          5883 => x"8a",
          5884 => x"98",
          5885 => x"71",
          5886 => x"c0",
          5887 => x"52",
          5888 => x"87",
          5889 => x"80",
          5890 => x"81",
          5891 => x"c0",
          5892 => x"53",
          5893 => x"82",
          5894 => x"71",
          5895 => x"19",
          5896 => x"81",
          5897 => x"ff",
          5898 => x"19",
          5899 => x"78",
          5900 => x"38",
          5901 => x"80",
          5902 => x"87",
          5903 => x"26",
          5904 => x"73",
          5905 => x"06",
          5906 => x"2e",
          5907 => x"52",
          5908 => x"82",
          5909 => x"8f",
          5910 => x"fa",
          5911 => x"02",
          5912 => x"05",
          5913 => x"05",
          5914 => x"71",
          5915 => x"57",
          5916 => x"82",
          5917 => x"81",
          5918 => x"54",
          5919 => x"38",
          5920 => x"c0",
          5921 => x"81",
          5922 => x"2e",
          5923 => x"71",
          5924 => x"38",
          5925 => x"87",
          5926 => x"11",
          5927 => x"80",
          5928 => x"80",
          5929 => x"83",
          5930 => x"38",
          5931 => x"72",
          5932 => x"2a",
          5933 => x"51",
          5934 => x"80",
          5935 => x"87",
          5936 => x"08",
          5937 => x"38",
          5938 => x"8c",
          5939 => x"96",
          5940 => x"0c",
          5941 => x"8c",
          5942 => x"08",
          5943 => x"51",
          5944 => x"38",
          5945 => x"56",
          5946 => x"80",
          5947 => x"85",
          5948 => x"77",
          5949 => x"83",
          5950 => x"75",
          5951 => x"e0",
          5952 => x"3d",
          5953 => x"3d",
          5954 => x"11",
          5955 => x"71",
          5956 => x"82",
          5957 => x"53",
          5958 => x"0d",
          5959 => x"0d",
          5960 => x"33",
          5961 => x"71",
          5962 => x"88",
          5963 => x"14",
          5964 => x"07",
          5965 => x"33",
          5966 => x"e0",
          5967 => x"53",
          5968 => x"52",
          5969 => x"04",
          5970 => x"73",
          5971 => x"92",
          5972 => x"52",
          5973 => x"81",
          5974 => x"70",
          5975 => x"70",
          5976 => x"3d",
          5977 => x"3d",
          5978 => x"52",
          5979 => x"70",
          5980 => x"34",
          5981 => x"51",
          5982 => x"81",
          5983 => x"70",
          5984 => x"70",
          5985 => x"05",
          5986 => x"88",
          5987 => x"72",
          5988 => x"0d",
          5989 => x"0d",
          5990 => x"54",
          5991 => x"80",
          5992 => x"71",
          5993 => x"53",
          5994 => x"81",
          5995 => x"ff",
          5996 => x"39",
          5997 => x"04",
          5998 => x"75",
          5999 => x"52",
          6000 => x"70",
          6001 => x"34",
          6002 => x"70",
          6003 => x"3d",
          6004 => x"3d",
          6005 => x"79",
          6006 => x"74",
          6007 => x"56",
          6008 => x"81",
          6009 => x"71",
          6010 => x"16",
          6011 => x"52",
          6012 => x"86",
          6013 => x"2e",
          6014 => x"82",
          6015 => x"86",
          6016 => x"fe",
          6017 => x"76",
          6018 => x"39",
          6019 => x"8a",
          6020 => x"51",
          6021 => x"71",
          6022 => x"33",
          6023 => x"0c",
          6024 => x"04",
          6025 => x"e0",
          6026 => x"fb",
          6027 => x"70",
          6028 => x"81",
          6029 => x"70",
          6030 => x"56",
          6031 => x"55",
          6032 => x"08",
          6033 => x"80",
          6034 => x"83",
          6035 => x"51",
          6036 => x"3f",
          6037 => x"08",
          6038 => x"06",
          6039 => x"2e",
          6040 => x"76",
          6041 => x"74",
          6042 => x"0c",
          6043 => x"04",
          6044 => x"7b",
          6045 => x"83",
          6046 => x"5a",
          6047 => x"80",
          6048 => x"54",
          6049 => x"53",
          6050 => x"53",
          6051 => x"52",
          6052 => x"3f",
          6053 => x"08",
          6054 => x"81",
          6055 => x"82",
          6056 => x"83",
          6057 => x"16",
          6058 => x"18",
          6059 => x"18",
          6060 => x"58",
          6061 => x"9f",
          6062 => x"33",
          6063 => x"2e",
          6064 => x"93",
          6065 => x"76",
          6066 => x"52",
          6067 => x"51",
          6068 => x"83",
          6069 => x"79",
          6070 => x"0c",
          6071 => x"04",
          6072 => x"78",
          6073 => x"80",
          6074 => x"17",
          6075 => x"38",
          6076 => x"fc",
          6077 => x"98",
          6078 => x"e0",
          6079 => x"38",
          6080 => x"53",
          6081 => x"81",
          6082 => x"f7",
          6083 => x"e0",
          6084 => x"2e",
          6085 => x"55",
          6086 => x"b4",
          6087 => x"82",
          6088 => x"88",
          6089 => x"f8",
          6090 => x"70",
          6091 => x"c0",
          6092 => x"98",
          6093 => x"e0",
          6094 => x"91",
          6095 => x"55",
          6096 => x"09",
          6097 => x"f0",
          6098 => x"33",
          6099 => x"2e",
          6100 => x"80",
          6101 => x"80",
          6102 => x"98",
          6103 => x"17",
          6104 => x"fc",
          6105 => x"d4",
          6106 => x"b6",
          6107 => x"d8",
          6108 => x"85",
          6109 => x"75",
          6110 => x"3f",
          6111 => x"e4",
          6112 => x"9c",
          6113 => x"de",
          6114 => x"08",
          6115 => x"17",
          6116 => x"3f",
          6117 => x"52",
          6118 => x"51",
          6119 => x"a4",
          6120 => x"05",
          6121 => x"0c",
          6122 => x"75",
          6123 => x"33",
          6124 => x"3f",
          6125 => x"34",
          6126 => x"52",
          6127 => x"51",
          6128 => x"82",
          6129 => x"80",
          6130 => x"81",
          6131 => x"e0",
          6132 => x"3d",
          6133 => x"3d",
          6134 => x"1a",
          6135 => x"fe",
          6136 => x"54",
          6137 => x"73",
          6138 => x"8a",
          6139 => x"71",
          6140 => x"08",
          6141 => x"75",
          6142 => x"0c",
          6143 => x"04",
          6144 => x"7a",
          6145 => x"56",
          6146 => x"77",
          6147 => x"38",
          6148 => x"08",
          6149 => x"38",
          6150 => x"54",
          6151 => x"2e",
          6152 => x"72",
          6153 => x"38",
          6154 => x"8d",
          6155 => x"39",
          6156 => x"81",
          6157 => x"b6",
          6158 => x"2a",
          6159 => x"2a",
          6160 => x"05",
          6161 => x"55",
          6162 => x"82",
          6163 => x"81",
          6164 => x"83",
          6165 => x"b8",
          6166 => x"17",
          6167 => x"a8",
          6168 => x"55",
          6169 => x"57",
          6170 => x"3f",
          6171 => x"08",
          6172 => x"74",
          6173 => x"14",
          6174 => x"70",
          6175 => x"07",
          6176 => x"71",
          6177 => x"52",
          6178 => x"72",
          6179 => x"75",
          6180 => x"58",
          6181 => x"76",
          6182 => x"15",
          6183 => x"73",
          6184 => x"3f",
          6185 => x"08",
          6186 => x"76",
          6187 => x"06",
          6188 => x"05",
          6189 => x"3f",
          6190 => x"08",
          6191 => x"06",
          6192 => x"76",
          6193 => x"15",
          6194 => x"73",
          6195 => x"3f",
          6196 => x"08",
          6197 => x"82",
          6198 => x"06",
          6199 => x"05",
          6200 => x"3f",
          6201 => x"08",
          6202 => x"58",
          6203 => x"58",
          6204 => x"98",
          6205 => x"0d",
          6206 => x"0d",
          6207 => x"5a",
          6208 => x"59",
          6209 => x"82",
          6210 => x"9c",
          6211 => x"82",
          6212 => x"33",
          6213 => x"2e",
          6214 => x"72",
          6215 => x"38",
          6216 => x"8d",
          6217 => x"39",
          6218 => x"81",
          6219 => x"f7",
          6220 => x"2a",
          6221 => x"2a",
          6222 => x"05",
          6223 => x"55",
          6224 => x"82",
          6225 => x"59",
          6226 => x"08",
          6227 => x"74",
          6228 => x"16",
          6229 => x"16",
          6230 => x"59",
          6231 => x"53",
          6232 => x"8f",
          6233 => x"2b",
          6234 => x"74",
          6235 => x"71",
          6236 => x"72",
          6237 => x"0b",
          6238 => x"74",
          6239 => x"17",
          6240 => x"75",
          6241 => x"3f",
          6242 => x"08",
          6243 => x"98",
          6244 => x"38",
          6245 => x"06",
          6246 => x"78",
          6247 => x"54",
          6248 => x"77",
          6249 => x"33",
          6250 => x"71",
          6251 => x"51",
          6252 => x"34",
          6253 => x"76",
          6254 => x"17",
          6255 => x"75",
          6256 => x"3f",
          6257 => x"08",
          6258 => x"98",
          6259 => x"38",
          6260 => x"ff",
          6261 => x"10",
          6262 => x"76",
          6263 => x"51",
          6264 => x"be",
          6265 => x"2a",
          6266 => x"05",
          6267 => x"f9",
          6268 => x"e0",
          6269 => x"82",
          6270 => x"ab",
          6271 => x"0a",
          6272 => x"2b",
          6273 => x"70",
          6274 => x"70",
          6275 => x"54",
          6276 => x"82",
          6277 => x"8f",
          6278 => x"07",
          6279 => x"f6",
          6280 => x"0b",
          6281 => x"78",
          6282 => x"0c",
          6283 => x"04",
          6284 => x"7a",
          6285 => x"08",
          6286 => x"59",
          6287 => x"a4",
          6288 => x"17",
          6289 => x"38",
          6290 => x"aa",
          6291 => x"73",
          6292 => x"fd",
          6293 => x"e0",
          6294 => x"82",
          6295 => x"80",
          6296 => x"39",
          6297 => x"eb",
          6298 => x"80",
          6299 => x"e0",
          6300 => x"80",
          6301 => x"52",
          6302 => x"84",
          6303 => x"98",
          6304 => x"e0",
          6305 => x"2e",
          6306 => x"82",
          6307 => x"81",
          6308 => x"82",
          6309 => x"ff",
          6310 => x"80",
          6311 => x"75",
          6312 => x"3f",
          6313 => x"08",
          6314 => x"16",
          6315 => x"94",
          6316 => x"55",
          6317 => x"27",
          6318 => x"15",
          6319 => x"84",
          6320 => x"07",
          6321 => x"17",
          6322 => x"76",
          6323 => x"a6",
          6324 => x"73",
          6325 => x"0c",
          6326 => x"04",
          6327 => x"7c",
          6328 => x"59",
          6329 => x"95",
          6330 => x"08",
          6331 => x"2e",
          6332 => x"17",
          6333 => x"b2",
          6334 => x"ae",
          6335 => x"7a",
          6336 => x"3f",
          6337 => x"82",
          6338 => x"27",
          6339 => x"82",
          6340 => x"55",
          6341 => x"08",
          6342 => x"d2",
          6343 => x"08",
          6344 => x"08",
          6345 => x"38",
          6346 => x"17",
          6347 => x"54",
          6348 => x"82",
          6349 => x"7a",
          6350 => x"06",
          6351 => x"81",
          6352 => x"17",
          6353 => x"83",
          6354 => x"75",
          6355 => x"f9",
          6356 => x"59",
          6357 => x"08",
          6358 => x"81",
          6359 => x"82",
          6360 => x"59",
          6361 => x"08",
          6362 => x"70",
          6363 => x"25",
          6364 => x"82",
          6365 => x"54",
          6366 => x"55",
          6367 => x"38",
          6368 => x"08",
          6369 => x"38",
          6370 => x"54",
          6371 => x"90",
          6372 => x"18",
          6373 => x"38",
          6374 => x"39",
          6375 => x"38",
          6376 => x"16",
          6377 => x"08",
          6378 => x"38",
          6379 => x"78",
          6380 => x"38",
          6381 => x"51",
          6382 => x"82",
          6383 => x"80",
          6384 => x"80",
          6385 => x"98",
          6386 => x"09",
          6387 => x"38",
          6388 => x"08",
          6389 => x"98",
          6390 => x"30",
          6391 => x"80",
          6392 => x"07",
          6393 => x"55",
          6394 => x"38",
          6395 => x"09",
          6396 => x"ae",
          6397 => x"80",
          6398 => x"53",
          6399 => x"51",
          6400 => x"82",
          6401 => x"82",
          6402 => x"30",
          6403 => x"98",
          6404 => x"25",
          6405 => x"79",
          6406 => x"38",
          6407 => x"8f",
          6408 => x"79",
          6409 => x"f9",
          6410 => x"e0",
          6411 => x"74",
          6412 => x"90",
          6413 => x"17",
          6414 => x"94",
          6415 => x"54",
          6416 => x"86",
          6417 => x"94",
          6418 => x"17",
          6419 => x"54",
          6420 => x"34",
          6421 => x"56",
          6422 => x"90",
          6423 => x"80",
          6424 => x"82",
          6425 => x"55",
          6426 => x"56",
          6427 => x"82",
          6428 => x"8c",
          6429 => x"f8",
          6430 => x"70",
          6431 => x"f0",
          6432 => x"98",
          6433 => x"56",
          6434 => x"08",
          6435 => x"7b",
          6436 => x"f6",
          6437 => x"e0",
          6438 => x"e0",
          6439 => x"17",
          6440 => x"80",
          6441 => x"b8",
          6442 => x"57",
          6443 => x"77",
          6444 => x"81",
          6445 => x"15",
          6446 => x"78",
          6447 => x"81",
          6448 => x"53",
          6449 => x"15",
          6450 => x"ab",
          6451 => x"98",
          6452 => x"df",
          6453 => x"22",
          6454 => x"30",
          6455 => x"70",
          6456 => x"51",
          6457 => x"82",
          6458 => x"8a",
          6459 => x"f8",
          6460 => x"7c",
          6461 => x"56",
          6462 => x"80",
          6463 => x"f1",
          6464 => x"06",
          6465 => x"e9",
          6466 => x"18",
          6467 => x"08",
          6468 => x"38",
          6469 => x"82",
          6470 => x"38",
          6471 => x"54",
          6472 => x"74",
          6473 => x"82",
          6474 => x"22",
          6475 => x"79",
          6476 => x"38",
          6477 => x"98",
          6478 => x"cd",
          6479 => x"22",
          6480 => x"54",
          6481 => x"26",
          6482 => x"52",
          6483 => x"b0",
          6484 => x"98",
          6485 => x"e0",
          6486 => x"2e",
          6487 => x"0b",
          6488 => x"08",
          6489 => x"9c",
          6490 => x"e0",
          6491 => x"85",
          6492 => x"bd",
          6493 => x"31",
          6494 => x"73",
          6495 => x"f4",
          6496 => x"e0",
          6497 => x"18",
          6498 => x"18",
          6499 => x"08",
          6500 => x"72",
          6501 => x"38",
          6502 => x"58",
          6503 => x"89",
          6504 => x"18",
          6505 => x"ff",
          6506 => x"05",
          6507 => x"80",
          6508 => x"e0",
          6509 => x"3d",
          6510 => x"3d",
          6511 => x"08",
          6512 => x"a0",
          6513 => x"54",
          6514 => x"77",
          6515 => x"80",
          6516 => x"0c",
          6517 => x"53",
          6518 => x"80",
          6519 => x"38",
          6520 => x"06",
          6521 => x"b5",
          6522 => x"98",
          6523 => x"14",
          6524 => x"92",
          6525 => x"2a",
          6526 => x"56",
          6527 => x"26",
          6528 => x"80",
          6529 => x"16",
          6530 => x"77",
          6531 => x"53",
          6532 => x"38",
          6533 => x"51",
          6534 => x"82",
          6535 => x"53",
          6536 => x"0b",
          6537 => x"08",
          6538 => x"38",
          6539 => x"e0",
          6540 => x"2e",
          6541 => x"9c",
          6542 => x"e0",
          6543 => x"80",
          6544 => x"8a",
          6545 => x"15",
          6546 => x"80",
          6547 => x"14",
          6548 => x"51",
          6549 => x"82",
          6550 => x"53",
          6551 => x"e0",
          6552 => x"2e",
          6553 => x"82",
          6554 => x"98",
          6555 => x"ba",
          6556 => x"82",
          6557 => x"ff",
          6558 => x"82",
          6559 => x"52",
          6560 => x"f3",
          6561 => x"98",
          6562 => x"72",
          6563 => x"72",
          6564 => x"f2",
          6565 => x"e0",
          6566 => x"15",
          6567 => x"15",
          6568 => x"b8",
          6569 => x"0c",
          6570 => x"82",
          6571 => x"8a",
          6572 => x"f7",
          6573 => x"7d",
          6574 => x"5b",
          6575 => x"76",
          6576 => x"3f",
          6577 => x"08",
          6578 => x"98",
          6579 => x"38",
          6580 => x"08",
          6581 => x"08",
          6582 => x"f0",
          6583 => x"e0",
          6584 => x"82",
          6585 => x"80",
          6586 => x"e0",
          6587 => x"18",
          6588 => x"51",
          6589 => x"81",
          6590 => x"81",
          6591 => x"81",
          6592 => x"98",
          6593 => x"83",
          6594 => x"77",
          6595 => x"72",
          6596 => x"38",
          6597 => x"75",
          6598 => x"81",
          6599 => x"a5",
          6600 => x"98",
          6601 => x"52",
          6602 => x"8e",
          6603 => x"98",
          6604 => x"e0",
          6605 => x"2e",
          6606 => x"73",
          6607 => x"81",
          6608 => x"87",
          6609 => x"e0",
          6610 => x"3d",
          6611 => x"3d",
          6612 => x"11",
          6613 => x"ae",
          6614 => x"98",
          6615 => x"ff",
          6616 => x"33",
          6617 => x"71",
          6618 => x"81",
          6619 => x"94",
          6620 => x"92",
          6621 => x"98",
          6622 => x"73",
          6623 => x"82",
          6624 => x"85",
          6625 => x"fc",
          6626 => x"79",
          6627 => x"ff",
          6628 => x"12",
          6629 => x"eb",
          6630 => x"70",
          6631 => x"72",
          6632 => x"81",
          6633 => x"73",
          6634 => x"94",
          6635 => x"98",
          6636 => x"0d",
          6637 => x"0d",
          6638 => x"51",
          6639 => x"81",
          6640 => x"80",
          6641 => x"70",
          6642 => x"33",
          6643 => x"81",
          6644 => x"16",
          6645 => x"51",
          6646 => x"70",
          6647 => x"0c",
          6648 => x"04",
          6649 => x"60",
          6650 => x"84",
          6651 => x"5b",
          6652 => x"5d",
          6653 => x"08",
          6654 => x"80",
          6655 => x"08",
          6656 => x"ed",
          6657 => x"e0",
          6658 => x"82",
          6659 => x"82",
          6660 => x"19",
          6661 => x"55",
          6662 => x"38",
          6663 => x"dc",
          6664 => x"33",
          6665 => x"81",
          6666 => x"53",
          6667 => x"34",
          6668 => x"08",
          6669 => x"e5",
          6670 => x"06",
          6671 => x"56",
          6672 => x"08",
          6673 => x"2e",
          6674 => x"83",
          6675 => x"75",
          6676 => x"72",
          6677 => x"e0",
          6678 => x"df",
          6679 => x"72",
          6680 => x"81",
          6681 => x"81",
          6682 => x"2e",
          6683 => x"ff",
          6684 => x"39",
          6685 => x"09",
          6686 => x"ca",
          6687 => x"2a",
          6688 => x"51",
          6689 => x"2e",
          6690 => x"15",
          6691 => x"bf",
          6692 => x"1c",
          6693 => x"0c",
          6694 => x"73",
          6695 => x"81",
          6696 => x"38",
          6697 => x"53",
          6698 => x"09",
          6699 => x"8f",
          6700 => x"08",
          6701 => x"5a",
          6702 => x"82",
          6703 => x"83",
          6704 => x"53",
          6705 => x"38",
          6706 => x"81",
          6707 => x"29",
          6708 => x"54",
          6709 => x"58",
          6710 => x"17",
          6711 => x"51",
          6712 => x"82",
          6713 => x"83",
          6714 => x"56",
          6715 => x"96",
          6716 => x"fe",
          6717 => x"38",
          6718 => x"76",
          6719 => x"73",
          6720 => x"54",
          6721 => x"83",
          6722 => x"09",
          6723 => x"38",
          6724 => x"8c",
          6725 => x"38",
          6726 => x"86",
          6727 => x"06",
          6728 => x"72",
          6729 => x"38",
          6730 => x"26",
          6731 => x"10",
          6732 => x"73",
          6733 => x"70",
          6734 => x"51",
          6735 => x"81",
          6736 => x"5c",
          6737 => x"93",
          6738 => x"fc",
          6739 => x"e0",
          6740 => x"ff",
          6741 => x"7d",
          6742 => x"ff",
          6743 => x"0c",
          6744 => x"52",
          6745 => x"d2",
          6746 => x"98",
          6747 => x"e0",
          6748 => x"38",
          6749 => x"fd",
          6750 => x"39",
          6751 => x"1a",
          6752 => x"e0",
          6753 => x"3d",
          6754 => x"3d",
          6755 => x"08",
          6756 => x"52",
          6757 => x"d7",
          6758 => x"98",
          6759 => x"e0",
          6760 => x"a4",
          6761 => x"70",
          6762 => x"0b",
          6763 => x"98",
          6764 => x"7e",
          6765 => x"3f",
          6766 => x"08",
          6767 => x"98",
          6768 => x"38",
          6769 => x"70",
          6770 => x"75",
          6771 => x"58",
          6772 => x"8b",
          6773 => x"06",
          6774 => x"06",
          6775 => x"86",
          6776 => x"81",
          6777 => x"c3",
          6778 => x"2a",
          6779 => x"51",
          6780 => x"2e",
          6781 => x"82",
          6782 => x"8f",
          6783 => x"06",
          6784 => x"ab",
          6785 => x"86",
          6786 => x"06",
          6787 => x"73",
          6788 => x"75",
          6789 => x"81",
          6790 => x"73",
          6791 => x"38",
          6792 => x"76",
          6793 => x"70",
          6794 => x"ac",
          6795 => x"5d",
          6796 => x"2e",
          6797 => x"81",
          6798 => x"17",
          6799 => x"76",
          6800 => x"06",
          6801 => x"8c",
          6802 => x"18",
          6803 => x"b6",
          6804 => x"98",
          6805 => x"ff",
          6806 => x"81",
          6807 => x"33",
          6808 => x"8d",
          6809 => x"59",
          6810 => x"5c",
          6811 => x"a8",
          6812 => x"05",
          6813 => x"3f",
          6814 => x"08",
          6815 => x"06",
          6816 => x"2e",
          6817 => x"81",
          6818 => x"e6",
          6819 => x"80",
          6820 => x"82",
          6821 => x"78",
          6822 => x"22",
          6823 => x"19",
          6824 => x"e1",
          6825 => x"82",
          6826 => x"2e",
          6827 => x"80",
          6828 => x"5a",
          6829 => x"83",
          6830 => x"09",
          6831 => x"38",
          6832 => x"8c",
          6833 => x"a5",
          6834 => x"70",
          6835 => x"81",
          6836 => x"57",
          6837 => x"90",
          6838 => x"2e",
          6839 => x"10",
          6840 => x"51",
          6841 => x"38",
          6842 => x"81",
          6843 => x"54",
          6844 => x"ff",
          6845 => x"bb",
          6846 => x"38",
          6847 => x"b5",
          6848 => x"98",
          6849 => x"06",
          6850 => x"2e",
          6851 => x"19",
          6852 => x"54",
          6853 => x"8b",
          6854 => x"52",
          6855 => x"51",
          6856 => x"82",
          6857 => x"80",
          6858 => x"81",
          6859 => x"0b",
          6860 => x"80",
          6861 => x"f5",
          6862 => x"e0",
          6863 => x"82",
          6864 => x"80",
          6865 => x"38",
          6866 => x"98",
          6867 => x"0d",
          6868 => x"0d",
          6869 => x"ab",
          6870 => x"a0",
          6871 => x"5a",
          6872 => x"85",
          6873 => x"8c",
          6874 => x"22",
          6875 => x"73",
          6876 => x"38",
          6877 => x"10",
          6878 => x"51",
          6879 => x"39",
          6880 => x"1a",
          6881 => x"3d",
          6882 => x"59",
          6883 => x"02",
          6884 => x"33",
          6885 => x"73",
          6886 => x"a8",
          6887 => x"0b",
          6888 => x"81",
          6889 => x"08",
          6890 => x"8b",
          6891 => x"78",
          6892 => x"3f",
          6893 => x"80",
          6894 => x"56",
          6895 => x"83",
          6896 => x"55",
          6897 => x"2e",
          6898 => x"83",
          6899 => x"82",
          6900 => x"8f",
          6901 => x"06",
          6902 => x"75",
          6903 => x"90",
          6904 => x"06",
          6905 => x"56",
          6906 => x"87",
          6907 => x"a0",
          6908 => x"ff",
          6909 => x"80",
          6910 => x"c0",
          6911 => x"87",
          6912 => x"bf",
          6913 => x"74",
          6914 => x"06",
          6915 => x"27",
          6916 => x"14",
          6917 => x"34",
          6918 => x"18",
          6919 => x"57",
          6920 => x"e3",
          6921 => x"ec",
          6922 => x"80",
          6923 => x"80",
          6924 => x"38",
          6925 => x"73",
          6926 => x"38",
          6927 => x"33",
          6928 => x"e0",
          6929 => x"98",
          6930 => x"8c",
          6931 => x"54",
          6932 => x"94",
          6933 => x"55",
          6934 => x"74",
          6935 => x"38",
          6936 => x"33",
          6937 => x"39",
          6938 => x"05",
          6939 => x"78",
          6940 => x"56",
          6941 => x"76",
          6942 => x"38",
          6943 => x"15",
          6944 => x"55",
          6945 => x"34",
          6946 => x"e3",
          6947 => x"f9",
          6948 => x"e0",
          6949 => x"38",
          6950 => x"80",
          6951 => x"fe",
          6952 => x"55",
          6953 => x"2e",
          6954 => x"82",
          6955 => x"55",
          6956 => x"08",
          6957 => x"81",
          6958 => x"38",
          6959 => x"05",
          6960 => x"34",
          6961 => x"05",
          6962 => x"2a",
          6963 => x"51",
          6964 => x"59",
          6965 => x"90",
          6966 => x"8c",
          6967 => x"eb",
          6968 => x"e0",
          6969 => x"59",
          6970 => x"51",
          6971 => x"82",
          6972 => x"57",
          6973 => x"08",
          6974 => x"ff",
          6975 => x"80",
          6976 => x"38",
          6977 => x"90",
          6978 => x"31",
          6979 => x"51",
          6980 => x"82",
          6981 => x"57",
          6982 => x"08",
          6983 => x"a0",
          6984 => x"91",
          6985 => x"98",
          6986 => x"06",
          6987 => x"08",
          6988 => x"e3",
          6989 => x"e0",
          6990 => x"82",
          6991 => x"81",
          6992 => x"1c",
          6993 => x"08",
          6994 => x"06",
          6995 => x"7c",
          6996 => x"8f",
          6997 => x"34",
          6998 => x"08",
          6999 => x"82",
          7000 => x"52",
          7001 => x"df",
          7002 => x"8d",
          7003 => x"77",
          7004 => x"83",
          7005 => x"8b",
          7006 => x"1b",
          7007 => x"17",
          7008 => x"73",
          7009 => x"a8",
          7010 => x"05",
          7011 => x"3f",
          7012 => x"83",
          7013 => x"81",
          7014 => x"77",
          7015 => x"73",
          7016 => x"2e",
          7017 => x"10",
          7018 => x"51",
          7019 => x"38",
          7020 => x"07",
          7021 => x"34",
          7022 => x"1d",
          7023 => x"79",
          7024 => x"3f",
          7025 => x"08",
          7026 => x"98",
          7027 => x"38",
          7028 => x"78",
          7029 => x"98",
          7030 => x"7b",
          7031 => x"3f",
          7032 => x"08",
          7033 => x"98",
          7034 => x"a0",
          7035 => x"98",
          7036 => x"1a",
          7037 => x"c0",
          7038 => x"a0",
          7039 => x"1a",
          7040 => x"91",
          7041 => x"08",
          7042 => x"98",
          7043 => x"73",
          7044 => x"81",
          7045 => x"34",
          7046 => x"82",
          7047 => x"94",
          7048 => x"fa",
          7049 => x"70",
          7050 => x"08",
          7051 => x"56",
          7052 => x"72",
          7053 => x"38",
          7054 => x"51",
          7055 => x"82",
          7056 => x"54",
          7057 => x"08",
          7058 => x"98",
          7059 => x"75",
          7060 => x"3f",
          7061 => x"08",
          7062 => x"98",
          7063 => x"9c",
          7064 => x"e5",
          7065 => x"0b",
          7066 => x"90",
          7067 => x"27",
          7068 => x"e0",
          7069 => x"74",
          7070 => x"3f",
          7071 => x"08",
          7072 => x"98",
          7073 => x"c3",
          7074 => x"2e",
          7075 => x"83",
          7076 => x"73",
          7077 => x"0c",
          7078 => x"04",
          7079 => x"7e",
          7080 => x"5f",
          7081 => x"0b",
          7082 => x"98",
          7083 => x"2e",
          7084 => x"ac",
          7085 => x"2e",
          7086 => x"80",
          7087 => x"8c",
          7088 => x"22",
          7089 => x"5c",
          7090 => x"2e",
          7091 => x"78",
          7092 => x"22",
          7093 => x"56",
          7094 => x"38",
          7095 => x"15",
          7096 => x"ff",
          7097 => x"72",
          7098 => x"86",
          7099 => x"80",
          7100 => x"18",
          7101 => x"ff",
          7102 => x"5b",
          7103 => x"52",
          7104 => x"75",
          7105 => x"d7",
          7106 => x"e0",
          7107 => x"ff",
          7108 => x"81",
          7109 => x"95",
          7110 => x"27",
          7111 => x"88",
          7112 => x"7a",
          7113 => x"15",
          7114 => x"9f",
          7115 => x"76",
          7116 => x"07",
          7117 => x"80",
          7118 => x"54",
          7119 => x"2e",
          7120 => x"57",
          7121 => x"7a",
          7122 => x"74",
          7123 => x"5b",
          7124 => x"79",
          7125 => x"22",
          7126 => x"72",
          7127 => x"7a",
          7128 => x"25",
          7129 => x"06",
          7130 => x"77",
          7131 => x"53",
          7132 => x"14",
          7133 => x"89",
          7134 => x"57",
          7135 => x"19",
          7136 => x"1b",
          7137 => x"74",
          7138 => x"38",
          7139 => x"09",
          7140 => x"38",
          7141 => x"78",
          7142 => x"30",
          7143 => x"80",
          7144 => x"54",
          7145 => x"90",
          7146 => x"2e",
          7147 => x"76",
          7148 => x"58",
          7149 => x"57",
          7150 => x"81",
          7151 => x"81",
          7152 => x"79",
          7153 => x"38",
          7154 => x"05",
          7155 => x"81",
          7156 => x"18",
          7157 => x"81",
          7158 => x"8b",
          7159 => x"96",
          7160 => x"57",
          7161 => x"72",
          7162 => x"33",
          7163 => x"72",
          7164 => x"d3",
          7165 => x"89",
          7166 => x"73",
          7167 => x"11",
          7168 => x"99",
          7169 => x"9c",
          7170 => x"11",
          7171 => x"88",
          7172 => x"38",
          7173 => x"53",
          7174 => x"83",
          7175 => x"81",
          7176 => x"80",
          7177 => x"a0",
          7178 => x"ff",
          7179 => x"53",
          7180 => x"81",
          7181 => x"81",
          7182 => x"81",
          7183 => x"56",
          7184 => x"72",
          7185 => x"77",
          7186 => x"53",
          7187 => x"14",
          7188 => x"08",
          7189 => x"51",
          7190 => x"38",
          7191 => x"34",
          7192 => x"53",
          7193 => x"88",
          7194 => x"1c",
          7195 => x"52",
          7196 => x"3f",
          7197 => x"08",
          7198 => x"13",
          7199 => x"3f",
          7200 => x"08",
          7201 => x"98",
          7202 => x"fa",
          7203 => x"98",
          7204 => x"23",
          7205 => x"04",
          7206 => x"62",
          7207 => x"5e",
          7208 => x"33",
          7209 => x"73",
          7210 => x"38",
          7211 => x"80",
          7212 => x"38",
          7213 => x"8d",
          7214 => x"05",
          7215 => x"0c",
          7216 => x"15",
          7217 => x"70",
          7218 => x"56",
          7219 => x"09",
          7220 => x"38",
          7221 => x"80",
          7222 => x"30",
          7223 => x"78",
          7224 => x"54",
          7225 => x"73",
          7226 => x"63",
          7227 => x"54",
          7228 => x"96",
          7229 => x"0b",
          7230 => x"80",
          7231 => x"e7",
          7232 => x"e0",
          7233 => x"87",
          7234 => x"41",
          7235 => x"11",
          7236 => x"80",
          7237 => x"fc",
          7238 => x"8f",
          7239 => x"98",
          7240 => x"82",
          7241 => x"ff",
          7242 => x"e0",
          7243 => x"92",
          7244 => x"1a",
          7245 => x"08",
          7246 => x"55",
          7247 => x"81",
          7248 => x"e0",
          7249 => x"ff",
          7250 => x"af",
          7251 => x"9f",
          7252 => x"80",
          7253 => x"51",
          7254 => x"b4",
          7255 => x"dc",
          7256 => x"75",
          7257 => x"91",
          7258 => x"82",
          7259 => x"d9",
          7260 => x"e0",
          7261 => x"de",
          7262 => x"fe",
          7263 => x"38",
          7264 => x"54",
          7265 => x"81",
          7266 => x"89",
          7267 => x"41",
          7268 => x"33",
          7269 => x"73",
          7270 => x"81",
          7271 => x"81",
          7272 => x"dc",
          7273 => x"70",
          7274 => x"07",
          7275 => x"73",
          7276 => x"44",
          7277 => x"82",
          7278 => x"81",
          7279 => x"06",
          7280 => x"22",
          7281 => x"2e",
          7282 => x"d2",
          7283 => x"2e",
          7284 => x"80",
          7285 => x"1a",
          7286 => x"ae",
          7287 => x"06",
          7288 => x"79",
          7289 => x"ae",
          7290 => x"06",
          7291 => x"10",
          7292 => x"74",
          7293 => x"a0",
          7294 => x"ae",
          7295 => x"26",
          7296 => x"54",
          7297 => x"81",
          7298 => x"81",
          7299 => x"78",
          7300 => x"76",
          7301 => x"73",
          7302 => x"84",
          7303 => x"80",
          7304 => x"78",
          7305 => x"05",
          7306 => x"fe",
          7307 => x"a0",
          7308 => x"70",
          7309 => x"51",
          7310 => x"54",
          7311 => x"84",
          7312 => x"38",
          7313 => x"78",
          7314 => x"19",
          7315 => x"56",
          7316 => x"78",
          7317 => x"56",
          7318 => x"76",
          7319 => x"83",
          7320 => x"7a",
          7321 => x"ff",
          7322 => x"56",
          7323 => x"2e",
          7324 => x"93",
          7325 => x"70",
          7326 => x"22",
          7327 => x"73",
          7328 => x"38",
          7329 => x"74",
          7330 => x"06",
          7331 => x"2e",
          7332 => x"85",
          7333 => x"07",
          7334 => x"2e",
          7335 => x"16",
          7336 => x"22",
          7337 => x"ae",
          7338 => x"78",
          7339 => x"05",
          7340 => x"59",
          7341 => x"8f",
          7342 => x"70",
          7343 => x"73",
          7344 => x"81",
          7345 => x"8b",
          7346 => x"a0",
          7347 => x"e8",
          7348 => x"59",
          7349 => x"7c",
          7350 => x"22",
          7351 => x"57",
          7352 => x"2e",
          7353 => x"75",
          7354 => x"38",
          7355 => x"70",
          7356 => x"25",
          7357 => x"7c",
          7358 => x"38",
          7359 => x"89",
          7360 => x"07",
          7361 => x"80",
          7362 => x"7e",
          7363 => x"38",
          7364 => x"79",
          7365 => x"70",
          7366 => x"25",
          7367 => x"51",
          7368 => x"73",
          7369 => x"38",
          7370 => x"fe",
          7371 => x"79",
          7372 => x"76",
          7373 => x"7c",
          7374 => x"be",
          7375 => x"88",
          7376 => x"82",
          7377 => x"06",
          7378 => x"8b",
          7379 => x"76",
          7380 => x"76",
          7381 => x"83",
          7382 => x"51",
          7383 => x"3f",
          7384 => x"08",
          7385 => x"06",
          7386 => x"70",
          7387 => x"55",
          7388 => x"2e",
          7389 => x"80",
          7390 => x"d2",
          7391 => x"57",
          7392 => x"76",
          7393 => x"ff",
          7394 => x"78",
          7395 => x"76",
          7396 => x"59",
          7397 => x"39",
          7398 => x"05",
          7399 => x"55",
          7400 => x"34",
          7401 => x"80",
          7402 => x"80",
          7403 => x"75",
          7404 => x"d0",
          7405 => x"3f",
          7406 => x"08",
          7407 => x"38",
          7408 => x"83",
          7409 => x"a4",
          7410 => x"16",
          7411 => x"26",
          7412 => x"82",
          7413 => x"9f",
          7414 => x"99",
          7415 => x"7b",
          7416 => x"17",
          7417 => x"ff",
          7418 => x"5c",
          7419 => x"05",
          7420 => x"34",
          7421 => x"fd",
          7422 => x"1e",
          7423 => x"81",
          7424 => x"81",
          7425 => x"85",
          7426 => x"34",
          7427 => x"09",
          7428 => x"38",
          7429 => x"81",
          7430 => x"7b",
          7431 => x"73",
          7432 => x"38",
          7433 => x"54",
          7434 => x"09",
          7435 => x"38",
          7436 => x"57",
          7437 => x"70",
          7438 => x"54",
          7439 => x"7b",
          7440 => x"73",
          7441 => x"38",
          7442 => x"57",
          7443 => x"70",
          7444 => x"54",
          7445 => x"85",
          7446 => x"07",
          7447 => x"1f",
          7448 => x"ea",
          7449 => x"e0",
          7450 => x"1f",
          7451 => x"82",
          7452 => x"80",
          7453 => x"82",
          7454 => x"84",
          7455 => x"06",
          7456 => x"74",
          7457 => x"81",
          7458 => x"2a",
          7459 => x"73",
          7460 => x"38",
          7461 => x"54",
          7462 => x"f8",
          7463 => x"80",
          7464 => x"34",
          7465 => x"c2",
          7466 => x"06",
          7467 => x"38",
          7468 => x"39",
          7469 => x"70",
          7470 => x"54",
          7471 => x"86",
          7472 => x"84",
          7473 => x"06",
          7474 => x"73",
          7475 => x"38",
          7476 => x"83",
          7477 => x"05",
          7478 => x"7f",
          7479 => x"3f",
          7480 => x"08",
          7481 => x"f8",
          7482 => x"82",
          7483 => x"92",
          7484 => x"f6",
          7485 => x"5b",
          7486 => x"70",
          7487 => x"59",
          7488 => x"73",
          7489 => x"c6",
          7490 => x"81",
          7491 => x"70",
          7492 => x"52",
          7493 => x"8d",
          7494 => x"38",
          7495 => x"09",
          7496 => x"a5",
          7497 => x"d0",
          7498 => x"ff",
          7499 => x"53",
          7500 => x"91",
          7501 => x"73",
          7502 => x"d0",
          7503 => x"71",
          7504 => x"f7",
          7505 => x"82",
          7506 => x"55",
          7507 => x"55",
          7508 => x"81",
          7509 => x"74",
          7510 => x"56",
          7511 => x"12",
          7512 => x"70",
          7513 => x"38",
          7514 => x"81",
          7515 => x"51",
          7516 => x"51",
          7517 => x"89",
          7518 => x"70",
          7519 => x"53",
          7520 => x"70",
          7521 => x"51",
          7522 => x"09",
          7523 => x"38",
          7524 => x"38",
          7525 => x"77",
          7526 => x"70",
          7527 => x"2a",
          7528 => x"07",
          7529 => x"51",
          7530 => x"8f",
          7531 => x"84",
          7532 => x"83",
          7533 => x"94",
          7534 => x"74",
          7535 => x"38",
          7536 => x"0c",
          7537 => x"86",
          7538 => x"f4",
          7539 => x"82",
          7540 => x"8c",
          7541 => x"fa",
          7542 => x"56",
          7543 => x"17",
          7544 => x"b4",
          7545 => x"52",
          7546 => x"f4",
          7547 => x"82",
          7548 => x"81",
          7549 => x"b6",
          7550 => x"8a",
          7551 => x"98",
          7552 => x"ff",
          7553 => x"55",
          7554 => x"d5",
          7555 => x"06",
          7556 => x"80",
          7557 => x"33",
          7558 => x"81",
          7559 => x"81",
          7560 => x"81",
          7561 => x"eb",
          7562 => x"70",
          7563 => x"07",
          7564 => x"73",
          7565 => x"81",
          7566 => x"81",
          7567 => x"83",
          7568 => x"d8",
          7569 => x"16",
          7570 => x"3f",
          7571 => x"08",
          7572 => x"98",
          7573 => x"9d",
          7574 => x"82",
          7575 => x"81",
          7576 => x"ce",
          7577 => x"e0",
          7578 => x"82",
          7579 => x"80",
          7580 => x"82",
          7581 => x"e0",
          7582 => x"3d",
          7583 => x"3d",
          7584 => x"84",
          7585 => x"05",
          7586 => x"80",
          7587 => x"51",
          7588 => x"82",
          7589 => x"58",
          7590 => x"0b",
          7591 => x"08",
          7592 => x"38",
          7593 => x"08",
          7594 => x"f7",
          7595 => x"08",
          7596 => x"56",
          7597 => x"87",
          7598 => x"75",
          7599 => x"fe",
          7600 => x"54",
          7601 => x"2e",
          7602 => x"14",
          7603 => x"a0",
          7604 => x"98",
          7605 => x"06",
          7606 => x"54",
          7607 => x"38",
          7608 => x"87",
          7609 => x"82",
          7610 => x"06",
          7611 => x"56",
          7612 => x"38",
          7613 => x"80",
          7614 => x"18",
          7615 => x"8c",
          7616 => x"15",
          7617 => x"81",
          7618 => x"c6",
          7619 => x"e0",
          7620 => x"ff",
          7621 => x"06",
          7622 => x"56",
          7623 => x"38",
          7624 => x"8f",
          7625 => x"2a",
          7626 => x"51",
          7627 => x"72",
          7628 => x"80",
          7629 => x"52",
          7630 => x"3f",
          7631 => x"08",
          7632 => x"57",
          7633 => x"93",
          7634 => x"26",
          7635 => x"82",
          7636 => x"33",
          7637 => x"2e",
          7638 => x"8c",
          7639 => x"59",
          7640 => x"fa",
          7641 => x"58",
          7642 => x"2e",
          7643 => x"fe",
          7644 => x"a9",
          7645 => x"98",
          7646 => x"79",
          7647 => x"5b",
          7648 => x"90",
          7649 => x"75",
          7650 => x"38",
          7651 => x"e0",
          7652 => x"70",
          7653 => x"2a",
          7654 => x"95",
          7655 => x"29",
          7656 => x"5a",
          7657 => x"57",
          7658 => x"5b",
          7659 => x"80",
          7660 => x"7a",
          7661 => x"fc",
          7662 => x"e0",
          7663 => x"ff",
          7664 => x"0b",
          7665 => x"1a",
          7666 => x"72",
          7667 => x"81",
          7668 => x"81",
          7669 => x"27",
          7670 => x"80",
          7671 => x"81",
          7672 => x"56",
          7673 => x"27",
          7674 => x"56",
          7675 => x"84",
          7676 => x"56",
          7677 => x"84",
          7678 => x"c3",
          7679 => x"86",
          7680 => x"98",
          7681 => x"ff",
          7682 => x"84",
          7683 => x"81",
          7684 => x"38",
          7685 => x"51",
          7686 => x"82",
          7687 => x"83",
          7688 => x"58",
          7689 => x"80",
          7690 => x"c9",
          7691 => x"e0",
          7692 => x"77",
          7693 => x"80",
          7694 => x"82",
          7695 => x"c8",
          7696 => x"11",
          7697 => x"06",
          7698 => x"8d",
          7699 => x"26",
          7700 => x"74",
          7701 => x"78",
          7702 => x"c5",
          7703 => x"59",
          7704 => x"15",
          7705 => x"2e",
          7706 => x"13",
          7707 => x"72",
          7708 => x"38",
          7709 => x"f2",
          7710 => x"14",
          7711 => x"3f",
          7712 => x"08",
          7713 => x"98",
          7714 => x"23",
          7715 => x"57",
          7716 => x"83",
          7717 => x"cb",
          7718 => x"ea",
          7719 => x"98",
          7720 => x"ff",
          7721 => x"8d",
          7722 => x"14",
          7723 => x"3f",
          7724 => x"08",
          7725 => x"14",
          7726 => x"3f",
          7727 => x"08",
          7728 => x"06",
          7729 => x"72",
          7730 => x"9e",
          7731 => x"22",
          7732 => x"84",
          7733 => x"5a",
          7734 => x"83",
          7735 => x"14",
          7736 => x"79",
          7737 => x"d3",
          7738 => x"e0",
          7739 => x"82",
          7740 => x"80",
          7741 => x"38",
          7742 => x"08",
          7743 => x"ff",
          7744 => x"38",
          7745 => x"83",
          7746 => x"83",
          7747 => x"74",
          7748 => x"85",
          7749 => x"89",
          7750 => x"76",
          7751 => x"ca",
          7752 => x"70",
          7753 => x"7b",
          7754 => x"73",
          7755 => x"17",
          7756 => x"b0",
          7757 => x"55",
          7758 => x"09",
          7759 => x"38",
          7760 => x"51",
          7761 => x"82",
          7762 => x"83",
          7763 => x"53",
          7764 => x"82",
          7765 => x"82",
          7766 => x"e4",
          7767 => x"bd",
          7768 => x"98",
          7769 => x"0c",
          7770 => x"53",
          7771 => x"56",
          7772 => x"81",
          7773 => x"13",
          7774 => x"74",
          7775 => x"82",
          7776 => x"74",
          7777 => x"81",
          7778 => x"06",
          7779 => x"83",
          7780 => x"2a",
          7781 => x"72",
          7782 => x"26",
          7783 => x"ff",
          7784 => x"0c",
          7785 => x"15",
          7786 => x"0b",
          7787 => x"76",
          7788 => x"81",
          7789 => x"38",
          7790 => x"51",
          7791 => x"82",
          7792 => x"83",
          7793 => x"53",
          7794 => x"09",
          7795 => x"f9",
          7796 => x"52",
          7797 => x"88",
          7798 => x"98",
          7799 => x"38",
          7800 => x"08",
          7801 => x"84",
          7802 => x"c6",
          7803 => x"e0",
          7804 => x"ff",
          7805 => x"72",
          7806 => x"2e",
          7807 => x"80",
          7808 => x"14",
          7809 => x"3f",
          7810 => x"08",
          7811 => x"a4",
          7812 => x"81",
          7813 => x"84",
          7814 => x"c6",
          7815 => x"e0",
          7816 => x"8a",
          7817 => x"2e",
          7818 => x"9d",
          7819 => x"14",
          7820 => x"3f",
          7821 => x"08",
          7822 => x"84",
          7823 => x"c5",
          7824 => x"e0",
          7825 => x"15",
          7826 => x"34",
          7827 => x"22",
          7828 => x"72",
          7829 => x"23",
          7830 => x"23",
          7831 => x"0b",
          7832 => x"80",
          7833 => x"0c",
          7834 => x"82",
          7835 => x"90",
          7836 => x"fb",
          7837 => x"54",
          7838 => x"80",
          7839 => x"73",
          7840 => x"80",
          7841 => x"72",
          7842 => x"80",
          7843 => x"86",
          7844 => x"15",
          7845 => x"71",
          7846 => x"81",
          7847 => x"81",
          7848 => x"ff",
          7849 => x"82",
          7850 => x"81",
          7851 => x"88",
          7852 => x"08",
          7853 => x"39",
          7854 => x"73",
          7855 => x"74",
          7856 => x"0c",
          7857 => x"04",
          7858 => x"02",
          7859 => x"7a",
          7860 => x"fc",
          7861 => x"f4",
          7862 => x"54",
          7863 => x"e0",
          7864 => x"bc",
          7865 => x"98",
          7866 => x"82",
          7867 => x"70",
          7868 => x"73",
          7869 => x"38",
          7870 => x"78",
          7871 => x"2e",
          7872 => x"74",
          7873 => x"0c",
          7874 => x"80",
          7875 => x"80",
          7876 => x"70",
          7877 => x"51",
          7878 => x"82",
          7879 => x"54",
          7880 => x"98",
          7881 => x"0d",
          7882 => x"0d",
          7883 => x"05",
          7884 => x"33",
          7885 => x"54",
          7886 => x"84",
          7887 => x"bf",
          7888 => x"99",
          7889 => x"53",
          7890 => x"05",
          7891 => x"ae",
          7892 => x"98",
          7893 => x"e0",
          7894 => x"a4",
          7895 => x"69",
          7896 => x"70",
          7897 => x"b0",
          7898 => x"98",
          7899 => x"e0",
          7900 => x"38",
          7901 => x"05",
          7902 => x"2b",
          7903 => x"80",
          7904 => x"86",
          7905 => x"06",
          7906 => x"2e",
          7907 => x"74",
          7908 => x"38",
          7909 => x"09",
          7910 => x"38",
          7911 => x"b1",
          7912 => x"98",
          7913 => x"39",
          7914 => x"33",
          7915 => x"73",
          7916 => x"77",
          7917 => x"81",
          7918 => x"73",
          7919 => x"38",
          7920 => x"bc",
          7921 => x"07",
          7922 => x"b4",
          7923 => x"2a",
          7924 => x"51",
          7925 => x"2e",
          7926 => x"62",
          7927 => x"d6",
          7928 => x"e0",
          7929 => x"82",
          7930 => x"52",
          7931 => x"51",
          7932 => x"62",
          7933 => x"8b",
          7934 => x"53",
          7935 => x"51",
          7936 => x"80",
          7937 => x"05",
          7938 => x"3f",
          7939 => x"0b",
          7940 => x"75",
          7941 => x"f1",
          7942 => x"11",
          7943 => x"80",
          7944 => x"98",
          7945 => x"51",
          7946 => x"82",
          7947 => x"55",
          7948 => x"08",
          7949 => x"b7",
          7950 => x"c4",
          7951 => x"05",
          7952 => x"2a",
          7953 => x"51",
          7954 => x"80",
          7955 => x"84",
          7956 => x"39",
          7957 => x"70",
          7958 => x"54",
          7959 => x"a9",
          7960 => x"06",
          7961 => x"2e",
          7962 => x"55",
          7963 => x"73",
          7964 => x"c4",
          7965 => x"e0",
          7966 => x"ff",
          7967 => x"0c",
          7968 => x"e0",
          7969 => x"f8",
          7970 => x"2a",
          7971 => x"51",
          7972 => x"2e",
          7973 => x"80",
          7974 => x"7a",
          7975 => x"a0",
          7976 => x"a4",
          7977 => x"53",
          7978 => x"d5",
          7979 => x"e0",
          7980 => x"e0",
          7981 => x"1b",
          7982 => x"05",
          7983 => x"dd",
          7984 => x"98",
          7985 => x"98",
          7986 => x"0c",
          7987 => x"56",
          7988 => x"84",
          7989 => x"90",
          7990 => x"0b",
          7991 => x"80",
          7992 => x"0c",
          7993 => x"1a",
          7994 => x"2a",
          7995 => x"51",
          7996 => x"2e",
          7997 => x"82",
          7998 => x"80",
          7999 => x"38",
          8000 => x"08",
          8001 => x"8a",
          8002 => x"89",
          8003 => x"59",
          8004 => x"76",
          8005 => x"c5",
          8006 => x"e0",
          8007 => x"82",
          8008 => x"81",
          8009 => x"82",
          8010 => x"98",
          8011 => x"09",
          8012 => x"38",
          8013 => x"78",
          8014 => x"30",
          8015 => x"80",
          8016 => x"77",
          8017 => x"38",
          8018 => x"06",
          8019 => x"c3",
          8020 => x"1a",
          8021 => x"38",
          8022 => x"06",
          8023 => x"2e",
          8024 => x"52",
          8025 => x"ee",
          8026 => x"98",
          8027 => x"82",
          8028 => x"75",
          8029 => x"e0",
          8030 => x"9c",
          8031 => x"39",
          8032 => x"74",
          8033 => x"e0",
          8034 => x"3d",
          8035 => x"3d",
          8036 => x"65",
          8037 => x"5d",
          8038 => x"0c",
          8039 => x"05",
          8040 => x"f9",
          8041 => x"e0",
          8042 => x"82",
          8043 => x"8a",
          8044 => x"33",
          8045 => x"2e",
          8046 => x"56",
          8047 => x"90",
          8048 => x"06",
          8049 => x"74",
          8050 => x"b9",
          8051 => x"82",
          8052 => x"34",
          8053 => x"ad",
          8054 => x"91",
          8055 => x"56",
          8056 => x"8c",
          8057 => x"1a",
          8058 => x"74",
          8059 => x"38",
          8060 => x"80",
          8061 => x"38",
          8062 => x"70",
          8063 => x"56",
          8064 => x"b4",
          8065 => x"11",
          8066 => x"77",
          8067 => x"5b",
          8068 => x"38",
          8069 => x"88",
          8070 => x"8f",
          8071 => x"08",
          8072 => x"c3",
          8073 => x"e0",
          8074 => x"81",
          8075 => x"9f",
          8076 => x"2e",
          8077 => x"74",
          8078 => x"98",
          8079 => x"7e",
          8080 => x"3f",
          8081 => x"08",
          8082 => x"83",
          8083 => x"98",
          8084 => x"89",
          8085 => x"77",
          8086 => x"d8",
          8087 => x"7f",
          8088 => x"58",
          8089 => x"75",
          8090 => x"75",
          8091 => x"77",
          8092 => x"7c",
          8093 => x"33",
          8094 => x"91",
          8095 => x"98",
          8096 => x"38",
          8097 => x"33",
          8098 => x"80",
          8099 => x"b4",
          8100 => x"31",
          8101 => x"27",
          8102 => x"80",
          8103 => x"52",
          8104 => x"77",
          8105 => x"7d",
          8106 => x"bd",
          8107 => x"89",
          8108 => x"39",
          8109 => x"0c",
          8110 => x"83",
          8111 => x"80",
          8112 => x"55",
          8113 => x"83",
          8114 => x"9c",
          8115 => x"7e",
          8116 => x"3f",
          8117 => x"08",
          8118 => x"75",
          8119 => x"08",
          8120 => x"1f",
          8121 => x"7c",
          8122 => x"a9",
          8123 => x"31",
          8124 => x"7f",
          8125 => x"94",
          8126 => x"94",
          8127 => x"5c",
          8128 => x"80",
          8129 => x"e0",
          8130 => x"3d",
          8131 => x"3d",
          8132 => x"65",
          8133 => x"5d",
          8134 => x"0c",
          8135 => x"05",
          8136 => x"f6",
          8137 => x"e0",
          8138 => x"82",
          8139 => x"8a",
          8140 => x"33",
          8141 => x"2e",
          8142 => x"56",
          8143 => x"90",
          8144 => x"81",
          8145 => x"06",
          8146 => x"87",
          8147 => x"2e",
          8148 => x"95",
          8149 => x"91",
          8150 => x"56",
          8151 => x"81",
          8152 => x"34",
          8153 => x"95",
          8154 => x"08",
          8155 => x"56",
          8156 => x"84",
          8157 => x"5c",
          8158 => x"82",
          8159 => x"18",
          8160 => x"ff",
          8161 => x"74",
          8162 => x"7e",
          8163 => x"ff",
          8164 => x"2a",
          8165 => x"7a",
          8166 => x"8c",
          8167 => x"08",
          8168 => x"38",
          8169 => x"39",
          8170 => x"52",
          8171 => x"ac",
          8172 => x"98",
          8173 => x"e0",
          8174 => x"2e",
          8175 => x"74",
          8176 => x"91",
          8177 => x"2e",
          8178 => x"74",
          8179 => x"88",
          8180 => x"38",
          8181 => x"0c",
          8182 => x"15",
          8183 => x"08",
          8184 => x"06",
          8185 => x"51",
          8186 => x"3f",
          8187 => x"08",
          8188 => x"98",
          8189 => x"7e",
          8190 => x"da",
          8191 => x"98",
          8192 => x"fe",
          8193 => x"e0",
          8194 => x"7c",
          8195 => x"57",
          8196 => x"80",
          8197 => x"1b",
          8198 => x"22",
          8199 => x"75",
          8200 => x"38",
          8201 => x"59",
          8202 => x"53",
          8203 => x"1a",
          8204 => x"b6",
          8205 => x"e0",
          8206 => x"a3",
          8207 => x"11",
          8208 => x"56",
          8209 => x"27",
          8210 => x"80",
          8211 => x"08",
          8212 => x"2b",
          8213 => x"b8",
          8214 => x"ba",
          8215 => x"55",
          8216 => x"16",
          8217 => x"2b",
          8218 => x"39",
          8219 => x"94",
          8220 => x"94",
          8221 => x"ff",
          8222 => x"82",
          8223 => x"fd",
          8224 => x"77",
          8225 => x"55",
          8226 => x"0c",
          8227 => x"83",
          8228 => x"80",
          8229 => x"55",
          8230 => x"83",
          8231 => x"9c",
          8232 => x"7e",
          8233 => x"b8",
          8234 => x"98",
          8235 => x"38",
          8236 => x"52",
          8237 => x"83",
          8238 => x"b8",
          8239 => x"b9",
          8240 => x"55",
          8241 => x"16",
          8242 => x"31",
          8243 => x"7f",
          8244 => x"94",
          8245 => x"70",
          8246 => x"8c",
          8247 => x"58",
          8248 => x"76",
          8249 => x"75",
          8250 => x"19",
          8251 => x"39",
          8252 => x"80",
          8253 => x"74",
          8254 => x"80",
          8255 => x"e0",
          8256 => x"3d",
          8257 => x"3d",
          8258 => x"3d",
          8259 => x"70",
          8260 => x"df",
          8261 => x"98",
          8262 => x"e0",
          8263 => x"80",
          8264 => x"33",
          8265 => x"70",
          8266 => x"55",
          8267 => x"2e",
          8268 => x"a0",
          8269 => x"78",
          8270 => x"a4",
          8271 => x"98",
          8272 => x"e0",
          8273 => x"d8",
          8274 => x"08",
          8275 => x"a0",
          8276 => x"73",
          8277 => x"88",
          8278 => x"74",
          8279 => x"51",
          8280 => x"8c",
          8281 => x"9c",
          8282 => x"b7",
          8283 => x"88",
          8284 => x"96",
          8285 => x"b7",
          8286 => x"52",
          8287 => x"ff",
          8288 => x"78",
          8289 => x"83",
          8290 => x"51",
          8291 => x"3f",
          8292 => x"08",
          8293 => x"81",
          8294 => x"57",
          8295 => x"34",
          8296 => x"98",
          8297 => x"0d",
          8298 => x"0d",
          8299 => x"54",
          8300 => x"82",
          8301 => x"53",
          8302 => x"08",
          8303 => x"3d",
          8304 => x"73",
          8305 => x"3f",
          8306 => x"08",
          8307 => x"98",
          8308 => x"82",
          8309 => x"74",
          8310 => x"e0",
          8311 => x"3d",
          8312 => x"3d",
          8313 => x"51",
          8314 => x"8b",
          8315 => x"82",
          8316 => x"24",
          8317 => x"e0",
          8318 => x"f7",
          8319 => x"52",
          8320 => x"98",
          8321 => x"0d",
          8322 => x"0d",
          8323 => x"3d",
          8324 => x"95",
          8325 => x"e6",
          8326 => x"98",
          8327 => x"e0",
          8328 => x"e0",
          8329 => x"64",
          8330 => x"d0",
          8331 => x"e8",
          8332 => x"98",
          8333 => x"e0",
          8334 => x"38",
          8335 => x"05",
          8336 => x"2b",
          8337 => x"80",
          8338 => x"76",
          8339 => x"0c",
          8340 => x"02",
          8341 => x"70",
          8342 => x"81",
          8343 => x"56",
          8344 => x"9e",
          8345 => x"53",
          8346 => x"c9",
          8347 => x"e0",
          8348 => x"15",
          8349 => x"82",
          8350 => x"84",
          8351 => x"06",
          8352 => x"55",
          8353 => x"98",
          8354 => x"0d",
          8355 => x"3d",
          8356 => x"3d",
          8357 => x"3d",
          8358 => x"80",
          8359 => x"53",
          8360 => x"fd",
          8361 => x"80",
          8362 => x"e7",
          8363 => x"e0",
          8364 => x"82",
          8365 => x"83",
          8366 => x"80",
          8367 => x"7a",
          8368 => x"08",
          8369 => x"0c",
          8370 => x"d5",
          8371 => x"73",
          8372 => x"83",
          8373 => x"80",
          8374 => x"52",
          8375 => x"3f",
          8376 => x"08",
          8377 => x"98",
          8378 => x"38",
          8379 => x"08",
          8380 => x"ff",
          8381 => x"82",
          8382 => x"57",
          8383 => x"08",
          8384 => x"80",
          8385 => x"52",
          8386 => x"c2",
          8387 => x"98",
          8388 => x"3d",
          8389 => x"74",
          8390 => x"3f",
          8391 => x"08",
          8392 => x"98",
          8393 => x"38",
          8394 => x"51",
          8395 => x"82",
          8396 => x"57",
          8397 => x"08",
          8398 => x"da",
          8399 => x"7b",
          8400 => x"3f",
          8401 => x"98",
          8402 => x"38",
          8403 => x"51",
          8404 => x"82",
          8405 => x"57",
          8406 => x"08",
          8407 => x"38",
          8408 => x"09",
          8409 => x"38",
          8410 => x"ee",
          8411 => x"ea",
          8412 => x"3d",
          8413 => x"52",
          8414 => x"a0",
          8415 => x"3d",
          8416 => x"11",
          8417 => x"5a",
          8418 => x"2e",
          8419 => x"80",
          8420 => x"81",
          8421 => x"70",
          8422 => x"56",
          8423 => x"81",
          8424 => x"78",
          8425 => x"38",
          8426 => x"9c",
          8427 => x"82",
          8428 => x"18",
          8429 => x"08",
          8430 => x"ff",
          8431 => x"55",
          8432 => x"74",
          8433 => x"38",
          8434 => x"e1",
          8435 => x"55",
          8436 => x"34",
          8437 => x"77",
          8438 => x"81",
          8439 => x"ff",
          8440 => x"3d",
          8441 => x"58",
          8442 => x"80",
          8443 => x"f4",
          8444 => x"29",
          8445 => x"05",
          8446 => x"33",
          8447 => x"56",
          8448 => x"2e",
          8449 => x"16",
          8450 => x"33",
          8451 => x"73",
          8452 => x"16",
          8453 => x"26",
          8454 => x"55",
          8455 => x"91",
          8456 => x"54",
          8457 => x"70",
          8458 => x"34",
          8459 => x"ec",
          8460 => x"70",
          8461 => x"34",
          8462 => x"09",
          8463 => x"38",
          8464 => x"39",
          8465 => x"08",
          8466 => x"59",
          8467 => x"7a",
          8468 => x"5c",
          8469 => x"26",
          8470 => x"7a",
          8471 => x"e0",
          8472 => x"df",
          8473 => x"f7",
          8474 => x"7d",
          8475 => x"05",
          8476 => x"57",
          8477 => x"3f",
          8478 => x"08",
          8479 => x"98",
          8480 => x"38",
          8481 => x"53",
          8482 => x"38",
          8483 => x"54",
          8484 => x"92",
          8485 => x"33",
          8486 => x"70",
          8487 => x"54",
          8488 => x"38",
          8489 => x"15",
          8490 => x"70",
          8491 => x"58",
          8492 => x"82",
          8493 => x"8a",
          8494 => x"89",
          8495 => x"53",
          8496 => x"b7",
          8497 => x"ff",
          8498 => x"bc",
          8499 => x"e0",
          8500 => x"15",
          8501 => x"53",
          8502 => x"bb",
          8503 => x"e0",
          8504 => x"26",
          8505 => x"30",
          8506 => x"70",
          8507 => x"77",
          8508 => x"18",
          8509 => x"51",
          8510 => x"88",
          8511 => x"73",
          8512 => x"52",
          8513 => x"bb",
          8514 => x"e0",
          8515 => x"82",
          8516 => x"81",
          8517 => x"38",
          8518 => x"08",
          8519 => x"9e",
          8520 => x"98",
          8521 => x"0c",
          8522 => x"0c",
          8523 => x"81",
          8524 => x"76",
          8525 => x"38",
          8526 => x"94",
          8527 => x"94",
          8528 => x"16",
          8529 => x"2a",
          8530 => x"51",
          8531 => x"72",
          8532 => x"38",
          8533 => x"51",
          8534 => x"3f",
          8535 => x"08",
          8536 => x"98",
          8537 => x"82",
          8538 => x"56",
          8539 => x"52",
          8540 => x"b5",
          8541 => x"e0",
          8542 => x"73",
          8543 => x"38",
          8544 => x"b0",
          8545 => x"73",
          8546 => x"27",
          8547 => x"98",
          8548 => x"9e",
          8549 => x"08",
          8550 => x"0c",
          8551 => x"06",
          8552 => x"2e",
          8553 => x"52",
          8554 => x"b4",
          8555 => x"e0",
          8556 => x"38",
          8557 => x"16",
          8558 => x"80",
          8559 => x"0b",
          8560 => x"81",
          8561 => x"75",
          8562 => x"e0",
          8563 => x"58",
          8564 => x"54",
          8565 => x"74",
          8566 => x"73",
          8567 => x"90",
          8568 => x"c0",
          8569 => x"90",
          8570 => x"83",
          8571 => x"72",
          8572 => x"38",
          8573 => x"08",
          8574 => x"77",
          8575 => x"80",
          8576 => x"e0",
          8577 => x"3d",
          8578 => x"3d",
          8579 => x"89",
          8580 => x"2e",
          8581 => x"80",
          8582 => x"fc",
          8583 => x"3d",
          8584 => x"e0",
          8585 => x"e0",
          8586 => x"82",
          8587 => x"80",
          8588 => x"76",
          8589 => x"75",
          8590 => x"3f",
          8591 => x"08",
          8592 => x"98",
          8593 => x"38",
          8594 => x"70",
          8595 => x"57",
          8596 => x"a2",
          8597 => x"33",
          8598 => x"70",
          8599 => x"55",
          8600 => x"2e",
          8601 => x"16",
          8602 => x"51",
          8603 => x"82",
          8604 => x"88",
          8605 => x"54",
          8606 => x"84",
          8607 => x"52",
          8608 => x"bc",
          8609 => x"e0",
          8610 => x"74",
          8611 => x"81",
          8612 => x"85",
          8613 => x"74",
          8614 => x"38",
          8615 => x"74",
          8616 => x"e0",
          8617 => x"3d",
          8618 => x"3d",
          8619 => x"3d",
          8620 => x"70",
          8621 => x"bb",
          8622 => x"98",
          8623 => x"82",
          8624 => x"73",
          8625 => x"0d",
          8626 => x"0d",
          8627 => x"3d",
          8628 => x"71",
          8629 => x"e7",
          8630 => x"e0",
          8631 => x"82",
          8632 => x"80",
          8633 => x"94",
          8634 => x"98",
          8635 => x"51",
          8636 => x"3f",
          8637 => x"08",
          8638 => x"39",
          8639 => x"08",
          8640 => x"c1",
          8641 => x"e0",
          8642 => x"82",
          8643 => x"84",
          8644 => x"06",
          8645 => x"53",
          8646 => x"e0",
          8647 => x"38",
          8648 => x"51",
          8649 => x"72",
          8650 => x"ff",
          8651 => x"82",
          8652 => x"84",
          8653 => x"70",
          8654 => x"2c",
          8655 => x"98",
          8656 => x"51",
          8657 => x"82",
          8658 => x"87",
          8659 => x"ed",
          8660 => x"57",
          8661 => x"3d",
          8662 => x"3d",
          8663 => x"9e",
          8664 => x"98",
          8665 => x"e0",
          8666 => x"38",
          8667 => x"51",
          8668 => x"82",
          8669 => x"55",
          8670 => x"08",
          8671 => x"80",
          8672 => x"70",
          8673 => x"58",
          8674 => x"85",
          8675 => x"8d",
          8676 => x"2e",
          8677 => x"52",
          8678 => x"80",
          8679 => x"e0",
          8680 => x"3d",
          8681 => x"3d",
          8682 => x"55",
          8683 => x"92",
          8684 => x"52",
          8685 => x"dd",
          8686 => x"e0",
          8687 => x"82",
          8688 => x"82",
          8689 => x"74",
          8690 => x"9c",
          8691 => x"11",
          8692 => x"59",
          8693 => x"75",
          8694 => x"38",
          8695 => x"81",
          8696 => x"5b",
          8697 => x"82",
          8698 => x"39",
          8699 => x"08",
          8700 => x"59",
          8701 => x"09",
          8702 => x"c0",
          8703 => x"5f",
          8704 => x"92",
          8705 => x"51",
          8706 => x"3f",
          8707 => x"08",
          8708 => x"38",
          8709 => x"08",
          8710 => x"38",
          8711 => x"08",
          8712 => x"e0",
          8713 => x"80",
          8714 => x"81",
          8715 => x"59",
          8716 => x"14",
          8717 => x"c9",
          8718 => x"39",
          8719 => x"82",
          8720 => x"57",
          8721 => x"38",
          8722 => x"18",
          8723 => x"ff",
          8724 => x"82",
          8725 => x"5b",
          8726 => x"08",
          8727 => x"7c",
          8728 => x"12",
          8729 => x"52",
          8730 => x"82",
          8731 => x"06",
          8732 => x"14",
          8733 => x"8e",
          8734 => x"98",
          8735 => x"ff",
          8736 => x"70",
          8737 => x"82",
          8738 => x"51",
          8739 => x"b8",
          8740 => x"a9",
          8741 => x"e0",
          8742 => x"0a",
          8743 => x"70",
          8744 => x"84",
          8745 => x"51",
          8746 => x"ff",
          8747 => x"56",
          8748 => x"38",
          8749 => x"7c",
          8750 => x"0c",
          8751 => x"81",
          8752 => x"74",
          8753 => x"7a",
          8754 => x"0c",
          8755 => x"04",
          8756 => x"79",
          8757 => x"05",
          8758 => x"57",
          8759 => x"82",
          8760 => x"56",
          8761 => x"08",
          8762 => x"91",
          8763 => x"75",
          8764 => x"90",
          8765 => x"81",
          8766 => x"06",
          8767 => x"87",
          8768 => x"2e",
          8769 => x"94",
          8770 => x"73",
          8771 => x"27",
          8772 => x"73",
          8773 => x"e0",
          8774 => x"88",
          8775 => x"76",
          8776 => x"8c",
          8777 => x"98",
          8778 => x"19",
          8779 => x"ca",
          8780 => x"08",
          8781 => x"ff",
          8782 => x"82",
          8783 => x"ff",
          8784 => x"06",
          8785 => x"56",
          8786 => x"08",
          8787 => x"81",
          8788 => x"82",
          8789 => x"75",
          8790 => x"54",
          8791 => x"08",
          8792 => x"27",
          8793 => x"17",
          8794 => x"e0",
          8795 => x"76",
          8796 => x"bc",
          8797 => x"98",
          8798 => x"17",
          8799 => x"0c",
          8800 => x"80",
          8801 => x"73",
          8802 => x"75",
          8803 => x"38",
          8804 => x"34",
          8805 => x"82",
          8806 => x"89",
          8807 => x"e0",
          8808 => x"53",
          8809 => x"9c",
          8810 => x"3d",
          8811 => x"3f",
          8812 => x"08",
          8813 => x"98",
          8814 => x"38",
          8815 => x"3d",
          8816 => x"3d",
          8817 => x"cd",
          8818 => x"e0",
          8819 => x"82",
          8820 => x"81",
          8821 => x"80",
          8822 => x"70",
          8823 => x"81",
          8824 => x"56",
          8825 => x"81",
          8826 => x"98",
          8827 => x"74",
          8828 => x"38",
          8829 => x"05",
          8830 => x"06",
          8831 => x"55",
          8832 => x"38",
          8833 => x"51",
          8834 => x"3f",
          8835 => x"08",
          8836 => x"70",
          8837 => x"55",
          8838 => x"2e",
          8839 => x"78",
          8840 => x"98",
          8841 => x"08",
          8842 => x"38",
          8843 => x"e0",
          8844 => x"76",
          8845 => x"70",
          8846 => x"b5",
          8847 => x"e0",
          8848 => x"82",
          8849 => x"80",
          8850 => x"e0",
          8851 => x"73",
          8852 => x"90",
          8853 => x"98",
          8854 => x"e0",
          8855 => x"38",
          8856 => x"d0",
          8857 => x"98",
          8858 => x"88",
          8859 => x"98",
          8860 => x"38",
          8861 => x"ab",
          8862 => x"98",
          8863 => x"98",
          8864 => x"82",
          8865 => x"07",
          8866 => x"55",
          8867 => x"2e",
          8868 => x"80",
          8869 => x"80",
          8870 => x"77",
          8871 => x"90",
          8872 => x"98",
          8873 => x"8c",
          8874 => x"ff",
          8875 => x"82",
          8876 => x"55",
          8877 => x"98",
          8878 => x"0d",
          8879 => x"0d",
          8880 => x"3d",
          8881 => x"52",
          8882 => x"d7",
          8883 => x"e0",
          8884 => x"82",
          8885 => x"82",
          8886 => x"5e",
          8887 => x"3d",
          8888 => x"cb",
          8889 => x"e0",
          8890 => x"82",
          8891 => x"86",
          8892 => x"82",
          8893 => x"e0",
          8894 => x"2e",
          8895 => x"82",
          8896 => x"80",
          8897 => x"70",
          8898 => x"06",
          8899 => x"54",
          8900 => x"38",
          8901 => x"52",
          8902 => x"52",
          8903 => x"bc",
          8904 => x"98",
          8905 => x"56",
          8906 => x"08",
          8907 => x"54",
          8908 => x"08",
          8909 => x"81",
          8910 => x"82",
          8911 => x"98",
          8912 => x"09",
          8913 => x"38",
          8914 => x"ba",
          8915 => x"b6",
          8916 => x"98",
          8917 => x"51",
          8918 => x"3f",
          8919 => x"08",
          8920 => x"98",
          8921 => x"38",
          8922 => x"52",
          8923 => x"ff",
          8924 => x"78",
          8925 => x"b8",
          8926 => x"54",
          8927 => x"c3",
          8928 => x"88",
          8929 => x"80",
          8930 => x"ff",
          8931 => x"75",
          8932 => x"11",
          8933 => x"b7",
          8934 => x"53",
          8935 => x"53",
          8936 => x"51",
          8937 => x"3f",
          8938 => x"0b",
          8939 => x"34",
          8940 => x"80",
          8941 => x"51",
          8942 => x"3f",
          8943 => x"0b",
          8944 => x"77",
          8945 => x"89",
          8946 => x"98",
          8947 => x"e0",
          8948 => x"38",
          8949 => x"0a",
          8950 => x"05",
          8951 => x"86",
          8952 => x"64",
          8953 => x"ff",
          8954 => x"64",
          8955 => x"8b",
          8956 => x"54",
          8957 => x"15",
          8958 => x"ff",
          8959 => x"82",
          8960 => x"54",
          8961 => x"53",
          8962 => x"51",
          8963 => x"3f",
          8964 => x"98",
          8965 => x"0d",
          8966 => x"0d",
          8967 => x"05",
          8968 => x"3f",
          8969 => x"3d",
          8970 => x"52",
          8971 => x"d4",
          8972 => x"e0",
          8973 => x"82",
          8974 => x"82",
          8975 => x"4e",
          8976 => x"52",
          8977 => x"52",
          8978 => x"3f",
          8979 => x"08",
          8980 => x"98",
          8981 => x"38",
          8982 => x"05",
          8983 => x"06",
          8984 => x"73",
          8985 => x"a0",
          8986 => x"08",
          8987 => x"ff",
          8988 => x"ff",
          8989 => x"b0",
          8990 => x"92",
          8991 => x"54",
          8992 => x"3f",
          8993 => x"52",
          8994 => x"8c",
          8995 => x"98",
          8996 => x"e0",
          8997 => x"38",
          8998 => x"08",
          8999 => x"06",
          9000 => x"a3",
          9001 => x"92",
          9002 => x"81",
          9003 => x"e0",
          9004 => x"2e",
          9005 => x"81",
          9006 => x"51",
          9007 => x"3f",
          9008 => x"08",
          9009 => x"98",
          9010 => x"38",
          9011 => x"53",
          9012 => x"8d",
          9013 => x"16",
          9014 => x"b9",
          9015 => x"05",
          9016 => x"34",
          9017 => x"70",
          9018 => x"81",
          9019 => x"55",
          9020 => x"74",
          9021 => x"73",
          9022 => x"78",
          9023 => x"83",
          9024 => x"16",
          9025 => x"2a",
          9026 => x"51",
          9027 => x"80",
          9028 => x"38",
          9029 => x"80",
          9030 => x"52",
          9031 => x"b4",
          9032 => x"e0",
          9033 => x"78",
          9034 => x"aa",
          9035 => x"82",
          9036 => x"80",
          9037 => x"38",
          9038 => x"08",
          9039 => x"ff",
          9040 => x"82",
          9041 => x"79",
          9042 => x"58",
          9043 => x"e0",
          9044 => x"c1",
          9045 => x"33",
          9046 => x"2e",
          9047 => x"9a",
          9048 => x"75",
          9049 => x"ff",
          9050 => x"78",
          9051 => x"83",
          9052 => x"39",
          9053 => x"08",
          9054 => x"51",
          9055 => x"82",
          9056 => x"55",
          9057 => x"08",
          9058 => x"51",
          9059 => x"3f",
          9060 => x"08",
          9061 => x"e0",
          9062 => x"3d",
          9063 => x"3d",
          9064 => x"df",
          9065 => x"84",
          9066 => x"05",
          9067 => x"82",
          9068 => x"cc",
          9069 => x"3d",
          9070 => x"3f",
          9071 => x"08",
          9072 => x"98",
          9073 => x"38",
          9074 => x"52",
          9075 => x"05",
          9076 => x"3f",
          9077 => x"08",
          9078 => x"98",
          9079 => x"02",
          9080 => x"33",
          9081 => x"54",
          9082 => x"aa",
          9083 => x"06",
          9084 => x"8b",
          9085 => x"06",
          9086 => x"07",
          9087 => x"56",
          9088 => x"34",
          9089 => x"0b",
          9090 => x"78",
          9091 => x"97",
          9092 => x"98",
          9093 => x"82",
          9094 => x"96",
          9095 => x"ee",
          9096 => x"56",
          9097 => x"3d",
          9098 => x"95",
          9099 => x"ce",
          9100 => x"98",
          9101 => x"e0",
          9102 => x"cb",
          9103 => x"64",
          9104 => x"d0",
          9105 => x"d0",
          9106 => x"98",
          9107 => x"e0",
          9108 => x"38",
          9109 => x"05",
          9110 => x"06",
          9111 => x"73",
          9112 => x"16",
          9113 => x"22",
          9114 => x"07",
          9115 => x"1f",
          9116 => x"f2",
          9117 => x"81",
          9118 => x"34",
          9119 => x"a1",
          9120 => x"e0",
          9121 => x"74",
          9122 => x"0c",
          9123 => x"04",
          9124 => x"6a",
          9125 => x"80",
          9126 => x"cc",
          9127 => x"3d",
          9128 => x"3f",
          9129 => x"08",
          9130 => x"08",
          9131 => x"e0",
          9132 => x"80",
          9133 => x"57",
          9134 => x"81",
          9135 => x"70",
          9136 => x"55",
          9137 => x"80",
          9138 => x"5d",
          9139 => x"52",
          9140 => x"52",
          9141 => x"97",
          9142 => x"98",
          9143 => x"e0",
          9144 => x"d2",
          9145 => x"73",
          9146 => x"f8",
          9147 => x"98",
          9148 => x"e0",
          9149 => x"38",
          9150 => x"08",
          9151 => x"08",
          9152 => x"56",
          9153 => x"19",
          9154 => x"59",
          9155 => x"74",
          9156 => x"56",
          9157 => x"ec",
          9158 => x"75",
          9159 => x"74",
          9160 => x"2e",
          9161 => x"16",
          9162 => x"33",
          9163 => x"73",
          9164 => x"38",
          9165 => x"84",
          9166 => x"06",
          9167 => x"7a",
          9168 => x"76",
          9169 => x"07",
          9170 => x"54",
          9171 => x"80",
          9172 => x"80",
          9173 => x"7b",
          9174 => x"53",
          9175 => x"80",
          9176 => x"98",
          9177 => x"e0",
          9178 => x"38",
          9179 => x"55",
          9180 => x"56",
          9181 => x"8b",
          9182 => x"56",
          9183 => x"83",
          9184 => x"75",
          9185 => x"51",
          9186 => x"3f",
          9187 => x"08",
          9188 => x"82",
          9189 => x"99",
          9190 => x"e6",
          9191 => x"53",
          9192 => x"b4",
          9193 => x"3d",
          9194 => x"3f",
          9195 => x"08",
          9196 => x"08",
          9197 => x"e0",
          9198 => x"dd",
          9199 => x"a0",
          9200 => x"70",
          9201 => x"9b",
          9202 => x"6d",
          9203 => x"55",
          9204 => x"27",
          9205 => x"77",
          9206 => x"51",
          9207 => x"3f",
          9208 => x"08",
          9209 => x"26",
          9210 => x"82",
          9211 => x"51",
          9212 => x"83",
          9213 => x"e0",
          9214 => x"95",
          9215 => x"e0",
          9216 => x"ff",
          9217 => x"74",
          9218 => x"38",
          9219 => x"d3",
          9220 => x"9b",
          9221 => x"e0",
          9222 => x"38",
          9223 => x"27",
          9224 => x"89",
          9225 => x"8b",
          9226 => x"27",
          9227 => x"55",
          9228 => x"81",
          9229 => x"8f",
          9230 => x"2a",
          9231 => x"70",
          9232 => x"34",
          9233 => x"74",
          9234 => x"05",
          9235 => x"16",
          9236 => x"51",
          9237 => x"9f",
          9238 => x"38",
          9239 => x"54",
          9240 => x"81",
          9241 => x"b1",
          9242 => x"2e",
          9243 => x"a3",
          9244 => x"15",
          9245 => x"54",
          9246 => x"09",
          9247 => x"38",
          9248 => x"75",
          9249 => x"40",
          9250 => x"52",
          9251 => x"52",
          9252 => x"db",
          9253 => x"98",
          9254 => x"e0",
          9255 => x"f7",
          9256 => x"74",
          9257 => x"bc",
          9258 => x"98",
          9259 => x"e0",
          9260 => x"38",
          9261 => x"38",
          9262 => x"74",
          9263 => x"39",
          9264 => x"08",
          9265 => x"81",
          9266 => x"38",
          9267 => x"74",
          9268 => x"38",
          9269 => x"51",
          9270 => x"3f",
          9271 => x"08",
          9272 => x"98",
          9273 => x"a0",
          9274 => x"98",
          9275 => x"51",
          9276 => x"3f",
          9277 => x"0b",
          9278 => x"8b",
          9279 => x"66",
          9280 => x"91",
          9281 => x"81",
          9282 => x"34",
          9283 => x"9c",
          9284 => x"e0",
          9285 => x"73",
          9286 => x"e0",
          9287 => x"3d",
          9288 => x"3d",
          9289 => x"02",
          9290 => x"cb",
          9291 => x"3d",
          9292 => x"72",
          9293 => x"5a",
          9294 => x"82",
          9295 => x"58",
          9296 => x"08",
          9297 => x"91",
          9298 => x"77",
          9299 => x"7c",
          9300 => x"38",
          9301 => x"59",
          9302 => x"90",
          9303 => x"81",
          9304 => x"06",
          9305 => x"73",
          9306 => x"54",
          9307 => x"82",
          9308 => x"39",
          9309 => x"8b",
          9310 => x"11",
          9311 => x"2b",
          9312 => x"54",
          9313 => x"fe",
          9314 => x"ff",
          9315 => x"70",
          9316 => x"07",
          9317 => x"e0",
          9318 => x"90",
          9319 => x"40",
          9320 => x"55",
          9321 => x"88",
          9322 => x"08",
          9323 => x"38",
          9324 => x"77",
          9325 => x"56",
          9326 => x"51",
          9327 => x"3f",
          9328 => x"55",
          9329 => x"08",
          9330 => x"38",
          9331 => x"e0",
          9332 => x"2e",
          9333 => x"82",
          9334 => x"ff",
          9335 => x"38",
          9336 => x"08",
          9337 => x"16",
          9338 => x"2e",
          9339 => x"87",
          9340 => x"74",
          9341 => x"74",
          9342 => x"81",
          9343 => x"38",
          9344 => x"ff",
          9345 => x"2e",
          9346 => x"7b",
          9347 => x"80",
          9348 => x"81",
          9349 => x"81",
          9350 => x"06",
          9351 => x"56",
          9352 => x"52",
          9353 => x"9d",
          9354 => x"e0",
          9355 => x"82",
          9356 => x"80",
          9357 => x"81",
          9358 => x"56",
          9359 => x"d3",
          9360 => x"ff",
          9361 => x"7c",
          9362 => x"55",
          9363 => x"b3",
          9364 => x"1b",
          9365 => x"1b",
          9366 => x"33",
          9367 => x"54",
          9368 => x"34",
          9369 => x"fe",
          9370 => x"08",
          9371 => x"74",
          9372 => x"75",
          9373 => x"16",
          9374 => x"33",
          9375 => x"73",
          9376 => x"77",
          9377 => x"e0",
          9378 => x"3d",
          9379 => x"3d",
          9380 => x"02",
          9381 => x"ef",
          9382 => x"3d",
          9383 => x"59",
          9384 => x"8b",
          9385 => x"82",
          9386 => x"24",
          9387 => x"82",
          9388 => x"84",
          9389 => x"e0",
          9390 => x"51",
          9391 => x"2e",
          9392 => x"75",
          9393 => x"98",
          9394 => x"98",
          9395 => x"e0",
          9396 => x"82",
          9397 => x"33",
          9398 => x"81",
          9399 => x"ff",
          9400 => x"82",
          9401 => x"81",
          9402 => x"81",
          9403 => x"83",
          9404 => x"da",
          9405 => x"2a",
          9406 => x"51",
          9407 => x"74",
          9408 => x"9a",
          9409 => x"53",
          9410 => x"51",
          9411 => x"3f",
          9412 => x"08",
          9413 => x"55",
          9414 => x"92",
          9415 => x"80",
          9416 => x"38",
          9417 => x"06",
          9418 => x"2e",
          9419 => x"49",
          9420 => x"87",
          9421 => x"79",
          9422 => x"78",
          9423 => x"26",
          9424 => x"19",
          9425 => x"74",
          9426 => x"38",
          9427 => x"fe",
          9428 => x"2a",
          9429 => x"70",
          9430 => x"59",
          9431 => x"7a",
          9432 => x"56",
          9433 => x"80",
          9434 => x"51",
          9435 => x"74",
          9436 => x"64",
          9437 => x"e0",
          9438 => x"74",
          9439 => x"7f",
          9440 => x"89",
          9441 => x"82",
          9442 => x"8b",
          9443 => x"fe",
          9444 => x"92",
          9445 => x"e0",
          9446 => x"ff",
          9447 => x"8e",
          9448 => x"d4",
          9449 => x"81",
          9450 => x"38",
          9451 => x"1b",
          9452 => x"33",
          9453 => x"80",
          9454 => x"38",
          9455 => x"51",
          9456 => x"3f",
          9457 => x"08",
          9458 => x"52",
          9459 => x"cd",
          9460 => x"98",
          9461 => x"39",
          9462 => x"05",
          9463 => x"7f",
          9464 => x"f7",
          9465 => x"82",
          9466 => x"8a",
          9467 => x"83",
          9468 => x"06",
          9469 => x"08",
          9470 => x"74",
          9471 => x"5f",
          9472 => x"56",
          9473 => x"8a",
          9474 => x"7f",
          9475 => x"56",
          9476 => x"27",
          9477 => x"93",
          9478 => x"80",
          9479 => x"38",
          9480 => x"70",
          9481 => x"44",
          9482 => x"95",
          9483 => x"06",
          9484 => x"2e",
          9485 => x"62",
          9486 => x"74",
          9487 => x"83",
          9488 => x"06",
          9489 => x"82",
          9490 => x"2e",
          9491 => x"78",
          9492 => x"2e",
          9493 => x"80",
          9494 => x"ae",
          9495 => x"2a",
          9496 => x"82",
          9497 => x"56",
          9498 => x"2e",
          9499 => x"77",
          9500 => x"82",
          9501 => x"79",
          9502 => x"70",
          9503 => x"5a",
          9504 => x"86",
          9505 => x"27",
          9506 => x"52",
          9507 => x"9c",
          9508 => x"e0",
          9509 => x"29",
          9510 => x"70",
          9511 => x"55",
          9512 => x"0b",
          9513 => x"08",
          9514 => x"05",
          9515 => x"ff",
          9516 => x"27",
          9517 => x"89",
          9518 => x"ae",
          9519 => x"2a",
          9520 => x"82",
          9521 => x"56",
          9522 => x"2e",
          9523 => x"77",
          9524 => x"82",
          9525 => x"79",
          9526 => x"70",
          9527 => x"5a",
          9528 => x"86",
          9529 => x"27",
          9530 => x"52",
          9531 => x"9b",
          9532 => x"e0",
          9533 => x"84",
          9534 => x"e0",
          9535 => x"f5",
          9536 => x"81",
          9537 => x"98",
          9538 => x"e0",
          9539 => x"71",
          9540 => x"83",
          9541 => x"5e",
          9542 => x"89",
          9543 => x"5c",
          9544 => x"1f",
          9545 => x"05",
          9546 => x"ff",
          9547 => x"70",
          9548 => x"31",
          9549 => x"57",
          9550 => x"83",
          9551 => x"06",
          9552 => x"1c",
          9553 => x"5c",
          9554 => x"1d",
          9555 => x"29",
          9556 => x"31",
          9557 => x"55",
          9558 => x"87",
          9559 => x"7c",
          9560 => x"7a",
          9561 => x"31",
          9562 => x"9a",
          9563 => x"e0",
          9564 => x"7d",
          9565 => x"81",
          9566 => x"82",
          9567 => x"83",
          9568 => x"80",
          9569 => x"87",
          9570 => x"81",
          9571 => x"fd",
          9572 => x"ad",
          9573 => x"2e",
          9574 => x"80",
          9575 => x"ff",
          9576 => x"e0",
          9577 => x"a0",
          9578 => x"38",
          9579 => x"74",
          9580 => x"86",
          9581 => x"fd",
          9582 => x"81",
          9583 => x"80",
          9584 => x"83",
          9585 => x"39",
          9586 => x"08",
          9587 => x"92",
          9588 => x"ed",
          9589 => x"59",
          9590 => x"27",
          9591 => x"86",
          9592 => x"55",
          9593 => x"09",
          9594 => x"38",
          9595 => x"f5",
          9596 => x"38",
          9597 => x"55",
          9598 => x"86",
          9599 => x"80",
          9600 => x"7a",
          9601 => x"b0",
          9602 => x"82",
          9603 => x"7a",
          9604 => x"81",
          9605 => x"52",
          9606 => x"ff",
          9607 => x"79",
          9608 => x"7b",
          9609 => x"06",
          9610 => x"51",
          9611 => x"3f",
          9612 => x"1c",
          9613 => x"32",
          9614 => x"96",
          9615 => x"06",
          9616 => x"91",
          9617 => x"8d",
          9618 => x"55",
          9619 => x"ff",
          9620 => x"74",
          9621 => x"06",
          9622 => x"51",
          9623 => x"3f",
          9624 => x"52",
          9625 => x"ff",
          9626 => x"f8",
          9627 => x"34",
          9628 => x"1b",
          9629 => x"d0",
          9630 => x"52",
          9631 => x"ff",
          9632 => x"7e",
          9633 => x"51",
          9634 => x"3f",
          9635 => x"09",
          9636 => x"cb",
          9637 => x"b2",
          9638 => x"c3",
          9639 => x"8d",
          9640 => x"52",
          9641 => x"ff",
          9642 => x"82",
          9643 => x"51",
          9644 => x"3f",
          9645 => x"1b",
          9646 => x"8c",
          9647 => x"b2",
          9648 => x"8d",
          9649 => x"80",
          9650 => x"1c",
          9651 => x"80",
          9652 => x"93",
          9653 => x"f0",
          9654 => x"1b",
          9655 => x"82",
          9656 => x"52",
          9657 => x"ff",
          9658 => x"7c",
          9659 => x"06",
          9660 => x"51",
          9661 => x"3f",
          9662 => x"a4",
          9663 => x"0b",
          9664 => x"93",
          9665 => x"84",
          9666 => x"51",
          9667 => x"3f",
          9668 => x"52",
          9669 => x"70",
          9670 => x"8c",
          9671 => x"54",
          9672 => x"52",
          9673 => x"88",
          9674 => x"56",
          9675 => x"08",
          9676 => x"7d",
          9677 => x"81",
          9678 => x"38",
          9679 => x"1f",
          9680 => x"7f",
          9681 => x"af",
          9682 => x"53",
          9683 => x"51",
          9684 => x"3f",
          9685 => x"a4",
          9686 => x"51",
          9687 => x"3f",
          9688 => x"e4",
          9689 => x"e4",
          9690 => x"8b",
          9691 => x"18",
          9692 => x"1b",
          9693 => x"ee",
          9694 => x"83",
          9695 => x"ff",
          9696 => x"82",
          9697 => x"78",
          9698 => x"bc",
          9699 => x"87",
          9700 => x"52",
          9701 => x"87",
          9702 => x"54",
          9703 => x"7a",
          9704 => x"ff",
          9705 => x"66",
          9706 => x"7a",
          9707 => x"88",
          9708 => x"80",
          9709 => x"2e",
          9710 => x"9a",
          9711 => x"7a",
          9712 => x"a2",
          9713 => x"84",
          9714 => x"8b",
          9715 => x"0a",
          9716 => x"51",
          9717 => x"ff",
          9718 => x"7d",
          9719 => x"38",
          9720 => x"52",
          9721 => x"8a",
          9722 => x"55",
          9723 => x"62",
          9724 => x"74",
          9725 => x"75",
          9726 => x"7f",
          9727 => x"f7",
          9728 => x"98",
          9729 => x"38",
          9730 => x"82",
          9731 => x"52",
          9732 => x"8b",
          9733 => x"16",
          9734 => x"56",
          9735 => x"38",
          9736 => x"77",
          9737 => x"8d",
          9738 => x"7d",
          9739 => x"38",
          9740 => x"57",
          9741 => x"83",
          9742 => x"76",
          9743 => x"7a",
          9744 => x"ff",
          9745 => x"82",
          9746 => x"81",
          9747 => x"16",
          9748 => x"56",
          9749 => x"38",
          9750 => x"83",
          9751 => x"86",
          9752 => x"ff",
          9753 => x"38",
          9754 => x"82",
          9755 => x"81",
          9756 => x"2e",
          9757 => x"54",
          9758 => x"52",
          9759 => x"84",
          9760 => x"56",
          9761 => x"08",
          9762 => x"64",
          9763 => x"55",
          9764 => x"16",
          9765 => x"82",
          9766 => x"53",
          9767 => x"51",
          9768 => x"3f",
          9769 => x"62",
          9770 => x"06",
          9771 => x"fd",
          9772 => x"53",
          9773 => x"51",
          9774 => x"3f",
          9775 => x"52",
          9776 => x"89",
          9777 => x"be",
          9778 => x"75",
          9779 => x"81",
          9780 => x"0b",
          9781 => x"77",
          9782 => x"76",
          9783 => x"67",
          9784 => x"fd",
          9785 => x"51",
          9786 => x"3f",
          9787 => x"16",
          9788 => x"98",
          9789 => x"bf",
          9790 => x"86",
          9791 => x"e0",
          9792 => x"16",
          9793 => x"83",
          9794 => x"ff",
          9795 => x"67",
          9796 => x"1b",
          9797 => x"ce",
          9798 => x"77",
          9799 => x"7f",
          9800 => x"d3",
          9801 => x"82",
          9802 => x"a2",
          9803 => x"80",
          9804 => x"ff",
          9805 => x"81",
          9806 => x"98",
          9807 => x"89",
          9808 => x"8a",
          9809 => x"86",
          9810 => x"98",
          9811 => x"82",
          9812 => x"9a",
          9813 => x"f5",
          9814 => x"60",
          9815 => x"79",
          9816 => x"5a",
          9817 => x"78",
          9818 => x"8d",
          9819 => x"55",
          9820 => x"fc",
          9821 => x"51",
          9822 => x"7a",
          9823 => x"81",
          9824 => x"8c",
          9825 => x"74",
          9826 => x"38",
          9827 => x"81",
          9828 => x"81",
          9829 => x"8a",
          9830 => x"06",
          9831 => x"76",
          9832 => x"76",
          9833 => x"55",
          9834 => x"98",
          9835 => x"0d",
          9836 => x"0d",
          9837 => x"05",
          9838 => x"59",
          9839 => x"2e",
          9840 => x"87",
          9841 => x"76",
          9842 => x"84",
          9843 => x"80",
          9844 => x"38",
          9845 => x"77",
          9846 => x"56",
          9847 => x"34",
          9848 => x"bb",
          9849 => x"38",
          9850 => x"05",
          9851 => x"8c",
          9852 => x"08",
          9853 => x"3f",
          9854 => x"70",
          9855 => x"07",
          9856 => x"30",
          9857 => x"56",
          9858 => x"0c",
          9859 => x"18",
          9860 => x"0d",
          9861 => x"0d",
          9862 => x"08",
          9863 => x"75",
          9864 => x"89",
          9865 => x"54",
          9866 => x"16",
          9867 => x"51",
          9868 => x"82",
          9869 => x"91",
          9870 => x"08",
          9871 => x"81",
          9872 => x"88",
          9873 => x"83",
          9874 => x"74",
          9875 => x"0c",
          9876 => x"04",
          9877 => x"75",
          9878 => x"53",
          9879 => x"51",
          9880 => x"3f",
          9881 => x"85",
          9882 => x"ea",
          9883 => x"80",
          9884 => x"6a",
          9885 => x"70",
          9886 => x"d8",
          9887 => x"72",
          9888 => x"3f",
          9889 => x"8d",
          9890 => x"0d",
          9891 => x"0d",
          9892 => x"05",
          9893 => x"55",
          9894 => x"72",
          9895 => x"8a",
          9896 => x"ff",
          9897 => x"80",
          9898 => x"ff",
          9899 => x"51",
          9900 => x"2e",
          9901 => x"b4",
          9902 => x"2e",
          9903 => x"d3",
          9904 => x"72",
          9905 => x"38",
          9906 => x"83",
          9907 => x"53",
          9908 => x"ff",
          9909 => x"71",
          9910 => x"ec",
          9911 => x"51",
          9912 => x"81",
          9913 => x"81",
          9914 => x"51",
          9915 => x"98",
          9916 => x"0d",
          9917 => x"0d",
          9918 => x"22",
          9919 => x"96",
          9920 => x"51",
          9921 => x"80",
          9922 => x"38",
          9923 => x"39",
          9924 => x"2e",
          9925 => x"91",
          9926 => x"ff",
          9927 => x"70",
          9928 => x"ec",
          9929 => x"54",
          9930 => x"e0",
          9931 => x"3d",
          9932 => x"3d",
          9933 => x"70",
          9934 => x"26",
          9935 => x"70",
          9936 => x"06",
          9937 => x"57",
          9938 => x"72",
          9939 => x"82",
          9940 => x"75",
          9941 => x"57",
          9942 => x"70",
          9943 => x"75",
          9944 => x"52",
          9945 => x"fb",
          9946 => x"82",
          9947 => x"70",
          9948 => x"81",
          9949 => x"18",
          9950 => x"53",
          9951 => x"80",
          9952 => x"88",
          9953 => x"38",
          9954 => x"82",
          9955 => x"51",
          9956 => x"71",
          9957 => x"76",
          9958 => x"54",
          9959 => x"c3",
          9960 => x"31",
          9961 => x"71",
          9962 => x"a4",
          9963 => x"51",
          9964 => x"12",
          9965 => x"d0",
          9966 => x"39",
          9967 => x"90",
          9968 => x"51",
          9969 => x"b0",
          9970 => x"39",
          9971 => x"51",
          9972 => x"ff",
          9973 => x"39",
          9974 => x"38",
          9975 => x"56",
          9976 => x"71",
          9977 => x"e0",
          9978 => x"3d",
          9979 => x"ff",
          9980 => x"00",
          9981 => x"ff",
          9982 => x"ff",
          9983 => x"00",
          9984 => x"00",
          9985 => x"00",
          9986 => x"00",
          9987 => x"00",
          9988 => x"00",
          9989 => x"00",
          9990 => x"00",
          9991 => x"00",
          9992 => x"00",
          9993 => x"00",
          9994 => x"00",
          9995 => x"00",
          9996 => x"00",
          9997 => x"00",
          9998 => x"00",
          9999 => x"00",
         10000 => x"00",
         10001 => x"00",
         10002 => x"00",
         10003 => x"00",
         10004 => x"00",
         10005 => x"00",
         10006 => x"00",
         10007 => x"00",
         10008 => x"00",
         10009 => x"00",
         10010 => x"00",
         10011 => x"00",
         10012 => x"00",
         10013 => x"00",
         10014 => x"00",
         10015 => x"00",
         10016 => x"00",
         10017 => x"00",
         10018 => x"00",
         10019 => x"00",
         10020 => x"00",
         10021 => x"00",
         10022 => x"00",
         10023 => x"00",
         10024 => x"00",
         10025 => x"00",
         10026 => x"00",
         10027 => x"00",
         10028 => x"00",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"00",
         10033 => x"00",
         10034 => x"00",
         10035 => x"00",
         10036 => x"00",
         10037 => x"00",
         10038 => x"00",
         10039 => x"00",
         10040 => x"00",
         10041 => x"00",
         10042 => x"00",
         10043 => x"00",
         10044 => x"00",
         10045 => x"00",
         10046 => x"00",
         10047 => x"00",
         10048 => x"00",
         10049 => x"00",
         10050 => x"00",
         10051 => x"00",
         10052 => x"00",
         10053 => x"00",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"00",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"00",
         10063 => x"00",
         10064 => x"00",
         10065 => x"00",
         10066 => x"00",
         10067 => x"00",
         10068 => x"00",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"00",
         10079 => x"00",
         10080 => x"00",
         10081 => x"00",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
         10086 => x"00",
         10087 => x"00",
         10088 => x"00",
         10089 => x"00",
         10090 => x"00",
         10091 => x"00",
         10092 => x"00",
         10093 => x"00",
         10094 => x"00",
         10095 => x"00",
         10096 => x"00",
         10097 => x"00",
         10098 => x"00",
         10099 => x"00",
         10100 => x"00",
         10101 => x"00",
         10102 => x"00",
         10103 => x"00",
         10104 => x"00",
         10105 => x"00",
         10106 => x"00",
         10107 => x"00",
         10108 => x"00",
         10109 => x"00",
         10110 => x"00",
         10111 => x"00",
         10112 => x"00",
         10113 => x"00",
         10114 => x"00",
         10115 => x"00",
         10116 => x"00",
         10117 => x"00",
         10118 => x"00",
         10119 => x"00",
         10120 => x"00",
         10121 => x"00",
         10122 => x"00",
         10123 => x"00",
         10124 => x"00",
         10125 => x"00",
         10126 => x"00",
         10127 => x"00",
         10128 => x"69",
         10129 => x"00",
         10130 => x"69",
         10131 => x"6c",
         10132 => x"69",
         10133 => x"00",
         10134 => x"6c",
         10135 => x"00",
         10136 => x"65",
         10137 => x"00",
         10138 => x"63",
         10139 => x"72",
         10140 => x"63",
         10141 => x"00",
         10142 => x"64",
         10143 => x"00",
         10144 => x"64",
         10145 => x"00",
         10146 => x"65",
         10147 => x"65",
         10148 => x"65",
         10149 => x"69",
         10150 => x"69",
         10151 => x"66",
         10152 => x"66",
         10153 => x"61",
         10154 => x"00",
         10155 => x"6d",
         10156 => x"65",
         10157 => x"72",
         10158 => x"65",
         10159 => x"00",
         10160 => x"6e",
         10161 => x"00",
         10162 => x"62",
         10163 => x"63",
         10164 => x"62",
         10165 => x"63",
         10166 => x"69",
         10167 => x"00",
         10168 => x"64",
         10169 => x"69",
         10170 => x"45",
         10171 => x"72",
         10172 => x"6e",
         10173 => x"6e",
         10174 => x"65",
         10175 => x"72",
         10176 => x"69",
         10177 => x"6e",
         10178 => x"72",
         10179 => x"79",
         10180 => x"6f",
         10181 => x"6c",
         10182 => x"6f",
         10183 => x"2e",
         10184 => x"6f",
         10185 => x"74",
         10186 => x"6f",
         10187 => x"2e",
         10188 => x"6e",
         10189 => x"69",
         10190 => x"69",
         10191 => x"61",
         10192 => x"00",
         10193 => x"63",
         10194 => x"73",
         10195 => x"6e",
         10196 => x"2e",
         10197 => x"69",
         10198 => x"61",
         10199 => x"61",
         10200 => x"65",
         10201 => x"74",
         10202 => x"00",
         10203 => x"69",
         10204 => x"68",
         10205 => x"6c",
         10206 => x"6e",
         10207 => x"69",
         10208 => x"00",
         10209 => x"44",
         10210 => x"20",
         10211 => x"74",
         10212 => x"72",
         10213 => x"63",
         10214 => x"2e",
         10215 => x"72",
         10216 => x"20",
         10217 => x"62",
         10218 => x"69",
         10219 => x"6e",
         10220 => x"69",
         10221 => x"00",
         10222 => x"69",
         10223 => x"6e",
         10224 => x"65",
         10225 => x"6c",
         10226 => x"00",
         10227 => x"6f",
         10228 => x"6d",
         10229 => x"69",
         10230 => x"20",
         10231 => x"65",
         10232 => x"74",
         10233 => x"66",
         10234 => x"64",
         10235 => x"20",
         10236 => x"6b",
         10237 => x"6f",
         10238 => x"74",
         10239 => x"6f",
         10240 => x"64",
         10241 => x"69",
         10242 => x"75",
         10243 => x"6f",
         10244 => x"61",
         10245 => x"6e",
         10246 => x"6e",
         10247 => x"6c",
         10248 => x"00",
         10249 => x"69",
         10250 => x"69",
         10251 => x"6f",
         10252 => x"64",
         10253 => x"6e",
         10254 => x"66",
         10255 => x"65",
         10256 => x"6d",
         10257 => x"72",
         10258 => x"00",
         10259 => x"6f",
         10260 => x"61",
         10261 => x"6f",
         10262 => x"20",
         10263 => x"65",
         10264 => x"00",
         10265 => x"61",
         10266 => x"65",
         10267 => x"73",
         10268 => x"63",
         10269 => x"65",
         10270 => x"00",
         10271 => x"75",
         10272 => x"73",
         10273 => x"00",
         10274 => x"6e",
         10275 => x"77",
         10276 => x"72",
         10277 => x"2e",
         10278 => x"25",
         10279 => x"62",
         10280 => x"73",
         10281 => x"20",
         10282 => x"25",
         10283 => x"62",
         10284 => x"73",
         10285 => x"63",
         10286 => x"00",
         10287 => x"65",
         10288 => x"00",
         10289 => x"30",
         10290 => x"00",
         10291 => x"20",
         10292 => x"30",
         10293 => x"00",
         10294 => x"20",
         10295 => x"20",
         10296 => x"00",
         10297 => x"30",
         10298 => x"00",
         10299 => x"20",
         10300 => x"7c",
         10301 => x"00",
         10302 => x"4f",
         10303 => x"2a",
         10304 => x"20",
         10305 => x"31",
         10306 => x"2f",
         10307 => x"30",
         10308 => x"31",
         10309 => x"00",
         10310 => x"5a",
         10311 => x"20",
         10312 => x"20",
         10313 => x"78",
         10314 => x"73",
         10315 => x"20",
         10316 => x"0a",
         10317 => x"50",
         10318 => x"6e",
         10319 => x"72",
         10320 => x"20",
         10321 => x"64",
         10322 => x"00",
         10323 => x"69",
         10324 => x"20",
         10325 => x"65",
         10326 => x"70",
         10327 => x"53",
         10328 => x"6e",
         10329 => x"72",
         10330 => x"00",
         10331 => x"4f",
         10332 => x"20",
         10333 => x"69",
         10334 => x"72",
         10335 => x"74",
         10336 => x"4f",
         10337 => x"20",
         10338 => x"69",
         10339 => x"72",
         10340 => x"74",
         10341 => x"41",
         10342 => x"20",
         10343 => x"69",
         10344 => x"72",
         10345 => x"74",
         10346 => x"41",
         10347 => x"20",
         10348 => x"69",
         10349 => x"72",
         10350 => x"74",
         10351 => x"41",
         10352 => x"20",
         10353 => x"69",
         10354 => x"72",
         10355 => x"74",
         10356 => x"41",
         10357 => x"20",
         10358 => x"69",
         10359 => x"72",
         10360 => x"74",
         10361 => x"65",
         10362 => x"6e",
         10363 => x"70",
         10364 => x"6d",
         10365 => x"2e",
         10366 => x"6e",
         10367 => x"69",
         10368 => x"74",
         10369 => x"72",
         10370 => x"00",
         10371 => x"75",
         10372 => x"78",
         10373 => x"62",
         10374 => x"00",
         10375 => x"4f",
         10376 => x"70",
         10377 => x"73",
         10378 => x"3a",
         10379 => x"61",
         10380 => x"64",
         10381 => x"20",
         10382 => x"74",
         10383 => x"69",
         10384 => x"73",
         10385 => x"61",
         10386 => x"30",
         10387 => x"6c",
         10388 => x"65",
         10389 => x"69",
         10390 => x"61",
         10391 => x"6c",
         10392 => x"00",
         10393 => x"20",
         10394 => x"6c",
         10395 => x"69",
         10396 => x"2e",
         10397 => x"00",
         10398 => x"6f",
         10399 => x"6e",
         10400 => x"2e",
         10401 => x"6f",
         10402 => x"72",
         10403 => x"2e",
         10404 => x"00",
         10405 => x"30",
         10406 => x"28",
         10407 => x"78",
         10408 => x"25",
         10409 => x"78",
         10410 => x"38",
         10411 => x"00",
         10412 => x"75",
         10413 => x"4d",
         10414 => x"72",
         10415 => x"43",
         10416 => x"6c",
         10417 => x"2e",
         10418 => x"30",
         10419 => x"20",
         10420 => x"58",
         10421 => x"3f",
         10422 => x"30",
         10423 => x"20",
         10424 => x"58",
         10425 => x"30",
         10426 => x"20",
         10427 => x"6c",
         10428 => x"00",
         10429 => x"78",
         10430 => x"74",
         10431 => x"20",
         10432 => x"65",
         10433 => x"25",
         10434 => x"78",
         10435 => x"2e",
         10436 => x"61",
         10437 => x"6e",
         10438 => x"6f",
         10439 => x"40",
         10440 => x"38",
         10441 => x"2e",
         10442 => x"00",
         10443 => x"61",
         10444 => x"72",
         10445 => x"72",
         10446 => x"20",
         10447 => x"65",
         10448 => x"64",
         10449 => x"00",
         10450 => x"65",
         10451 => x"72",
         10452 => x"67",
         10453 => x"70",
         10454 => x"61",
         10455 => x"6e",
         10456 => x"00",
         10457 => x"6f",
         10458 => x"72",
         10459 => x"6f",
         10460 => x"67",
         10461 => x"00",
         10462 => x"50",
         10463 => x"69",
         10464 => x"64",
         10465 => x"73",
         10466 => x"2e",
         10467 => x"00",
         10468 => x"64",
         10469 => x"73",
         10470 => x"00",
         10471 => x"64",
         10472 => x"73",
         10473 => x"61",
         10474 => x"6f",
         10475 => x"6e",
         10476 => x"00",
         10477 => x"65",
         10478 => x"79",
         10479 => x"68",
         10480 => x"74",
         10481 => x"20",
         10482 => x"6e",
         10483 => x"70",
         10484 => x"65",
         10485 => x"63",
         10486 => x"61",
         10487 => x"00",
         10488 => x"75",
         10489 => x"6e",
         10490 => x"2e",
         10491 => x"6e",
         10492 => x"69",
         10493 => x"69",
         10494 => x"72",
         10495 => x"74",
         10496 => x"2e",
         10497 => x"64",
         10498 => x"2f",
         10499 => x"25",
         10500 => x"64",
         10501 => x"2e",
         10502 => x"64",
         10503 => x"6f",
         10504 => x"6f",
         10505 => x"67",
         10506 => x"74",
         10507 => x"00",
         10508 => x"28",
         10509 => x"6d",
         10510 => x"43",
         10511 => x"6e",
         10512 => x"29",
         10513 => x"0a",
         10514 => x"69",
         10515 => x"20",
         10516 => x"6c",
         10517 => x"6e",
         10518 => x"3a",
         10519 => x"20",
         10520 => x"42",
         10521 => x"52",
         10522 => x"20",
         10523 => x"38",
         10524 => x"30",
         10525 => x"2e",
         10526 => x"20",
         10527 => x"44",
         10528 => x"20",
         10529 => x"20",
         10530 => x"38",
         10531 => x"30",
         10532 => x"2e",
         10533 => x"20",
         10534 => x"4e",
         10535 => x"42",
         10536 => x"20",
         10537 => x"38",
         10538 => x"30",
         10539 => x"2e",
         10540 => x"20",
         10541 => x"52",
         10542 => x"20",
         10543 => x"20",
         10544 => x"38",
         10545 => x"30",
         10546 => x"2e",
         10547 => x"20",
         10548 => x"41",
         10549 => x"20",
         10550 => x"20",
         10551 => x"38",
         10552 => x"30",
         10553 => x"2e",
         10554 => x"20",
         10555 => x"44",
         10556 => x"52",
         10557 => x"20",
         10558 => x"76",
         10559 => x"73",
         10560 => x"30",
         10561 => x"2e",
         10562 => x"20",
         10563 => x"49",
         10564 => x"31",
         10565 => x"20",
         10566 => x"6d",
         10567 => x"20",
         10568 => x"30",
         10569 => x"2e",
         10570 => x"20",
         10571 => x"4e",
         10572 => x"43",
         10573 => x"20",
         10574 => x"61",
         10575 => x"6c",
         10576 => x"30",
         10577 => x"2e",
         10578 => x"20",
         10579 => x"49",
         10580 => x"4f",
         10581 => x"42",
         10582 => x"00",
         10583 => x"20",
         10584 => x"42",
         10585 => x"43",
         10586 => x"20",
         10587 => x"4f",
         10588 => x"00",
         10589 => x"20",
         10590 => x"53",
         10591 => x"20",
         10592 => x"50",
         10593 => x"64",
         10594 => x"73",
         10595 => x"3a",
         10596 => x"20",
         10597 => x"50",
         10598 => x"65",
         10599 => x"20",
         10600 => x"74",
         10601 => x"41",
         10602 => x"65",
         10603 => x"3d",
         10604 => x"38",
         10605 => x"00",
         10606 => x"20",
         10607 => x"50",
         10608 => x"65",
         10609 => x"79",
         10610 => x"61",
         10611 => x"41",
         10612 => x"65",
         10613 => x"3d",
         10614 => x"38",
         10615 => x"00",
         10616 => x"20",
         10617 => x"74",
         10618 => x"20",
         10619 => x"72",
         10620 => x"64",
         10621 => x"73",
         10622 => x"20",
         10623 => x"3d",
         10624 => x"38",
         10625 => x"00",
         10626 => x"69",
         10627 => x"00",
         10628 => x"20",
         10629 => x"50",
         10630 => x"64",
         10631 => x"20",
         10632 => x"20",
         10633 => x"20",
         10634 => x"20",
         10635 => x"3d",
         10636 => x"34",
         10637 => x"00",
         10638 => x"20",
         10639 => x"79",
         10640 => x"6d",
         10641 => x"6f",
         10642 => x"46",
         10643 => x"20",
         10644 => x"20",
         10645 => x"3d",
         10646 => x"2e",
         10647 => x"64",
         10648 => x"0a",
         10649 => x"20",
         10650 => x"44",
         10651 => x"20",
         10652 => x"63",
         10653 => x"72",
         10654 => x"20",
         10655 => x"20",
         10656 => x"3d",
         10657 => x"2e",
         10658 => x"64",
         10659 => x"0a",
         10660 => x"20",
         10661 => x"69",
         10662 => x"6f",
         10663 => x"53",
         10664 => x"4d",
         10665 => x"6f",
         10666 => x"46",
         10667 => x"3d",
         10668 => x"2e",
         10669 => x"64",
         10670 => x"0a",
         10671 => x"6d",
         10672 => x"00",
         10673 => x"65",
         10674 => x"6d",
         10675 => x"6c",
         10676 => x"00",
         10677 => x"56",
         10678 => x"56",
         10679 => x"00",
         10680 => x"6e",
         10681 => x"77",
         10682 => x"00",
         10683 => x"00",
         10684 => x"00",
         10685 => x"00",
         10686 => x"00",
         10687 => x"00",
         10688 => x"00",
         10689 => x"00",
         10690 => x"00",
         10691 => x"00",
         10692 => x"00",
         10693 => x"00",
         10694 => x"00",
         10695 => x"00",
         10696 => x"00",
         10697 => x"00",
         10698 => x"00",
         10699 => x"00",
         10700 => x"00",
         10701 => x"00",
         10702 => x"00",
         10703 => x"00",
         10704 => x"00",
         10705 => x"00",
         10706 => x"00",
         10707 => x"00",
         10708 => x"00",
         10709 => x"00",
         10710 => x"00",
         10711 => x"00",
         10712 => x"00",
         10713 => x"00",
         10714 => x"00",
         10715 => x"00",
         10716 => x"00",
         10717 => x"00",
         10718 => x"00",
         10719 => x"00",
         10720 => x"00",
         10721 => x"00",
         10722 => x"00",
         10723 => x"00",
         10724 => x"00",
         10725 => x"00",
         10726 => x"00",
         10727 => x"00",
         10728 => x"00",
         10729 => x"00",
         10730 => x"00",
         10731 => x"00",
         10732 => x"00",
         10733 => x"00",
         10734 => x"00",
         10735 => x"00",
         10736 => x"00",
         10737 => x"00",
         10738 => x"00",
         10739 => x"00",
         10740 => x"00",
         10741 => x"00",
         10742 => x"00",
         10743 => x"00",
         10744 => x"00",
         10745 => x"00",
         10746 => x"00",
         10747 => x"00",
         10748 => x"5b",
         10749 => x"5b",
         10750 => x"5b",
         10751 => x"5b",
         10752 => x"5b",
         10753 => x"5b",
         10754 => x"5b",
         10755 => x"30",
         10756 => x"5b",
         10757 => x"5b",
         10758 => x"5b",
         10759 => x"00",
         10760 => x"00",
         10761 => x"00",
         10762 => x"00",
         10763 => x"00",
         10764 => x"00",
         10765 => x"00",
         10766 => x"00",
         10767 => x"00",
         10768 => x"00",
         10769 => x"00",
         10770 => x"69",
         10771 => x"72",
         10772 => x"69",
         10773 => x"00",
         10774 => x"00",
         10775 => x"30",
         10776 => x"20",
         10777 => x"0a",
         10778 => x"61",
         10779 => x"64",
         10780 => x"20",
         10781 => x"65",
         10782 => x"68",
         10783 => x"69",
         10784 => x"72",
         10785 => x"69",
         10786 => x"74",
         10787 => x"4f",
         10788 => x"00",
         10789 => x"61",
         10790 => x"74",
         10791 => x"65",
         10792 => x"72",
         10793 => x"65",
         10794 => x"73",
         10795 => x"79",
         10796 => x"6c",
         10797 => x"64",
         10798 => x"62",
         10799 => x"67",
         10800 => x"44",
         10801 => x"2a",
         10802 => x"3f",
         10803 => x"00",
         10804 => x"2c",
         10805 => x"5d",
         10806 => x"41",
         10807 => x"41",
         10808 => x"00",
         10809 => x"fe",
         10810 => x"44",
         10811 => x"2e",
         10812 => x"4f",
         10813 => x"4d",
         10814 => x"20",
         10815 => x"54",
         10816 => x"20",
         10817 => x"4f",
         10818 => x"4d",
         10819 => x"20",
         10820 => x"54",
         10821 => x"20",
         10822 => x"00",
         10823 => x"00",
         10824 => x"00",
         10825 => x"00",
         10826 => x"03",
         10827 => x"0e",
         10828 => x"16",
         10829 => x"00",
         10830 => x"9a",
         10831 => x"41",
         10832 => x"45",
         10833 => x"49",
         10834 => x"92",
         10835 => x"4f",
         10836 => x"99",
         10837 => x"9d",
         10838 => x"49",
         10839 => x"a5",
         10840 => x"a9",
         10841 => x"ad",
         10842 => x"b1",
         10843 => x"b5",
         10844 => x"b9",
         10845 => x"bd",
         10846 => x"c1",
         10847 => x"c5",
         10848 => x"c9",
         10849 => x"cd",
         10850 => x"d1",
         10851 => x"d5",
         10852 => x"d9",
         10853 => x"dd",
         10854 => x"e1",
         10855 => x"e5",
         10856 => x"e9",
         10857 => x"ed",
         10858 => x"f1",
         10859 => x"f5",
         10860 => x"f9",
         10861 => x"fd",
         10862 => x"2e",
         10863 => x"5b",
         10864 => x"22",
         10865 => x"3e",
         10866 => x"00",
         10867 => x"01",
         10868 => x"10",
         10869 => x"00",
         10870 => x"00",
         10871 => x"01",
         10872 => x"04",
         10873 => x"10",
         10874 => x"00",
         10875 => x"c7",
         10876 => x"e9",
         10877 => x"e4",
         10878 => x"e5",
         10879 => x"ea",
         10880 => x"e8",
         10881 => x"ee",
         10882 => x"c4",
         10883 => x"c9",
         10884 => x"c6",
         10885 => x"f6",
         10886 => x"fb",
         10887 => x"ff",
         10888 => x"dc",
         10889 => x"a3",
         10890 => x"a7",
         10891 => x"e1",
         10892 => x"f3",
         10893 => x"f1",
         10894 => x"aa",
         10895 => x"bf",
         10896 => x"ac",
         10897 => x"bc",
         10898 => x"ab",
         10899 => x"91",
         10900 => x"93",
         10901 => x"24",
         10902 => x"62",
         10903 => x"55",
         10904 => x"51",
         10905 => x"5d",
         10906 => x"5b",
         10907 => x"14",
         10908 => x"2c",
         10909 => x"00",
         10910 => x"5e",
         10911 => x"5a",
         10912 => x"69",
         10913 => x"60",
         10914 => x"6c",
         10915 => x"68",
         10916 => x"65",
         10917 => x"58",
         10918 => x"53",
         10919 => x"6a",
         10920 => x"0c",
         10921 => x"84",
         10922 => x"90",
         10923 => x"b1",
         10924 => x"93",
         10925 => x"a3",
         10926 => x"b5",
         10927 => x"a6",
         10928 => x"a9",
         10929 => x"1e",
         10930 => x"b5",
         10931 => x"61",
         10932 => x"65",
         10933 => x"20",
         10934 => x"f7",
         10935 => x"b0",
         10936 => x"b7",
         10937 => x"7f",
         10938 => x"a0",
         10939 => x"61",
         10940 => x"e0",
         10941 => x"f8",
         10942 => x"ff",
         10943 => x"78",
         10944 => x"30",
         10945 => x"06",
         10946 => x"10",
         10947 => x"2e",
         10948 => x"06",
         10949 => x"4d",
         10950 => x"81",
         10951 => x"82",
         10952 => x"84",
         10953 => x"87",
         10954 => x"89",
         10955 => x"8b",
         10956 => x"8d",
         10957 => x"8f",
         10958 => x"91",
         10959 => x"93",
         10960 => x"f6",
         10961 => x"97",
         10962 => x"98",
         10963 => x"9b",
         10964 => x"9d",
         10965 => x"9f",
         10966 => x"a0",
         10967 => x"a2",
         10968 => x"a4",
         10969 => x"a7",
         10970 => x"a9",
         10971 => x"ab",
         10972 => x"ac",
         10973 => x"af",
         10974 => x"b1",
         10975 => x"b3",
         10976 => x"b5",
         10977 => x"b7",
         10978 => x"b8",
         10979 => x"bb",
         10980 => x"bc",
         10981 => x"f7",
         10982 => x"c1",
         10983 => x"c3",
         10984 => x"c5",
         10985 => x"c7",
         10986 => x"c7",
         10987 => x"cb",
         10988 => x"cd",
         10989 => x"dd",
         10990 => x"8e",
         10991 => x"12",
         10992 => x"03",
         10993 => x"f4",
         10994 => x"f8",
         10995 => x"22",
         10996 => x"3a",
         10997 => x"65",
         10998 => x"3b",
         10999 => x"66",
         11000 => x"40",
         11001 => x"41",
         11002 => x"0a",
         11003 => x"40",
         11004 => x"86",
         11005 => x"89",
         11006 => x"58",
         11007 => x"5a",
         11008 => x"5c",
         11009 => x"5e",
         11010 => x"93",
         11011 => x"62",
         11012 => x"64",
         11013 => x"66",
         11014 => x"97",
         11015 => x"6a",
         11016 => x"6c",
         11017 => x"6e",
         11018 => x"70",
         11019 => x"9d",
         11020 => x"74",
         11021 => x"76",
         11022 => x"78",
         11023 => x"7a",
         11024 => x"7c",
         11025 => x"7e",
         11026 => x"a6",
         11027 => x"82",
         11028 => x"84",
         11029 => x"86",
         11030 => x"ae",
         11031 => x"b1",
         11032 => x"45",
         11033 => x"8e",
         11034 => x"90",
         11035 => x"b7",
         11036 => x"03",
         11037 => x"fe",
         11038 => x"ac",
         11039 => x"86",
         11040 => x"89",
         11041 => x"b1",
         11042 => x"c2",
         11043 => x"a3",
         11044 => x"c4",
         11045 => x"cc",
         11046 => x"8c",
         11047 => x"8f",
         11048 => x"18",
         11049 => x"0a",
         11050 => x"f3",
         11051 => x"f5",
         11052 => x"f7",
         11053 => x"f9",
         11054 => x"fa",
         11055 => x"20",
         11056 => x"10",
         11057 => x"22",
         11058 => x"36",
         11059 => x"0e",
         11060 => x"01",
         11061 => x"d0",
         11062 => x"61",
         11063 => x"00",
         11064 => x"7d",
         11065 => x"63",
         11066 => x"96",
         11067 => x"5a",
         11068 => x"08",
         11069 => x"06",
         11070 => x"08",
         11071 => x"08",
         11072 => x"06",
         11073 => x"07",
         11074 => x"52",
         11075 => x"54",
         11076 => x"56",
         11077 => x"60",
         11078 => x"70",
         11079 => x"ba",
         11080 => x"c8",
         11081 => x"ca",
         11082 => x"da",
         11083 => x"f8",
         11084 => x"ea",
         11085 => x"fa",
         11086 => x"80",
         11087 => x"90",
         11088 => x"a0",
         11089 => x"b0",
         11090 => x"b8",
         11091 => x"b2",
         11092 => x"cc",
         11093 => x"c3",
         11094 => x"02",
         11095 => x"02",
         11096 => x"01",
         11097 => x"f3",
         11098 => x"fc",
         11099 => x"01",
         11100 => x"70",
         11101 => x"84",
         11102 => x"83",
         11103 => x"1a",
         11104 => x"2f",
         11105 => x"02",
         11106 => x"06",
         11107 => x"02",
         11108 => x"64",
         11109 => x"26",
         11110 => x"1a",
         11111 => x"00",
         11112 => x"00",
         11113 => x"02",
         11114 => x"00",
         11115 => x"00",
         11116 => x"00",
         11117 => x"04",
         11118 => x"00",
         11119 => x"00",
         11120 => x"00",
         11121 => x"14",
         11122 => x"00",
         11123 => x"00",
         11124 => x"00",
         11125 => x"2b",
         11126 => x"00",
         11127 => x"00",
         11128 => x"00",
         11129 => x"30",
         11130 => x"00",
         11131 => x"00",
         11132 => x"00",
         11133 => x"3c",
         11134 => x"00",
         11135 => x"00",
         11136 => x"00",
         11137 => x"3d",
         11138 => x"00",
         11139 => x"00",
         11140 => x"00",
         11141 => x"3f",
         11142 => x"00",
         11143 => x"00",
         11144 => x"00",
         11145 => x"40",
         11146 => x"00",
         11147 => x"00",
         11148 => x"00",
         11149 => x"41",
         11150 => x"00",
         11151 => x"00",
         11152 => x"00",
         11153 => x"42",
         11154 => x"00",
         11155 => x"00",
         11156 => x"00",
         11157 => x"43",
         11158 => x"00",
         11159 => x"00",
         11160 => x"00",
         11161 => x"50",
         11162 => x"00",
         11163 => x"00",
         11164 => x"00",
         11165 => x"51",
         11166 => x"00",
         11167 => x"00",
         11168 => x"00",
         11169 => x"54",
         11170 => x"00",
         11171 => x"00",
         11172 => x"00",
         11173 => x"55",
         11174 => x"00",
         11175 => x"00",
         11176 => x"00",
         11177 => x"79",
         11178 => x"00",
         11179 => x"00",
         11180 => x"00",
         11181 => x"78",
         11182 => x"00",
         11183 => x"00",
         11184 => x"00",
         11185 => x"82",
         11186 => x"00",
         11187 => x"00",
         11188 => x"00",
         11189 => x"83",
         11190 => x"00",
         11191 => x"00",
         11192 => x"00",
         11193 => x"85",
         11194 => x"00",
         11195 => x"00",
         11196 => x"00",
         11197 => x"8c",
         11198 => x"00",
         11199 => x"00",
         11200 => x"00",
         11201 => x"8d",
         11202 => x"00",
         11203 => x"00",
         11204 => x"00",
         11205 => x"8e",
         11206 => x"00",
         11207 => x"00",
         11208 => x"00",
         11209 => x"8f",
         11210 => x"00",
         11211 => x"00",
         11212 => x"00",
         11213 => x"00",
         11214 => x"00",
         11215 => x"00",
         11216 => x"00",
         11217 => x"01",
         11218 => x"00",
         11219 => x"01",
         11220 => x"81",
         11221 => x"00",
         11222 => x"7f",
         11223 => x"00",
         11224 => x"00",
         11225 => x"00",
         11226 => x"00",
         11227 => x"f5",
         11228 => x"f5",
         11229 => x"f5",
         11230 => x"00",
         11231 => x"01",
         11232 => x"01",
         11233 => x"01",
         11234 => x"00",
         11235 => x"00",
         11236 => x"00",
         11237 => x"00",
         11238 => x"00",
         11239 => x"00",
         11240 => x"00",
         11241 => x"00",
         11242 => x"00",
         11243 => x"00",
         11244 => x"00",
         11245 => x"00",
         11246 => x"00",
         11247 => x"00",
         11248 => x"00",
         11249 => x"00",
         11250 => x"00",
         11251 => x"00",
         11252 => x"00",
         11253 => x"00",
         11254 => x"00",
         11255 => x"00",
         11256 => x"00",
         11257 => x"00",
         11258 => x"00",
         11259 => x"00",
         11260 => x"00",
         11261 => x"00",
         11262 => x"00",
         11263 => x"00",
         11264 => x"00",
         11265 => x"00",
         11266 => x"00",
         11267 => x"01",
         11268 => x"03",
         11269 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"f8",
             2 => x"0b",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"d1",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"ec",
           163 => x"10",
           164 => x"06",
           165 => x"93",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"fe",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"fc",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"ff",
           252 => x"ff",
           253 => x"ff",
           254 => x"ff",
           255 => x"ff",
           256 => x"00",
           257 => x"ff",
           258 => x"ff",
           259 => x"ff",
           260 => x"ff",
           261 => x"ff",
           262 => x"ff",
           263 => x"ff",
           264 => x"0b",
           265 => x"81",
           266 => x"0b",
           267 => x"0b",
           268 => x"96",
           269 => x"0b",
           270 => x"0b",
           271 => x"b6",
           272 => x"0b",
           273 => x"0b",
           274 => x"d6",
           275 => x"0b",
           276 => x"0b",
           277 => x"f7",
           278 => x"0b",
           279 => x"0b",
           280 => x"98",
           281 => x"0b",
           282 => x"0b",
           283 => x"b8",
           284 => x"0b",
           285 => x"0b",
           286 => x"da",
           287 => x"0b",
           288 => x"0b",
           289 => x"fc",
           290 => x"0b",
           291 => x"0b",
           292 => x"9e",
           293 => x"0b",
           294 => x"0b",
           295 => x"c0",
           296 => x"0b",
           297 => x"0b",
           298 => x"e2",
           299 => x"0b",
           300 => x"0b",
           301 => x"84",
           302 => x"0b",
           303 => x"0b",
           304 => x"a6",
           305 => x"0b",
           306 => x"0b",
           307 => x"c8",
           308 => x"0b",
           309 => x"0b",
           310 => x"ea",
           311 => x"0b",
           312 => x"0b",
           313 => x"8c",
           314 => x"0b",
           315 => x"0b",
           316 => x"ae",
           317 => x"0b",
           318 => x"0b",
           319 => x"d0",
           320 => x"0b",
           321 => x"0b",
           322 => x"f2",
           323 => x"0b",
           324 => x"0b",
           325 => x"94",
           326 => x"0b",
           327 => x"0b",
           328 => x"b6",
           329 => x"0b",
           330 => x"0b",
           331 => x"d8",
           332 => x"0b",
           333 => x"0b",
           334 => x"fa",
           335 => x"0b",
           336 => x"0b",
           337 => x"9c",
           338 => x"0b",
           339 => x"0b",
           340 => x"be",
           341 => x"0b",
           342 => x"0b",
           343 => x"e0",
           344 => x"0b",
           345 => x"0b",
           346 => x"82",
           347 => x"ff",
           348 => x"ff",
           349 => x"ff",
           350 => x"ff",
           351 => x"ff",
           352 => x"ff",
           353 => x"ff",
           354 => x"ff",
           355 => x"ff",
           356 => x"ff",
           357 => x"ff",
           358 => x"ff",
           359 => x"ff",
           360 => x"ff",
           361 => x"ff",
           362 => x"ff",
           363 => x"ff",
           364 => x"ff",
           365 => x"ff",
           366 => x"ff",
           367 => x"ff",
           368 => x"ff",
           369 => x"ff",
           370 => x"ff",
           371 => x"ff",
           372 => x"ff",
           373 => x"ff",
           374 => x"ff",
           375 => x"ff",
           376 => x"ff",
           377 => x"ff",
           378 => x"ff",
           379 => x"ff",
           380 => x"ff",
           381 => x"ff",
           382 => x"ff",
           383 => x"ff",
           384 => x"04",
           385 => x"04",
           386 => x"0c",
           387 => x"2d",
           388 => x"08",
           389 => x"90",
           390 => x"a4",
           391 => x"2d",
           392 => x"08",
           393 => x"90",
           394 => x"a4",
           395 => x"2d",
           396 => x"08",
           397 => x"90",
           398 => x"a4",
           399 => x"2d",
           400 => x"08",
           401 => x"90",
           402 => x"a4",
           403 => x"2d",
           404 => x"08",
           405 => x"90",
           406 => x"a4",
           407 => x"2d",
           408 => x"08",
           409 => x"90",
           410 => x"a4",
           411 => x"9f",
           412 => x"a4",
           413 => x"80",
           414 => x"e0",
           415 => x"d4",
           416 => x"e0",
           417 => x"c0",
           418 => x"82",
           419 => x"94",
           420 => x"e0",
           421 => x"c0",
           422 => x"82",
           423 => x"96",
           424 => x"e0",
           425 => x"c0",
           426 => x"82",
           427 => x"98",
           428 => x"e0",
           429 => x"c0",
           430 => x"82",
           431 => x"80",
           432 => x"82",
           433 => x"80",
           434 => x"04",
           435 => x"0c",
           436 => x"2d",
           437 => x"08",
           438 => x"90",
           439 => x"a4",
           440 => x"dd",
           441 => x"a4",
           442 => x"80",
           443 => x"e0",
           444 => x"fd",
           445 => x"e0",
           446 => x"c0",
           447 => x"82",
           448 => x"80",
           449 => x"82",
           450 => x"80",
           451 => x"04",
           452 => x"0c",
           453 => x"2d",
           454 => x"08",
           455 => x"90",
           456 => x"a4",
           457 => x"a7",
           458 => x"a4",
           459 => x"80",
           460 => x"e0",
           461 => x"fb",
           462 => x"e0",
           463 => x"c0",
           464 => x"82",
           465 => x"81",
           466 => x"82",
           467 => x"80",
           468 => x"04",
           469 => x"0c",
           470 => x"2d",
           471 => x"08",
           472 => x"90",
           473 => x"a4",
           474 => x"ce",
           475 => x"a4",
           476 => x"80",
           477 => x"e0",
           478 => x"82",
           479 => x"e0",
           480 => x"c0",
           481 => x"82",
           482 => x"82",
           483 => x"82",
           484 => x"80",
           485 => x"04",
           486 => x"0c",
           487 => x"2d",
           488 => x"08",
           489 => x"90",
           490 => x"a4",
           491 => x"c7",
           492 => x"a4",
           493 => x"80",
           494 => x"e0",
           495 => x"95",
           496 => x"e0",
           497 => x"c0",
           498 => x"82",
           499 => x"82",
           500 => x"82",
           501 => x"80",
           502 => x"04",
           503 => x"0c",
           504 => x"2d",
           505 => x"08",
           506 => x"90",
           507 => x"a4",
           508 => x"cd",
           509 => x"a4",
           510 => x"80",
           511 => x"e0",
           512 => x"9b",
           513 => x"e0",
           514 => x"c0",
           515 => x"82",
           516 => x"82",
           517 => x"82",
           518 => x"80",
           519 => x"04",
           520 => x"0c",
           521 => x"2d",
           522 => x"08",
           523 => x"90",
           524 => x"a4",
           525 => x"e0",
           526 => x"a4",
           527 => x"80",
           528 => x"e0",
           529 => x"85",
           530 => x"e0",
           531 => x"c0",
           532 => x"82",
           533 => x"82",
           534 => x"82",
           535 => x"80",
           536 => x"04",
           537 => x"0c",
           538 => x"2d",
           539 => x"08",
           540 => x"90",
           541 => x"a4",
           542 => x"99",
           543 => x"a4",
           544 => x"80",
           545 => x"e0",
           546 => x"a2",
           547 => x"e0",
           548 => x"c0",
           549 => x"82",
           550 => x"81",
           551 => x"82",
           552 => x"80",
           553 => x"04",
           554 => x"0c",
           555 => x"2d",
           556 => x"08",
           557 => x"90",
           558 => x"a4",
           559 => x"e9",
           560 => x"a4",
           561 => x"80",
           562 => x"e0",
           563 => x"b2",
           564 => x"e0",
           565 => x"c0",
           566 => x"82",
           567 => x"81",
           568 => x"82",
           569 => x"80",
           570 => x"04",
           571 => x"0c",
           572 => x"2d",
           573 => x"08",
           574 => x"90",
           575 => x"a4",
           576 => x"d9",
           577 => x"a4",
           578 => x"80",
           579 => x"e0",
           580 => x"fb",
           581 => x"e0",
           582 => x"c0",
           583 => x"82",
           584 => x"80",
           585 => x"82",
           586 => x"80",
           587 => x"04",
           588 => x"0c",
           589 => x"2d",
           590 => x"08",
           591 => x"90",
           592 => x"a4",
           593 => x"ef",
           594 => x"a4",
           595 => x"80",
           596 => x"e0",
           597 => x"af",
           598 => x"e0",
           599 => x"c0",
           600 => x"82",
           601 => x"81",
           602 => x"82",
           603 => x"80",
           604 => x"04",
           605 => x"0c",
           606 => x"2d",
           607 => x"08",
           608 => x"90",
           609 => x"a4",
           610 => x"89",
           611 => x"a4",
           612 => x"80",
           613 => x"04",
           614 => x"10",
           615 => x"10",
           616 => x"10",
           617 => x"10",
           618 => x"10",
           619 => x"10",
           620 => x"10",
           621 => x"53",
           622 => x"00",
           623 => x"06",
           624 => x"09",
           625 => x"05",
           626 => x"2b",
           627 => x"06",
           628 => x"04",
           629 => x"72",
           630 => x"05",
           631 => x"05",
           632 => x"72",
           633 => x"53",
           634 => x"51",
           635 => x"04",
           636 => x"70",
           637 => x"27",
           638 => x"71",
           639 => x"53",
           640 => x"0b",
           641 => x"8c",
           642 => x"fa",
           643 => x"82",
           644 => x"02",
           645 => x"0c",
           646 => x"82",
           647 => x"8c",
           648 => x"e0",
           649 => x"05",
           650 => x"a4",
           651 => x"08",
           652 => x"a4",
           653 => x"08",
           654 => x"fc",
           655 => x"84",
           656 => x"e0",
           657 => x"82",
           658 => x"f8",
           659 => x"e0",
           660 => x"05",
           661 => x"e0",
           662 => x"54",
           663 => x"82",
           664 => x"04",
           665 => x"08",
           666 => x"a4",
           667 => x"0d",
           668 => x"08",
           669 => x"85",
           670 => x"81",
           671 => x"06",
           672 => x"52",
           673 => x"80",
           674 => x"a4",
           675 => x"08",
           676 => x"8d",
           677 => x"82",
           678 => x"f4",
           679 => x"c4",
           680 => x"a4",
           681 => x"08",
           682 => x"e0",
           683 => x"05",
           684 => x"82",
           685 => x"f8",
           686 => x"e0",
           687 => x"05",
           688 => x"a4",
           689 => x"0c",
           690 => x"08",
           691 => x"8a",
           692 => x"38",
           693 => x"e0",
           694 => x"05",
           695 => x"e9",
           696 => x"a4",
           697 => x"08",
           698 => x"3f",
           699 => x"08",
           700 => x"a4",
           701 => x"0c",
           702 => x"a4",
           703 => x"08",
           704 => x"81",
           705 => x"80",
           706 => x"a4",
           707 => x"0c",
           708 => x"82",
           709 => x"fc",
           710 => x"e0",
           711 => x"05",
           712 => x"71",
           713 => x"e0",
           714 => x"05",
           715 => x"82",
           716 => x"8c",
           717 => x"e0",
           718 => x"05",
           719 => x"82",
           720 => x"fc",
           721 => x"80",
           722 => x"a4",
           723 => x"08",
           724 => x"34",
           725 => x"08",
           726 => x"70",
           727 => x"08",
           728 => x"52",
           729 => x"08",
           730 => x"82",
           731 => x"87",
           732 => x"e0",
           733 => x"82",
           734 => x"02",
           735 => x"0c",
           736 => x"86",
           737 => x"a4",
           738 => x"34",
           739 => x"08",
           740 => x"82",
           741 => x"e0",
           742 => x"0a",
           743 => x"a4",
           744 => x"0c",
           745 => x"08",
           746 => x"82",
           747 => x"fc",
           748 => x"e0",
           749 => x"05",
           750 => x"e0",
           751 => x"05",
           752 => x"e0",
           753 => x"05",
           754 => x"54",
           755 => x"82",
           756 => x"70",
           757 => x"08",
           758 => x"82",
           759 => x"ec",
           760 => x"e0",
           761 => x"05",
           762 => x"54",
           763 => x"82",
           764 => x"dc",
           765 => x"82",
           766 => x"54",
           767 => x"82",
           768 => x"04",
           769 => x"08",
           770 => x"a4",
           771 => x"0d",
           772 => x"08",
           773 => x"82",
           774 => x"fc",
           775 => x"e0",
           776 => x"05",
           777 => x"e0",
           778 => x"05",
           779 => x"e0",
           780 => x"05",
           781 => x"a3",
           782 => x"98",
           783 => x"e0",
           784 => x"05",
           785 => x"a4",
           786 => x"08",
           787 => x"98",
           788 => x"87",
           789 => x"e0",
           790 => x"82",
           791 => x"02",
           792 => x"0c",
           793 => x"80",
           794 => x"a4",
           795 => x"23",
           796 => x"08",
           797 => x"53",
           798 => x"14",
           799 => x"a4",
           800 => x"08",
           801 => x"70",
           802 => x"81",
           803 => x"06",
           804 => x"51",
           805 => x"2e",
           806 => x"0b",
           807 => x"08",
           808 => x"96",
           809 => x"e0",
           810 => x"05",
           811 => x"33",
           812 => x"e0",
           813 => x"05",
           814 => x"ff",
           815 => x"80",
           816 => x"38",
           817 => x"08",
           818 => x"81",
           819 => x"a4",
           820 => x"0c",
           821 => x"08",
           822 => x"70",
           823 => x"53",
           824 => x"95",
           825 => x"e0",
           826 => x"05",
           827 => x"73",
           828 => x"38",
           829 => x"08",
           830 => x"53",
           831 => x"81",
           832 => x"e0",
           833 => x"05",
           834 => x"b0",
           835 => x"06",
           836 => x"82",
           837 => x"e8",
           838 => x"98",
           839 => x"2c",
           840 => x"72",
           841 => x"e0",
           842 => x"05",
           843 => x"2a",
           844 => x"70",
           845 => x"51",
           846 => x"80",
           847 => x"82",
           848 => x"e4",
           849 => x"82",
           850 => x"53",
           851 => x"a4",
           852 => x"23",
           853 => x"82",
           854 => x"e8",
           855 => x"98",
           856 => x"2c",
           857 => x"2b",
           858 => x"11",
           859 => x"53",
           860 => x"72",
           861 => x"08",
           862 => x"82",
           863 => x"e8",
           864 => x"82",
           865 => x"f8",
           866 => x"15",
           867 => x"51",
           868 => x"e0",
           869 => x"05",
           870 => x"a4",
           871 => x"33",
           872 => x"70",
           873 => x"51",
           874 => x"25",
           875 => x"ff",
           876 => x"a4",
           877 => x"34",
           878 => x"08",
           879 => x"70",
           880 => x"81",
           881 => x"53",
           882 => x"38",
           883 => x"08",
           884 => x"70",
           885 => x"90",
           886 => x"2c",
           887 => x"51",
           888 => x"53",
           889 => x"a4",
           890 => x"23",
           891 => x"82",
           892 => x"e4",
           893 => x"83",
           894 => x"06",
           895 => x"72",
           896 => x"38",
           897 => x"08",
           898 => x"70",
           899 => x"98",
           900 => x"53",
           901 => x"81",
           902 => x"a4",
           903 => x"34",
           904 => x"08",
           905 => x"e0",
           906 => x"a4",
           907 => x"0c",
           908 => x"a4",
           909 => x"08",
           910 => x"92",
           911 => x"e0",
           912 => x"05",
           913 => x"2b",
           914 => x"11",
           915 => x"51",
           916 => x"04",
           917 => x"08",
           918 => x"70",
           919 => x"53",
           920 => x"a4",
           921 => x"23",
           922 => x"08",
           923 => x"70",
           924 => x"53",
           925 => x"a4",
           926 => x"23",
           927 => x"82",
           928 => x"e4",
           929 => x"81",
           930 => x"53",
           931 => x"a4",
           932 => x"23",
           933 => x"82",
           934 => x"e4",
           935 => x"80",
           936 => x"53",
           937 => x"a4",
           938 => x"23",
           939 => x"82",
           940 => x"e4",
           941 => x"88",
           942 => x"72",
           943 => x"08",
           944 => x"80",
           945 => x"a4",
           946 => x"34",
           947 => x"82",
           948 => x"e4",
           949 => x"84",
           950 => x"72",
           951 => x"08",
           952 => x"fb",
           953 => x"0b",
           954 => x"08",
           955 => x"82",
           956 => x"ec",
           957 => x"11",
           958 => x"82",
           959 => x"ec",
           960 => x"e3",
           961 => x"a4",
           962 => x"34",
           963 => x"82",
           964 => x"90",
           965 => x"e0",
           966 => x"05",
           967 => x"82",
           968 => x"90",
           969 => x"08",
           970 => x"82",
           971 => x"fc",
           972 => x"e0",
           973 => x"05",
           974 => x"51",
           975 => x"e0",
           976 => x"05",
           977 => x"39",
           978 => x"08",
           979 => x"82",
           980 => x"90",
           981 => x"05",
           982 => x"08",
           983 => x"70",
           984 => x"a4",
           985 => x"0c",
           986 => x"08",
           987 => x"70",
           988 => x"81",
           989 => x"51",
           990 => x"2e",
           991 => x"e0",
           992 => x"05",
           993 => x"2b",
           994 => x"2c",
           995 => x"a4",
           996 => x"08",
           997 => x"83",
           998 => x"98",
           999 => x"82",
          1000 => x"f4",
          1001 => x"39",
          1002 => x"08",
          1003 => x"51",
          1004 => x"82",
          1005 => x"53",
          1006 => x"a4",
          1007 => x"23",
          1008 => x"08",
          1009 => x"53",
          1010 => x"08",
          1011 => x"73",
          1012 => x"54",
          1013 => x"a4",
          1014 => x"23",
          1015 => x"82",
          1016 => x"90",
          1017 => x"e0",
          1018 => x"05",
          1019 => x"82",
          1020 => x"90",
          1021 => x"08",
          1022 => x"08",
          1023 => x"82",
          1024 => x"e4",
          1025 => x"83",
          1026 => x"06",
          1027 => x"53",
          1028 => x"ab",
          1029 => x"a4",
          1030 => x"33",
          1031 => x"53",
          1032 => x"53",
          1033 => x"08",
          1034 => x"52",
          1035 => x"3f",
          1036 => x"08",
          1037 => x"e0",
          1038 => x"05",
          1039 => x"82",
          1040 => x"fc",
          1041 => x"9b",
          1042 => x"e0",
          1043 => x"72",
          1044 => x"08",
          1045 => x"82",
          1046 => x"ec",
          1047 => x"82",
          1048 => x"f4",
          1049 => x"71",
          1050 => x"72",
          1051 => x"08",
          1052 => x"8a",
          1053 => x"e0",
          1054 => x"05",
          1055 => x"2a",
          1056 => x"51",
          1057 => x"80",
          1058 => x"82",
          1059 => x"90",
          1060 => x"e0",
          1061 => x"05",
          1062 => x"82",
          1063 => x"90",
          1064 => x"08",
          1065 => x"08",
          1066 => x"53",
          1067 => x"e0",
          1068 => x"05",
          1069 => x"a4",
          1070 => x"08",
          1071 => x"e0",
          1072 => x"05",
          1073 => x"82",
          1074 => x"dc",
          1075 => x"82",
          1076 => x"dc",
          1077 => x"e0",
          1078 => x"05",
          1079 => x"a4",
          1080 => x"08",
          1081 => x"38",
          1082 => x"08",
          1083 => x"70",
          1084 => x"53",
          1085 => x"a4",
          1086 => x"23",
          1087 => x"08",
          1088 => x"30",
          1089 => x"08",
          1090 => x"82",
          1091 => x"e4",
          1092 => x"ff",
          1093 => x"53",
          1094 => x"a4",
          1095 => x"23",
          1096 => x"88",
          1097 => x"a4",
          1098 => x"23",
          1099 => x"e0",
          1100 => x"05",
          1101 => x"c0",
          1102 => x"72",
          1103 => x"08",
          1104 => x"80",
          1105 => x"e0",
          1106 => x"05",
          1107 => x"82",
          1108 => x"f4",
          1109 => x"e0",
          1110 => x"05",
          1111 => x"2a",
          1112 => x"51",
          1113 => x"80",
          1114 => x"82",
          1115 => x"90",
          1116 => x"e0",
          1117 => x"05",
          1118 => x"82",
          1119 => x"90",
          1120 => x"08",
          1121 => x"08",
          1122 => x"53",
          1123 => x"e0",
          1124 => x"05",
          1125 => x"a4",
          1126 => x"08",
          1127 => x"e0",
          1128 => x"05",
          1129 => x"82",
          1130 => x"d8",
          1131 => x"82",
          1132 => x"d8",
          1133 => x"e0",
          1134 => x"05",
          1135 => x"a4",
          1136 => x"22",
          1137 => x"51",
          1138 => x"e0",
          1139 => x"05",
          1140 => x"a8",
          1141 => x"a4",
          1142 => x"0c",
          1143 => x"08",
          1144 => x"82",
          1145 => x"f4",
          1146 => x"e0",
          1147 => x"05",
          1148 => x"70",
          1149 => x"55",
          1150 => x"82",
          1151 => x"53",
          1152 => x"82",
          1153 => x"f0",
          1154 => x"e0",
          1155 => x"05",
          1156 => x"a4",
          1157 => x"08",
          1158 => x"53",
          1159 => x"a4",
          1160 => x"a4",
          1161 => x"08",
          1162 => x"54",
          1163 => x"08",
          1164 => x"70",
          1165 => x"51",
          1166 => x"82",
          1167 => x"d0",
          1168 => x"39",
          1169 => x"08",
          1170 => x"53",
          1171 => x"11",
          1172 => x"82",
          1173 => x"d0",
          1174 => x"e0",
          1175 => x"05",
          1176 => x"e0",
          1177 => x"05",
          1178 => x"82",
          1179 => x"f0",
          1180 => x"05",
          1181 => x"08",
          1182 => x"82",
          1183 => x"f4",
          1184 => x"53",
          1185 => x"08",
          1186 => x"52",
          1187 => x"3f",
          1188 => x"08",
          1189 => x"a4",
          1190 => x"0c",
          1191 => x"a4",
          1192 => x"08",
          1193 => x"38",
          1194 => x"82",
          1195 => x"f0",
          1196 => x"e0",
          1197 => x"72",
          1198 => x"75",
          1199 => x"72",
          1200 => x"08",
          1201 => x"82",
          1202 => x"e4",
          1203 => x"b2",
          1204 => x"72",
          1205 => x"38",
          1206 => x"08",
          1207 => x"ff",
          1208 => x"72",
          1209 => x"08",
          1210 => x"82",
          1211 => x"e4",
          1212 => x"86",
          1213 => x"06",
          1214 => x"72",
          1215 => x"e7",
          1216 => x"a4",
          1217 => x"22",
          1218 => x"82",
          1219 => x"cc",
          1220 => x"e0",
          1221 => x"05",
          1222 => x"82",
          1223 => x"cc",
          1224 => x"e0",
          1225 => x"05",
          1226 => x"72",
          1227 => x"81",
          1228 => x"82",
          1229 => x"cc",
          1230 => x"05",
          1231 => x"e0",
          1232 => x"05",
          1233 => x"82",
          1234 => x"cc",
          1235 => x"05",
          1236 => x"e0",
          1237 => x"05",
          1238 => x"a4",
          1239 => x"22",
          1240 => x"08",
          1241 => x"82",
          1242 => x"e4",
          1243 => x"83",
          1244 => x"06",
          1245 => x"72",
          1246 => x"d0",
          1247 => x"a4",
          1248 => x"33",
          1249 => x"70",
          1250 => x"e0",
          1251 => x"05",
          1252 => x"51",
          1253 => x"24",
          1254 => x"e0",
          1255 => x"05",
          1256 => x"06",
          1257 => x"82",
          1258 => x"e4",
          1259 => x"39",
          1260 => x"08",
          1261 => x"53",
          1262 => x"08",
          1263 => x"73",
          1264 => x"54",
          1265 => x"a4",
          1266 => x"34",
          1267 => x"08",
          1268 => x"70",
          1269 => x"81",
          1270 => x"53",
          1271 => x"b1",
          1272 => x"a4",
          1273 => x"33",
          1274 => x"70",
          1275 => x"90",
          1276 => x"2c",
          1277 => x"51",
          1278 => x"82",
          1279 => x"ec",
          1280 => x"75",
          1281 => x"72",
          1282 => x"08",
          1283 => x"af",
          1284 => x"a4",
          1285 => x"33",
          1286 => x"70",
          1287 => x"90",
          1288 => x"2c",
          1289 => x"51",
          1290 => x"82",
          1291 => x"ec",
          1292 => x"75",
          1293 => x"72",
          1294 => x"08",
          1295 => x"82",
          1296 => x"e4",
          1297 => x"83",
          1298 => x"53",
          1299 => x"82",
          1300 => x"ec",
          1301 => x"11",
          1302 => x"82",
          1303 => x"ec",
          1304 => x"90",
          1305 => x"2c",
          1306 => x"73",
          1307 => x"82",
          1308 => x"88",
          1309 => x"a0",
          1310 => x"3f",
          1311 => x"e0",
          1312 => x"05",
          1313 => x"2a",
          1314 => x"51",
          1315 => x"80",
          1316 => x"82",
          1317 => x"88",
          1318 => x"ad",
          1319 => x"3f",
          1320 => x"82",
          1321 => x"e4",
          1322 => x"84",
          1323 => x"06",
          1324 => x"72",
          1325 => x"38",
          1326 => x"08",
          1327 => x"52",
          1328 => x"a5",
          1329 => x"82",
          1330 => x"e4",
          1331 => x"85",
          1332 => x"06",
          1333 => x"72",
          1334 => x"38",
          1335 => x"08",
          1336 => x"52",
          1337 => x"81",
          1338 => x"a4",
          1339 => x"22",
          1340 => x"70",
          1341 => x"51",
          1342 => x"2e",
          1343 => x"e0",
          1344 => x"05",
          1345 => x"51",
          1346 => x"82",
          1347 => x"f4",
          1348 => x"72",
          1349 => x"81",
          1350 => x"82",
          1351 => x"88",
          1352 => x"82",
          1353 => x"f8",
          1354 => x"89",
          1355 => x"e0",
          1356 => x"05",
          1357 => x"2a",
          1358 => x"51",
          1359 => x"80",
          1360 => x"82",
          1361 => x"ec",
          1362 => x"11",
          1363 => x"82",
          1364 => x"ec",
          1365 => x"90",
          1366 => x"2c",
          1367 => x"73",
          1368 => x"82",
          1369 => x"88",
          1370 => x"b0",
          1371 => x"3f",
          1372 => x"e0",
          1373 => x"05",
          1374 => x"2a",
          1375 => x"51",
          1376 => x"80",
          1377 => x"82",
          1378 => x"e8",
          1379 => x"11",
          1380 => x"82",
          1381 => x"e8",
          1382 => x"98",
          1383 => x"2c",
          1384 => x"73",
          1385 => x"82",
          1386 => x"88",
          1387 => x"b0",
          1388 => x"3f",
          1389 => x"e0",
          1390 => x"05",
          1391 => x"2a",
          1392 => x"51",
          1393 => x"b0",
          1394 => x"a4",
          1395 => x"22",
          1396 => x"54",
          1397 => x"a4",
          1398 => x"23",
          1399 => x"70",
          1400 => x"53",
          1401 => x"90",
          1402 => x"a4",
          1403 => x"08",
          1404 => x"87",
          1405 => x"39",
          1406 => x"08",
          1407 => x"53",
          1408 => x"2e",
          1409 => x"97",
          1410 => x"a4",
          1411 => x"08",
          1412 => x"a4",
          1413 => x"33",
          1414 => x"3f",
          1415 => x"82",
          1416 => x"f8",
          1417 => x"72",
          1418 => x"09",
          1419 => x"cb",
          1420 => x"a4",
          1421 => x"22",
          1422 => x"53",
          1423 => x"a4",
          1424 => x"23",
          1425 => x"ff",
          1426 => x"83",
          1427 => x"81",
          1428 => x"e0",
          1429 => x"05",
          1430 => x"e0",
          1431 => x"05",
          1432 => x"52",
          1433 => x"08",
          1434 => x"81",
          1435 => x"a4",
          1436 => x"0c",
          1437 => x"3f",
          1438 => x"82",
          1439 => x"f8",
          1440 => x"72",
          1441 => x"09",
          1442 => x"cb",
          1443 => x"a4",
          1444 => x"22",
          1445 => x"53",
          1446 => x"a4",
          1447 => x"23",
          1448 => x"ff",
          1449 => x"83",
          1450 => x"80",
          1451 => x"e0",
          1452 => x"05",
          1453 => x"e0",
          1454 => x"05",
          1455 => x"52",
          1456 => x"3f",
          1457 => x"08",
          1458 => x"81",
          1459 => x"a4",
          1460 => x"0c",
          1461 => x"82",
          1462 => x"f0",
          1463 => x"e0",
          1464 => x"38",
          1465 => x"08",
          1466 => x"52",
          1467 => x"08",
          1468 => x"ff",
          1469 => x"a4",
          1470 => x"0c",
          1471 => x"08",
          1472 => x"70",
          1473 => x"85",
          1474 => x"39",
          1475 => x"08",
          1476 => x"70",
          1477 => x"81",
          1478 => x"53",
          1479 => x"80",
          1480 => x"e0",
          1481 => x"05",
          1482 => x"54",
          1483 => x"e0",
          1484 => x"05",
          1485 => x"2b",
          1486 => x"51",
          1487 => x"25",
          1488 => x"e0",
          1489 => x"05",
          1490 => x"51",
          1491 => x"d2",
          1492 => x"a4",
          1493 => x"08",
          1494 => x"a4",
          1495 => x"33",
          1496 => x"3f",
          1497 => x"e0",
          1498 => x"05",
          1499 => x"39",
          1500 => x"08",
          1501 => x"53",
          1502 => x"09",
          1503 => x"38",
          1504 => x"e0",
          1505 => x"05",
          1506 => x"82",
          1507 => x"ec",
          1508 => x"0b",
          1509 => x"08",
          1510 => x"8a",
          1511 => x"a4",
          1512 => x"23",
          1513 => x"82",
          1514 => x"88",
          1515 => x"82",
          1516 => x"f8",
          1517 => x"84",
          1518 => x"ea",
          1519 => x"a4",
          1520 => x"08",
          1521 => x"70",
          1522 => x"08",
          1523 => x"51",
          1524 => x"a4",
          1525 => x"08",
          1526 => x"0c",
          1527 => x"82",
          1528 => x"04",
          1529 => x"08",
          1530 => x"a4",
          1531 => x"0d",
          1532 => x"08",
          1533 => x"a4",
          1534 => x"08",
          1535 => x"a4",
          1536 => x"08",
          1537 => x"3f",
          1538 => x"08",
          1539 => x"98",
          1540 => x"3d",
          1541 => x"a4",
          1542 => x"e0",
          1543 => x"82",
          1544 => x"fb",
          1545 => x"0b",
          1546 => x"08",
          1547 => x"82",
          1548 => x"85",
          1549 => x"81",
          1550 => x"32",
          1551 => x"51",
          1552 => x"53",
          1553 => x"8d",
          1554 => x"82",
          1555 => x"f4",
          1556 => x"92",
          1557 => x"a4",
          1558 => x"08",
          1559 => x"82",
          1560 => x"88",
          1561 => x"05",
          1562 => x"08",
          1563 => x"53",
          1564 => x"a4",
          1565 => x"34",
          1566 => x"06",
          1567 => x"2e",
          1568 => x"fb",
          1569 => x"fb",
          1570 => x"82",
          1571 => x"fc",
          1572 => x"90",
          1573 => x"53",
          1574 => x"e0",
          1575 => x"72",
          1576 => x"b1",
          1577 => x"82",
          1578 => x"f8",
          1579 => x"a5",
          1580 => x"fc",
          1581 => x"fc",
          1582 => x"8a",
          1583 => x"08",
          1584 => x"82",
          1585 => x"53",
          1586 => x"8a",
          1587 => x"82",
          1588 => x"f8",
          1589 => x"e0",
          1590 => x"05",
          1591 => x"e0",
          1592 => x"05",
          1593 => x"e0",
          1594 => x"05",
          1595 => x"98",
          1596 => x"0d",
          1597 => x"0c",
          1598 => x"a4",
          1599 => x"e0",
          1600 => x"3d",
          1601 => x"82",
          1602 => x"f8",
          1603 => x"e0",
          1604 => x"05",
          1605 => x"33",
          1606 => x"70",
          1607 => x"81",
          1608 => x"51",
          1609 => x"80",
          1610 => x"ff",
          1611 => x"a4",
          1612 => x"0c",
          1613 => x"82",
          1614 => x"88",
          1615 => x"72",
          1616 => x"a4",
          1617 => x"08",
          1618 => x"e0",
          1619 => x"05",
          1620 => x"82",
          1621 => x"fc",
          1622 => x"81",
          1623 => x"72",
          1624 => x"38",
          1625 => x"08",
          1626 => x"82",
          1627 => x"8c",
          1628 => x"82",
          1629 => x"fc",
          1630 => x"90",
          1631 => x"53",
          1632 => x"e0",
          1633 => x"72",
          1634 => x"ab",
          1635 => x"82",
          1636 => x"f8",
          1637 => x"9f",
          1638 => x"a4",
          1639 => x"08",
          1640 => x"a4",
          1641 => x"0c",
          1642 => x"a4",
          1643 => x"08",
          1644 => x"0c",
          1645 => x"82",
          1646 => x"04",
          1647 => x"08",
          1648 => x"a4",
          1649 => x"0d",
          1650 => x"08",
          1651 => x"a4",
          1652 => x"08",
          1653 => x"82",
          1654 => x"70",
          1655 => x"0c",
          1656 => x"0d",
          1657 => x"0c",
          1658 => x"a4",
          1659 => x"e0",
          1660 => x"3d",
          1661 => x"a4",
          1662 => x"08",
          1663 => x"70",
          1664 => x"81",
          1665 => x"06",
          1666 => x"51",
          1667 => x"2e",
          1668 => x"0b",
          1669 => x"08",
          1670 => x"81",
          1671 => x"e0",
          1672 => x"05",
          1673 => x"33",
          1674 => x"70",
          1675 => x"51",
          1676 => x"80",
          1677 => x"38",
          1678 => x"08",
          1679 => x"82",
          1680 => x"8c",
          1681 => x"54",
          1682 => x"88",
          1683 => x"9f",
          1684 => x"a4",
          1685 => x"08",
          1686 => x"82",
          1687 => x"88",
          1688 => x"57",
          1689 => x"75",
          1690 => x"81",
          1691 => x"82",
          1692 => x"8c",
          1693 => x"11",
          1694 => x"8c",
          1695 => x"e0",
          1696 => x"05",
          1697 => x"e0",
          1698 => x"05",
          1699 => x"80",
          1700 => x"e0",
          1701 => x"05",
          1702 => x"a4",
          1703 => x"08",
          1704 => x"a4",
          1705 => x"08",
          1706 => x"06",
          1707 => x"08",
          1708 => x"72",
          1709 => x"98",
          1710 => x"a3",
          1711 => x"a4",
          1712 => x"08",
          1713 => x"81",
          1714 => x"0c",
          1715 => x"08",
          1716 => x"70",
          1717 => x"08",
          1718 => x"51",
          1719 => x"ff",
          1720 => x"a4",
          1721 => x"0c",
          1722 => x"08",
          1723 => x"82",
          1724 => x"87",
          1725 => x"e0",
          1726 => x"82",
          1727 => x"02",
          1728 => x"0c",
          1729 => x"82",
          1730 => x"88",
          1731 => x"11",
          1732 => x"32",
          1733 => x"51",
          1734 => x"71",
          1735 => x"38",
          1736 => x"e0",
          1737 => x"05",
          1738 => x"39",
          1739 => x"08",
          1740 => x"85",
          1741 => x"86",
          1742 => x"06",
          1743 => x"52",
          1744 => x"80",
          1745 => x"e0",
          1746 => x"05",
          1747 => x"a4",
          1748 => x"08",
          1749 => x"12",
          1750 => x"bf",
          1751 => x"71",
          1752 => x"82",
          1753 => x"88",
          1754 => x"11",
          1755 => x"8c",
          1756 => x"e0",
          1757 => x"05",
          1758 => x"33",
          1759 => x"a4",
          1760 => x"0c",
          1761 => x"82",
          1762 => x"e0",
          1763 => x"05",
          1764 => x"33",
          1765 => x"70",
          1766 => x"51",
          1767 => x"80",
          1768 => x"38",
          1769 => x"08",
          1770 => x"70",
          1771 => x"82",
          1772 => x"fc",
          1773 => x"52",
          1774 => x"08",
          1775 => x"a9",
          1776 => x"a4",
          1777 => x"08",
          1778 => x"08",
          1779 => x"53",
          1780 => x"33",
          1781 => x"51",
          1782 => x"14",
          1783 => x"82",
          1784 => x"f8",
          1785 => x"d7",
          1786 => x"a4",
          1787 => x"08",
          1788 => x"05",
          1789 => x"81",
          1790 => x"e0",
          1791 => x"05",
          1792 => x"a4",
          1793 => x"08",
          1794 => x"08",
          1795 => x"2d",
          1796 => x"08",
          1797 => x"a4",
          1798 => x"0c",
          1799 => x"a4",
          1800 => x"08",
          1801 => x"f2",
          1802 => x"a4",
          1803 => x"08",
          1804 => x"08",
          1805 => x"82",
          1806 => x"88",
          1807 => x"11",
          1808 => x"a4",
          1809 => x"0c",
          1810 => x"a4",
          1811 => x"08",
          1812 => x"81",
          1813 => x"82",
          1814 => x"f0",
          1815 => x"07",
          1816 => x"e0",
          1817 => x"05",
          1818 => x"82",
          1819 => x"f0",
          1820 => x"07",
          1821 => x"e0",
          1822 => x"05",
          1823 => x"a4",
          1824 => x"08",
          1825 => x"a4",
          1826 => x"33",
          1827 => x"ff",
          1828 => x"a4",
          1829 => x"0c",
          1830 => x"e0",
          1831 => x"05",
          1832 => x"08",
          1833 => x"12",
          1834 => x"a4",
          1835 => x"08",
          1836 => x"06",
          1837 => x"a4",
          1838 => x"0c",
          1839 => x"82",
          1840 => x"f8",
          1841 => x"e0",
          1842 => x"3d",
          1843 => x"a4",
          1844 => x"e0",
          1845 => x"82",
          1846 => x"fd",
          1847 => x"e0",
          1848 => x"05",
          1849 => x"a4",
          1850 => x"0c",
          1851 => x"08",
          1852 => x"82",
          1853 => x"f8",
          1854 => x"e0",
          1855 => x"05",
          1856 => x"82",
          1857 => x"e0",
          1858 => x"05",
          1859 => x"a4",
          1860 => x"08",
          1861 => x"38",
          1862 => x"08",
          1863 => x"82",
          1864 => x"90",
          1865 => x"51",
          1866 => x"08",
          1867 => x"71",
          1868 => x"38",
          1869 => x"08",
          1870 => x"82",
          1871 => x"90",
          1872 => x"82",
          1873 => x"fc",
          1874 => x"e0",
          1875 => x"05",
          1876 => x"a4",
          1877 => x"08",
          1878 => x"a4",
          1879 => x"0c",
          1880 => x"08",
          1881 => x"81",
          1882 => x"a4",
          1883 => x"0c",
          1884 => x"08",
          1885 => x"ff",
          1886 => x"a4",
          1887 => x"0c",
          1888 => x"08",
          1889 => x"80",
          1890 => x"38",
          1891 => x"08",
          1892 => x"ff",
          1893 => x"a4",
          1894 => x"0c",
          1895 => x"08",
          1896 => x"ff",
          1897 => x"a4",
          1898 => x"0c",
          1899 => x"08",
          1900 => x"82",
          1901 => x"f8",
          1902 => x"51",
          1903 => x"34",
          1904 => x"82",
          1905 => x"90",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"90",
          1910 => x"05",
          1911 => x"08",
          1912 => x"82",
          1913 => x"90",
          1914 => x"2e",
          1915 => x"e0",
          1916 => x"05",
          1917 => x"33",
          1918 => x"08",
          1919 => x"81",
          1920 => x"a4",
          1921 => x"0c",
          1922 => x"08",
          1923 => x"52",
          1924 => x"34",
          1925 => x"08",
          1926 => x"81",
          1927 => x"a4",
          1928 => x"0c",
          1929 => x"82",
          1930 => x"88",
          1931 => x"82",
          1932 => x"51",
          1933 => x"82",
          1934 => x"04",
          1935 => x"08",
          1936 => x"a4",
          1937 => x"0d",
          1938 => x"08",
          1939 => x"82",
          1940 => x"fc",
          1941 => x"e0",
          1942 => x"05",
          1943 => x"33",
          1944 => x"08",
          1945 => x"81",
          1946 => x"a4",
          1947 => x"0c",
          1948 => x"06",
          1949 => x"80",
          1950 => x"da",
          1951 => x"a4",
          1952 => x"08",
          1953 => x"e0",
          1954 => x"05",
          1955 => x"a4",
          1956 => x"08",
          1957 => x"08",
          1958 => x"31",
          1959 => x"98",
          1960 => x"3d",
          1961 => x"a4",
          1962 => x"e0",
          1963 => x"82",
          1964 => x"fe",
          1965 => x"e0",
          1966 => x"05",
          1967 => x"a4",
          1968 => x"0c",
          1969 => x"08",
          1970 => x"52",
          1971 => x"e0",
          1972 => x"05",
          1973 => x"82",
          1974 => x"8c",
          1975 => x"e0",
          1976 => x"05",
          1977 => x"70",
          1978 => x"e0",
          1979 => x"05",
          1980 => x"82",
          1981 => x"fc",
          1982 => x"81",
          1983 => x"70",
          1984 => x"38",
          1985 => x"82",
          1986 => x"88",
          1987 => x"82",
          1988 => x"51",
          1989 => x"82",
          1990 => x"04",
          1991 => x"08",
          1992 => x"a4",
          1993 => x"0d",
          1994 => x"08",
          1995 => x"82",
          1996 => x"fc",
          1997 => x"e0",
          1998 => x"05",
          1999 => x"a4",
          2000 => x"0c",
          2001 => x"08",
          2002 => x"80",
          2003 => x"38",
          2004 => x"08",
          2005 => x"81",
          2006 => x"a4",
          2007 => x"0c",
          2008 => x"08",
          2009 => x"ff",
          2010 => x"a4",
          2011 => x"0c",
          2012 => x"08",
          2013 => x"80",
          2014 => x"82",
          2015 => x"f8",
          2016 => x"70",
          2017 => x"a4",
          2018 => x"08",
          2019 => x"e0",
          2020 => x"05",
          2021 => x"a4",
          2022 => x"08",
          2023 => x"71",
          2024 => x"a4",
          2025 => x"08",
          2026 => x"e0",
          2027 => x"05",
          2028 => x"39",
          2029 => x"08",
          2030 => x"70",
          2031 => x"0c",
          2032 => x"0d",
          2033 => x"0c",
          2034 => x"a4",
          2035 => x"e0",
          2036 => x"3d",
          2037 => x"a4",
          2038 => x"08",
          2039 => x"f4",
          2040 => x"a4",
          2041 => x"08",
          2042 => x"82",
          2043 => x"8c",
          2044 => x"05",
          2045 => x"08",
          2046 => x"82",
          2047 => x"88",
          2048 => x"33",
          2049 => x"06",
          2050 => x"51",
          2051 => x"84",
          2052 => x"39",
          2053 => x"08",
          2054 => x"52",
          2055 => x"e0",
          2056 => x"05",
          2057 => x"82",
          2058 => x"88",
          2059 => x"81",
          2060 => x"51",
          2061 => x"80",
          2062 => x"a4",
          2063 => x"0c",
          2064 => x"82",
          2065 => x"90",
          2066 => x"05",
          2067 => x"08",
          2068 => x"82",
          2069 => x"90",
          2070 => x"2e",
          2071 => x"81",
          2072 => x"a4",
          2073 => x"08",
          2074 => x"e8",
          2075 => x"a4",
          2076 => x"08",
          2077 => x"53",
          2078 => x"ff",
          2079 => x"a4",
          2080 => x"0c",
          2081 => x"82",
          2082 => x"8c",
          2083 => x"05",
          2084 => x"08",
          2085 => x"82",
          2086 => x"8c",
          2087 => x"33",
          2088 => x"8c",
          2089 => x"82",
          2090 => x"fc",
          2091 => x"39",
          2092 => x"08",
          2093 => x"70",
          2094 => x"a4",
          2095 => x"08",
          2096 => x"71",
          2097 => x"e0",
          2098 => x"05",
          2099 => x"52",
          2100 => x"39",
          2101 => x"e0",
          2102 => x"05",
          2103 => x"a4",
          2104 => x"08",
          2105 => x"0c",
          2106 => x"82",
          2107 => x"04",
          2108 => x"08",
          2109 => x"a4",
          2110 => x"0d",
          2111 => x"08",
          2112 => x"52",
          2113 => x"08",
          2114 => x"51",
          2115 => x"82",
          2116 => x"70",
          2117 => x"08",
          2118 => x"82",
          2119 => x"f8",
          2120 => x"05",
          2121 => x"54",
          2122 => x"3f",
          2123 => x"08",
          2124 => x"a4",
          2125 => x"0c",
          2126 => x"a4",
          2127 => x"08",
          2128 => x"0b",
          2129 => x"08",
          2130 => x"bc",
          2131 => x"a4",
          2132 => x"08",
          2133 => x"08",
          2134 => x"05",
          2135 => x"34",
          2136 => x"08",
          2137 => x"53",
          2138 => x"08",
          2139 => x"52",
          2140 => x"08",
          2141 => x"51",
          2142 => x"82",
          2143 => x"70",
          2144 => x"08",
          2145 => x"54",
          2146 => x"08",
          2147 => x"82",
          2148 => x"88",
          2149 => x"e0",
          2150 => x"82",
          2151 => x"02",
          2152 => x"0c",
          2153 => x"82",
          2154 => x"88",
          2155 => x"e0",
          2156 => x"05",
          2157 => x"a4",
          2158 => x"08",
          2159 => x"0b",
          2160 => x"08",
          2161 => x"80",
          2162 => x"e0",
          2163 => x"05",
          2164 => x"33",
          2165 => x"08",
          2166 => x"81",
          2167 => x"a4",
          2168 => x"0c",
          2169 => x"06",
          2170 => x"80",
          2171 => x"82",
          2172 => x"8c",
          2173 => x"05",
          2174 => x"08",
          2175 => x"82",
          2176 => x"8c",
          2177 => x"2e",
          2178 => x"be",
          2179 => x"a4",
          2180 => x"08",
          2181 => x"e0",
          2182 => x"05",
          2183 => x"a4",
          2184 => x"08",
          2185 => x"08",
          2186 => x"31",
          2187 => x"a4",
          2188 => x"0c",
          2189 => x"a4",
          2190 => x"08",
          2191 => x"0c",
          2192 => x"82",
          2193 => x"04",
          2194 => x"08",
          2195 => x"a4",
          2196 => x"0d",
          2197 => x"08",
          2198 => x"82",
          2199 => x"fc",
          2200 => x"e0",
          2201 => x"05",
          2202 => x"80",
          2203 => x"e0",
          2204 => x"05",
          2205 => x"82",
          2206 => x"90",
          2207 => x"e0",
          2208 => x"05",
          2209 => x"82",
          2210 => x"90",
          2211 => x"e0",
          2212 => x"05",
          2213 => x"a9",
          2214 => x"a4",
          2215 => x"08",
          2216 => x"e0",
          2217 => x"05",
          2218 => x"71",
          2219 => x"e0",
          2220 => x"05",
          2221 => x"82",
          2222 => x"fc",
          2223 => x"be",
          2224 => x"a4",
          2225 => x"08",
          2226 => x"98",
          2227 => x"3d",
          2228 => x"a4",
          2229 => x"e0",
          2230 => x"82",
          2231 => x"fe",
          2232 => x"e0",
          2233 => x"05",
          2234 => x"e0",
          2235 => x"05",
          2236 => x"3f",
          2237 => x"08",
          2238 => x"98",
          2239 => x"3d",
          2240 => x"a4",
          2241 => x"e0",
          2242 => x"82",
          2243 => x"f6",
          2244 => x"0b",
          2245 => x"08",
          2246 => x"82",
          2247 => x"8c",
          2248 => x"2e",
          2249 => x"e0",
          2250 => x"05",
          2251 => x"fc",
          2252 => x"98",
          2253 => x"e0",
          2254 => x"05",
          2255 => x"39",
          2256 => x"08",
          2257 => x"82",
          2258 => x"e4",
          2259 => x"e0",
          2260 => x"05",
          2261 => x"a3",
          2262 => x"a4",
          2263 => x"08",
          2264 => x"3f",
          2265 => x"08",
          2266 => x"08",
          2267 => x"71",
          2268 => x"a4",
          2269 => x"0c",
          2270 => x"82",
          2271 => x"e4",
          2272 => x"e0",
          2273 => x"05",
          2274 => x"e0",
          2275 => x"05",
          2276 => x"a4",
          2277 => x"08",
          2278 => x"08",
          2279 => x"82",
          2280 => x"fc",
          2281 => x"05",
          2282 => x"e0",
          2283 => x"05",
          2284 => x"38",
          2285 => x"e0",
          2286 => x"05",
          2287 => x"39",
          2288 => x"08",
          2289 => x"ff",
          2290 => x"82",
          2291 => x"f8",
          2292 => x"09",
          2293 => x"38",
          2294 => x"08",
          2295 => x"70",
          2296 => x"08",
          2297 => x"52",
          2298 => x"82",
          2299 => x"f8",
          2300 => x"05",
          2301 => x"08",
          2302 => x"82",
          2303 => x"88",
          2304 => x"e0",
          2305 => x"05",
          2306 => x"e0",
          2307 => x"05",
          2308 => x"a4",
          2309 => x"08",
          2310 => x"08",
          2311 => x"31",
          2312 => x"08",
          2313 => x"71",
          2314 => x"a4",
          2315 => x"0c",
          2316 => x"82",
          2317 => x"f0",
          2318 => x"e0",
          2319 => x"05",
          2320 => x"81",
          2321 => x"e0",
          2322 => x"05",
          2323 => x"e0",
          2324 => x"05",
          2325 => x"82",
          2326 => x"88",
          2327 => x"2a",
          2328 => x"82",
          2329 => x"f4",
          2330 => x"e0",
          2331 => x"05",
          2332 => x"82",
          2333 => x"f0",
          2334 => x"82",
          2335 => x"88",
          2336 => x"e0",
          2337 => x"05",
          2338 => x"a4",
          2339 => x"08",
          2340 => x"82",
          2341 => x"fc",
          2342 => x"05",
          2343 => x"82",
          2344 => x"ec",
          2345 => x"e0",
          2346 => x"05",
          2347 => x"82",
          2348 => x"f0",
          2349 => x"e0",
          2350 => x"05",
          2351 => x"a4",
          2352 => x"08",
          2353 => x"a4",
          2354 => x"08",
          2355 => x"e0",
          2356 => x"05",
          2357 => x"a4",
          2358 => x"08",
          2359 => x"e0",
          2360 => x"05",
          2361 => x"55",
          2362 => x"53",
          2363 => x"39",
          2364 => x"08",
          2365 => x"10",
          2366 => x"a4",
          2367 => x"08",
          2368 => x"a4",
          2369 => x"0c",
          2370 => x"08",
          2371 => x"70",
          2372 => x"08",
          2373 => x"51",
          2374 => x"a4",
          2375 => x"08",
          2376 => x"0c",
          2377 => x"82",
          2378 => x"04",
          2379 => x"08",
          2380 => x"a4",
          2381 => x"0d",
          2382 => x"08",
          2383 => x"82",
          2384 => x"fc",
          2385 => x"e0",
          2386 => x"05",
          2387 => x"80",
          2388 => x"8c",
          2389 => x"82",
          2390 => x"f0",
          2391 => x"39",
          2392 => x"e0",
          2393 => x"05",
          2394 => x"a4",
          2395 => x"08",
          2396 => x"08",
          2397 => x"90",
          2398 => x"a4",
          2399 => x"08",
          2400 => x"a4",
          2401 => x"08",
          2402 => x"e0",
          2403 => x"05",
          2404 => x"a4",
          2405 => x"08",
          2406 => x"08",
          2407 => x"82",
          2408 => x"fc",
          2409 => x"fe",
          2410 => x"51",
          2411 => x"88",
          2412 => x"a4",
          2413 => x"0c",
          2414 => x"0b",
          2415 => x"08",
          2416 => x"82",
          2417 => x"ec",
          2418 => x"e0",
          2419 => x"05",
          2420 => x"82",
          2421 => x"f8",
          2422 => x"82",
          2423 => x"fc",
          2424 => x"2a",
          2425 => x"08",
          2426 => x"82",
          2427 => x"f4",
          2428 => x"e0",
          2429 => x"05",
          2430 => x"e0",
          2431 => x"05",
          2432 => x"a4",
          2433 => x"08",
          2434 => x"51",
          2435 => x"38",
          2436 => x"e0",
          2437 => x"05",
          2438 => x"80",
          2439 => x"a4",
          2440 => x"0c",
          2441 => x"08",
          2442 => x"82",
          2443 => x"f8",
          2444 => x"0b",
          2445 => x"08",
          2446 => x"31",
          2447 => x"08",
          2448 => x"71",
          2449 => x"a4",
          2450 => x"0c",
          2451 => x"08",
          2452 => x"82",
          2453 => x"f8",
          2454 => x"82",
          2455 => x"f4",
          2456 => x"e0",
          2457 => x"05",
          2458 => x"51",
          2459 => x"38",
          2460 => x"e0",
          2461 => x"05",
          2462 => x"80",
          2463 => x"a4",
          2464 => x"0c",
          2465 => x"08",
          2466 => x"82",
          2467 => x"f8",
          2468 => x"0b",
          2469 => x"08",
          2470 => x"31",
          2471 => x"08",
          2472 => x"71",
          2473 => x"a4",
          2474 => x"0c",
          2475 => x"08",
          2476 => x"82",
          2477 => x"f8",
          2478 => x"82",
          2479 => x"f4",
          2480 => x"0b",
          2481 => x"08",
          2482 => x"31",
          2483 => x"08",
          2484 => x"81",
          2485 => x"32",
          2486 => x"70",
          2487 => x"06",
          2488 => x"08",
          2489 => x"11",
          2490 => x"e0",
          2491 => x"51",
          2492 => x"51",
          2493 => x"8a",
          2494 => x"e0",
          2495 => x"82",
          2496 => x"02",
          2497 => x"0c",
          2498 => x"82",
          2499 => x"8c",
          2500 => x"82",
          2501 => x"88",
          2502 => x"84",
          2503 => x"e0",
          2504 => x"82",
          2505 => x"8c",
          2506 => x"82",
          2507 => x"88",
          2508 => x"31",
          2509 => x"98",
          2510 => x"53",
          2511 => x"82",
          2512 => x"04",
          2513 => x"08",
          2514 => x"a4",
          2515 => x"0d",
          2516 => x"08",
          2517 => x"52",
          2518 => x"08",
          2519 => x"51",
          2520 => x"e0",
          2521 => x"82",
          2522 => x"53",
          2523 => x"82",
          2524 => x"04",
          2525 => x"08",
          2526 => x"a4",
          2527 => x"0d",
          2528 => x"e0",
          2529 => x"05",
          2530 => x"a4",
          2531 => x"08",
          2532 => x"38",
          2533 => x"08",
          2534 => x"51",
          2535 => x"82",
          2536 => x"70",
          2537 => x"08",
          2538 => x"52",
          2539 => x"e0",
          2540 => x"05",
          2541 => x"a4",
          2542 => x"0c",
          2543 => x"08",
          2544 => x"80",
          2545 => x"82",
          2546 => x"88",
          2547 => x"fa",
          2548 => x"e0",
          2549 => x"e0",
          2550 => x"05",
          2551 => x"82",
          2552 => x"e0",
          2553 => x"97",
          2554 => x"a4",
          2555 => x"08",
          2556 => x"08",
          2557 => x"31",
          2558 => x"08",
          2559 => x"82",
          2560 => x"e0",
          2561 => x"e0",
          2562 => x"05",
          2563 => x"a4",
          2564 => x"08",
          2565 => x"71",
          2566 => x"08",
          2567 => x"27",
          2568 => x"e0",
          2569 => x"05",
          2570 => x"e0",
          2571 => x"05",
          2572 => x"ba",
          2573 => x"a4",
          2574 => x"08",
          2575 => x"71",
          2576 => x"08",
          2577 => x"2e",
          2578 => x"8d",
          2579 => x"82",
          2580 => x"e8",
          2581 => x"96",
          2582 => x"a4",
          2583 => x"08",
          2584 => x"e0",
          2585 => x"05",
          2586 => x"a4",
          2587 => x"08",
          2588 => x"08",
          2589 => x"2a",
          2590 => x"08",
          2591 => x"82",
          2592 => x"fc",
          2593 => x"e0",
          2594 => x"05",
          2595 => x"e0",
          2596 => x"05",
          2597 => x"82",
          2598 => x"88",
          2599 => x"80",
          2600 => x"a4",
          2601 => x"0c",
          2602 => x"08",
          2603 => x"80",
          2604 => x"38",
          2605 => x"08",
          2606 => x"10",
          2607 => x"08",
          2608 => x"ff",
          2609 => x"a4",
          2610 => x"08",
          2611 => x"73",
          2612 => x"a4",
          2613 => x"0c",
          2614 => x"08",
          2615 => x"10",
          2616 => x"a4",
          2617 => x"08",
          2618 => x"a4",
          2619 => x"0c",
          2620 => x"08",
          2621 => x"82",
          2622 => x"f4",
          2623 => x"ff",
          2624 => x"a4",
          2625 => x"08",
          2626 => x"71",
          2627 => x"a4",
          2628 => x"0c",
          2629 => x"08",
          2630 => x"81",
          2631 => x"a4",
          2632 => x"0c",
          2633 => x"08",
          2634 => x"82",
          2635 => x"ec",
          2636 => x"82",
          2637 => x"f4",
          2638 => x"31",
          2639 => x"08",
          2640 => x"82",
          2641 => x"f8",
          2642 => x"05",
          2643 => x"08",
          2644 => x"51",
          2645 => x"51",
          2646 => x"fe",
          2647 => x"e0",
          2648 => x"05",
          2649 => x"e0",
          2650 => x"05",
          2651 => x"e0",
          2652 => x"05",
          2653 => x"98",
          2654 => x"0d",
          2655 => x"0c",
          2656 => x"a4",
          2657 => x"e0",
          2658 => x"3d",
          2659 => x"82",
          2660 => x"fc",
          2661 => x"e0",
          2662 => x"05",
          2663 => x"a4",
          2664 => x"08",
          2665 => x"a4",
          2666 => x"0c",
          2667 => x"08",
          2668 => x"82",
          2669 => x"fc",
          2670 => x"82",
          2671 => x"f4",
          2672 => x"e0",
          2673 => x"05",
          2674 => x"a4",
          2675 => x"08",
          2676 => x"e0",
          2677 => x"05",
          2678 => x"e0",
          2679 => x"05",
          2680 => x"a4",
          2681 => x"08",
          2682 => x"08",
          2683 => x"32",
          2684 => x"a4",
          2685 => x"08",
          2686 => x"a4",
          2687 => x"0c",
          2688 => x"08",
          2689 => x"82",
          2690 => x"f4",
          2691 => x"82",
          2692 => x"f8",
          2693 => x"e0",
          2694 => x"05",
          2695 => x"e0",
          2696 => x"05",
          2697 => x"53",
          2698 => x"82",
          2699 => x"70",
          2700 => x"08",
          2701 => x"32",
          2702 => x"a4",
          2703 => x"08",
          2704 => x"e0",
          2705 => x"51",
          2706 => x"0d",
          2707 => x"0c",
          2708 => x"a4",
          2709 => x"e0",
          2710 => x"3d",
          2711 => x"82",
          2712 => x"f0",
          2713 => x"e0",
          2714 => x"05",
          2715 => x"73",
          2716 => x"a4",
          2717 => x"08",
          2718 => x"53",
          2719 => x"72",
          2720 => x"08",
          2721 => x"72",
          2722 => x"53",
          2723 => x"09",
          2724 => x"38",
          2725 => x"08",
          2726 => x"70",
          2727 => x"71",
          2728 => x"39",
          2729 => x"08",
          2730 => x"53",
          2731 => x"09",
          2732 => x"38",
          2733 => x"e0",
          2734 => x"05",
          2735 => x"a4",
          2736 => x"08",
          2737 => x"05",
          2738 => x"08",
          2739 => x"33",
          2740 => x"08",
          2741 => x"82",
          2742 => x"f8",
          2743 => x"72",
          2744 => x"81",
          2745 => x"38",
          2746 => x"08",
          2747 => x"70",
          2748 => x"71",
          2749 => x"51",
          2750 => x"82",
          2751 => x"f8",
          2752 => x"e0",
          2753 => x"05",
          2754 => x"a4",
          2755 => x"0c",
          2756 => x"08",
          2757 => x"80",
          2758 => x"38",
          2759 => x"08",
          2760 => x"80",
          2761 => x"38",
          2762 => x"90",
          2763 => x"a4",
          2764 => x"34",
          2765 => x"08",
          2766 => x"70",
          2767 => x"71",
          2768 => x"51",
          2769 => x"82",
          2770 => x"f8",
          2771 => x"a4",
          2772 => x"82",
          2773 => x"f4",
          2774 => x"e0",
          2775 => x"05",
          2776 => x"81",
          2777 => x"70",
          2778 => x"72",
          2779 => x"a4",
          2780 => x"34",
          2781 => x"82",
          2782 => x"f8",
          2783 => x"72",
          2784 => x"38",
          2785 => x"e0",
          2786 => x"05",
          2787 => x"39",
          2788 => x"08",
          2789 => x"53",
          2790 => x"90",
          2791 => x"a4",
          2792 => x"33",
          2793 => x"26",
          2794 => x"39",
          2795 => x"e0",
          2796 => x"05",
          2797 => x"39",
          2798 => x"e0",
          2799 => x"05",
          2800 => x"82",
          2801 => x"f8",
          2802 => x"af",
          2803 => x"38",
          2804 => x"08",
          2805 => x"53",
          2806 => x"83",
          2807 => x"80",
          2808 => x"a4",
          2809 => x"0c",
          2810 => x"8a",
          2811 => x"a4",
          2812 => x"34",
          2813 => x"e0",
          2814 => x"05",
          2815 => x"a4",
          2816 => x"33",
          2817 => x"27",
          2818 => x"82",
          2819 => x"f8",
          2820 => x"80",
          2821 => x"94",
          2822 => x"a4",
          2823 => x"33",
          2824 => x"53",
          2825 => x"a4",
          2826 => x"34",
          2827 => x"08",
          2828 => x"d0",
          2829 => x"72",
          2830 => x"08",
          2831 => x"82",
          2832 => x"f8",
          2833 => x"90",
          2834 => x"38",
          2835 => x"08",
          2836 => x"f9",
          2837 => x"72",
          2838 => x"08",
          2839 => x"82",
          2840 => x"f8",
          2841 => x"72",
          2842 => x"38",
          2843 => x"e0",
          2844 => x"05",
          2845 => x"39",
          2846 => x"08",
          2847 => x"82",
          2848 => x"f4",
          2849 => x"54",
          2850 => x"8d",
          2851 => x"82",
          2852 => x"ec",
          2853 => x"f7",
          2854 => x"a4",
          2855 => x"33",
          2856 => x"a4",
          2857 => x"08",
          2858 => x"a4",
          2859 => x"33",
          2860 => x"e0",
          2861 => x"05",
          2862 => x"a4",
          2863 => x"08",
          2864 => x"05",
          2865 => x"08",
          2866 => x"55",
          2867 => x"82",
          2868 => x"f8",
          2869 => x"a5",
          2870 => x"a4",
          2871 => x"33",
          2872 => x"2e",
          2873 => x"e0",
          2874 => x"05",
          2875 => x"e0",
          2876 => x"05",
          2877 => x"a4",
          2878 => x"08",
          2879 => x"08",
          2880 => x"71",
          2881 => x"0b",
          2882 => x"08",
          2883 => x"82",
          2884 => x"ec",
          2885 => x"e0",
          2886 => x"3d",
          2887 => x"a4",
          2888 => x"e0",
          2889 => x"82",
          2890 => x"f7",
          2891 => x"0b",
          2892 => x"08",
          2893 => x"82",
          2894 => x"8c",
          2895 => x"80",
          2896 => x"e0",
          2897 => x"05",
          2898 => x"51",
          2899 => x"53",
          2900 => x"a4",
          2901 => x"34",
          2902 => x"06",
          2903 => x"2e",
          2904 => x"91",
          2905 => x"a4",
          2906 => x"08",
          2907 => x"05",
          2908 => x"ce",
          2909 => x"a4",
          2910 => x"33",
          2911 => x"2e",
          2912 => x"a4",
          2913 => x"82",
          2914 => x"f0",
          2915 => x"e0",
          2916 => x"05",
          2917 => x"81",
          2918 => x"70",
          2919 => x"72",
          2920 => x"a4",
          2921 => x"34",
          2922 => x"08",
          2923 => x"53",
          2924 => x"09",
          2925 => x"dc",
          2926 => x"a4",
          2927 => x"08",
          2928 => x"05",
          2929 => x"08",
          2930 => x"33",
          2931 => x"08",
          2932 => x"82",
          2933 => x"f8",
          2934 => x"e0",
          2935 => x"05",
          2936 => x"a4",
          2937 => x"08",
          2938 => x"b6",
          2939 => x"a4",
          2940 => x"08",
          2941 => x"84",
          2942 => x"39",
          2943 => x"e0",
          2944 => x"05",
          2945 => x"a4",
          2946 => x"08",
          2947 => x"05",
          2948 => x"08",
          2949 => x"33",
          2950 => x"08",
          2951 => x"81",
          2952 => x"0b",
          2953 => x"08",
          2954 => x"82",
          2955 => x"88",
          2956 => x"08",
          2957 => x"0c",
          2958 => x"53",
          2959 => x"e0",
          2960 => x"05",
          2961 => x"39",
          2962 => x"08",
          2963 => x"53",
          2964 => x"8d",
          2965 => x"82",
          2966 => x"ec",
          2967 => x"80",
          2968 => x"a4",
          2969 => x"33",
          2970 => x"27",
          2971 => x"e0",
          2972 => x"05",
          2973 => x"b9",
          2974 => x"8d",
          2975 => x"82",
          2976 => x"ec",
          2977 => x"d8",
          2978 => x"82",
          2979 => x"f4",
          2980 => x"39",
          2981 => x"08",
          2982 => x"53",
          2983 => x"90",
          2984 => x"a4",
          2985 => x"33",
          2986 => x"26",
          2987 => x"39",
          2988 => x"e0",
          2989 => x"05",
          2990 => x"39",
          2991 => x"e0",
          2992 => x"05",
          2993 => x"82",
          2994 => x"fc",
          2995 => x"e0",
          2996 => x"05",
          2997 => x"73",
          2998 => x"38",
          2999 => x"08",
          3000 => x"53",
          3001 => x"27",
          3002 => x"e0",
          3003 => x"05",
          3004 => x"51",
          3005 => x"e0",
          3006 => x"05",
          3007 => x"a4",
          3008 => x"33",
          3009 => x"53",
          3010 => x"a4",
          3011 => x"34",
          3012 => x"08",
          3013 => x"53",
          3014 => x"ad",
          3015 => x"a4",
          3016 => x"33",
          3017 => x"53",
          3018 => x"a4",
          3019 => x"34",
          3020 => x"08",
          3021 => x"53",
          3022 => x"8d",
          3023 => x"82",
          3024 => x"ec",
          3025 => x"98",
          3026 => x"a4",
          3027 => x"33",
          3028 => x"08",
          3029 => x"54",
          3030 => x"26",
          3031 => x"0b",
          3032 => x"08",
          3033 => x"80",
          3034 => x"e0",
          3035 => x"05",
          3036 => x"e0",
          3037 => x"05",
          3038 => x"e0",
          3039 => x"05",
          3040 => x"82",
          3041 => x"fc",
          3042 => x"e0",
          3043 => x"05",
          3044 => x"81",
          3045 => x"70",
          3046 => x"52",
          3047 => x"33",
          3048 => x"08",
          3049 => x"fe",
          3050 => x"e0",
          3051 => x"05",
          3052 => x"80",
          3053 => x"82",
          3054 => x"fc",
          3055 => x"82",
          3056 => x"fc",
          3057 => x"e0",
          3058 => x"05",
          3059 => x"a4",
          3060 => x"08",
          3061 => x"81",
          3062 => x"a4",
          3063 => x"0c",
          3064 => x"08",
          3065 => x"82",
          3066 => x"8b",
          3067 => x"e0",
          3068 => x"f8",
          3069 => x"70",
          3070 => x"56",
          3071 => x"2e",
          3072 => x"8c",
          3073 => x"79",
          3074 => x"33",
          3075 => x"39",
          3076 => x"73",
          3077 => x"81",
          3078 => x"81",
          3079 => x"39",
          3080 => x"90",
          3081 => x"a0",
          3082 => x"52",
          3083 => x"3f",
          3084 => x"08",
          3085 => x"08",
          3086 => x"76",
          3087 => x"df",
          3088 => x"e0",
          3089 => x"38",
          3090 => x"54",
          3091 => x"ff",
          3092 => x"17",
          3093 => x"06",
          3094 => x"77",
          3095 => x"ff",
          3096 => x"e0",
          3097 => x"3d",
          3098 => x"a0",
          3099 => x"98",
          3100 => x"3d",
          3101 => x"71",
          3102 => x"8e",
          3103 => x"29",
          3104 => x"05",
          3105 => x"04",
          3106 => x"51",
          3107 => x"82",
          3108 => x"80",
          3109 => x"be",
          3110 => x"f2",
          3111 => x"90",
          3112 => x"39",
          3113 => x"51",
          3114 => x"82",
          3115 => x"80",
          3116 => x"be",
          3117 => x"d6",
          3118 => x"d4",
          3119 => x"39",
          3120 => x"51",
          3121 => x"82",
          3122 => x"80",
          3123 => x"bf",
          3124 => x"39",
          3125 => x"51",
          3126 => x"bf",
          3127 => x"39",
          3128 => x"51",
          3129 => x"c0",
          3130 => x"39",
          3131 => x"51",
          3132 => x"c0",
          3133 => x"39",
          3134 => x"51",
          3135 => x"c0",
          3136 => x"39",
          3137 => x"51",
          3138 => x"c1",
          3139 => x"8a",
          3140 => x"0d",
          3141 => x"0d",
          3142 => x"56",
          3143 => x"26",
          3144 => x"52",
          3145 => x"29",
          3146 => x"87",
          3147 => x"51",
          3148 => x"82",
          3149 => x"52",
          3150 => x"9a",
          3151 => x"98",
          3152 => x"53",
          3153 => x"c1",
          3154 => x"b1",
          3155 => x"3d",
          3156 => x"3d",
          3157 => x"84",
          3158 => x"05",
          3159 => x"80",
          3160 => x"70",
          3161 => x"25",
          3162 => x"59",
          3163 => x"87",
          3164 => x"38",
          3165 => x"76",
          3166 => x"ff",
          3167 => x"93",
          3168 => x"82",
          3169 => x"76",
          3170 => x"70",
          3171 => x"93",
          3172 => x"e0",
          3173 => x"82",
          3174 => x"b9",
          3175 => x"98",
          3176 => x"98",
          3177 => x"e0",
          3178 => x"96",
          3179 => x"54",
          3180 => x"77",
          3181 => x"81",
          3182 => x"82",
          3183 => x"57",
          3184 => x"08",
          3185 => x"55",
          3186 => x"89",
          3187 => x"75",
          3188 => x"d7",
          3189 => x"d8",
          3190 => x"9f",
          3191 => x"30",
          3192 => x"80",
          3193 => x"70",
          3194 => x"06",
          3195 => x"56",
          3196 => x"90",
          3197 => x"bc",
          3198 => x"98",
          3199 => x"78",
          3200 => x"3f",
          3201 => x"82",
          3202 => x"96",
          3203 => x"f8",
          3204 => x"02",
          3205 => x"05",
          3206 => x"ff",
          3207 => x"7b",
          3208 => x"fe",
          3209 => x"e0",
          3210 => x"38",
          3211 => x"88",
          3212 => x"2e",
          3213 => x"39",
          3214 => x"56",
          3215 => x"54",
          3216 => x"53",
          3217 => x"51",
          3218 => x"e0",
          3219 => x"83",
          3220 => x"77",
          3221 => x"0c",
          3222 => x"04",
          3223 => x"7f",
          3224 => x"8c",
          3225 => x"05",
          3226 => x"15",
          3227 => x"5d",
          3228 => x"5e",
          3229 => x"fb",
          3230 => x"e0",
          3231 => x"ff",
          3232 => x"58",
          3233 => x"92",
          3234 => x"72",
          3235 => x"8a",
          3236 => x"80",
          3237 => x"39",
          3238 => x"52",
          3239 => x"51",
          3240 => x"3f",
          3241 => x"51",
          3242 => x"3f",
          3243 => x"78",
          3244 => x"38",
          3245 => x"89",
          3246 => x"2e",
          3247 => x"c6",
          3248 => x"53",
          3249 => x"8e",
          3250 => x"52",
          3251 => x"51",
          3252 => x"3f",
          3253 => x"c1",
          3254 => x"ae",
          3255 => x"15",
          3256 => x"39",
          3257 => x"72",
          3258 => x"38",
          3259 => x"82",
          3260 => x"ff",
          3261 => x"89",
          3262 => x"d8",
          3263 => x"8f",
          3264 => x"55",
          3265 => x"19",
          3266 => x"27",
          3267 => x"33",
          3268 => x"e4",
          3269 => x"f7",
          3270 => x"82",
          3271 => x"ff",
          3272 => x"81",
          3273 => x"fb",
          3274 => x"a0",
          3275 => x"3f",
          3276 => x"82",
          3277 => x"ff",
          3278 => x"80",
          3279 => x"27",
          3280 => x"74",
          3281 => x"55",
          3282 => x"72",
          3283 => x"38",
          3284 => x"53",
          3285 => x"83",
          3286 => x"75",
          3287 => x"81",
          3288 => x"53",
          3289 => x"90",
          3290 => x"fe",
          3291 => x"82",
          3292 => x"52",
          3293 => x"39",
          3294 => x"08",
          3295 => x"cc",
          3296 => x"15",
          3297 => x"39",
          3298 => x"51",
          3299 => x"77",
          3300 => x"5c",
          3301 => x"98",
          3302 => x"e0",
          3303 => x"2b",
          3304 => x"51",
          3305 => x"2e",
          3306 => x"ac",
          3307 => x"98",
          3308 => x"e0",
          3309 => x"2b",
          3310 => x"70",
          3311 => x"30",
          3312 => x"70",
          3313 => x"07",
          3314 => x"06",
          3315 => x"59",
          3316 => x"80",
          3317 => x"38",
          3318 => x"fd",
          3319 => x"1e",
          3320 => x"26",
          3321 => x"ff",
          3322 => x"e0",
          3323 => x"3d",
          3324 => x"3d",
          3325 => x"05",
          3326 => x"51",
          3327 => x"82",
          3328 => x"82",
          3329 => x"ff",
          3330 => x"82",
          3331 => x"51",
          3332 => x"82",
          3333 => x"82",
          3334 => x"82",
          3335 => x"52",
          3336 => x"51",
          3337 => x"3f",
          3338 => x"84",
          3339 => x"3f",
          3340 => x"04",
          3341 => x"87",
          3342 => x"08",
          3343 => x"3f",
          3344 => x"bf",
          3345 => x"b4",
          3346 => x"3f",
          3347 => x"b3",
          3348 => x"2a",
          3349 => x"51",
          3350 => x"2e",
          3351 => x"51",
          3352 => x"82",
          3353 => x"9a",
          3354 => x"51",
          3355 => x"72",
          3356 => x"81",
          3357 => x"71",
          3358 => x"38",
          3359 => x"83",
          3360 => x"dc",
          3361 => x"3f",
          3362 => x"f7",
          3363 => x"2a",
          3364 => x"51",
          3365 => x"2e",
          3366 => x"51",
          3367 => x"82",
          3368 => x"99",
          3369 => x"51",
          3370 => x"72",
          3371 => x"81",
          3372 => x"71",
          3373 => x"38",
          3374 => x"c7",
          3375 => x"80",
          3376 => x"3f",
          3377 => x"bb",
          3378 => x"2a",
          3379 => x"51",
          3380 => x"2e",
          3381 => x"51",
          3382 => x"82",
          3383 => x"99",
          3384 => x"51",
          3385 => x"72",
          3386 => x"81",
          3387 => x"71",
          3388 => x"38",
          3389 => x"8b",
          3390 => x"a8",
          3391 => x"3f",
          3392 => x"ff",
          3393 => x"2a",
          3394 => x"51",
          3395 => x"2e",
          3396 => x"51",
          3397 => x"82",
          3398 => x"99",
          3399 => x"51",
          3400 => x"72",
          3401 => x"81",
          3402 => x"71",
          3403 => x"38",
          3404 => x"cf",
          3405 => x"d0",
          3406 => x"3f",
          3407 => x"c3",
          3408 => x"3f",
          3409 => x"04",
          3410 => x"77",
          3411 => x"a3",
          3412 => x"55",
          3413 => x"52",
          3414 => x"ec",
          3415 => x"82",
          3416 => x"54",
          3417 => x"81",
          3418 => x"8c",
          3419 => x"a8",
          3420 => x"b6",
          3421 => x"98",
          3422 => x"82",
          3423 => x"07",
          3424 => x"71",
          3425 => x"54",
          3426 => x"82",
          3427 => x"0b",
          3428 => x"9c",
          3429 => x"81",
          3430 => x"06",
          3431 => x"f7",
          3432 => x"52",
          3433 => x"c7",
          3434 => x"e0",
          3435 => x"2e",
          3436 => x"e0",
          3437 => x"c4",
          3438 => x"39",
          3439 => x"51",
          3440 => x"3f",
          3441 => x"0b",
          3442 => x"34",
          3443 => x"db",
          3444 => x"73",
          3445 => x"81",
          3446 => x"82",
          3447 => x"74",
          3448 => x"aa",
          3449 => x"0b",
          3450 => x"0c",
          3451 => x"04",
          3452 => x"80",
          3453 => x"ff",
          3454 => x"a4",
          3455 => x"52",
          3456 => x"c8",
          3457 => x"e0",
          3458 => x"ff",
          3459 => x"7e",
          3460 => x"06",
          3461 => x"3d",
          3462 => x"82",
          3463 => x"78",
          3464 => x"3f",
          3465 => x"52",
          3466 => x"51",
          3467 => x"3f",
          3468 => x"08",
          3469 => x"38",
          3470 => x"51",
          3471 => x"81",
          3472 => x"82",
          3473 => x"ff",
          3474 => x"97",
          3475 => x"5a",
          3476 => x"79",
          3477 => x"3f",
          3478 => x"84",
          3479 => x"93",
          3480 => x"98",
          3481 => x"70",
          3482 => x"59",
          3483 => x"2e",
          3484 => x"78",
          3485 => x"b2",
          3486 => x"2e",
          3487 => x"78",
          3488 => x"38",
          3489 => x"ff",
          3490 => x"bc",
          3491 => x"38",
          3492 => x"78",
          3493 => x"83",
          3494 => x"80",
          3495 => x"ce",
          3496 => x"2e",
          3497 => x"8a",
          3498 => x"80",
          3499 => x"df",
          3500 => x"f9",
          3501 => x"78",
          3502 => x"88",
          3503 => x"80",
          3504 => x"a7",
          3505 => x"39",
          3506 => x"2e",
          3507 => x"78",
          3508 => x"8b",
          3509 => x"82",
          3510 => x"38",
          3511 => x"78",
          3512 => x"8a",
          3513 => x"86",
          3514 => x"ff",
          3515 => x"ff",
          3516 => x"ec",
          3517 => x"e0",
          3518 => x"2e",
          3519 => x"b5",
          3520 => x"11",
          3521 => x"05",
          3522 => x"3f",
          3523 => x"08",
          3524 => x"af",
          3525 => x"fe",
          3526 => x"ff",
          3527 => x"ec",
          3528 => x"e0",
          3529 => x"38",
          3530 => x"08",
          3531 => x"e8",
          3532 => x"db",
          3533 => x"5c",
          3534 => x"27",
          3535 => x"62",
          3536 => x"70",
          3537 => x"0c",
          3538 => x"f5",
          3539 => x"39",
          3540 => x"80",
          3541 => x"84",
          3542 => x"c6",
          3543 => x"98",
          3544 => x"fd",
          3545 => x"3d",
          3546 => x"53",
          3547 => x"51",
          3548 => x"82",
          3549 => x"80",
          3550 => x"38",
          3551 => x"f8",
          3552 => x"84",
          3553 => x"9a",
          3554 => x"98",
          3555 => x"fd",
          3556 => x"c4",
          3557 => x"a4",
          3558 => x"5a",
          3559 => x"81",
          3560 => x"59",
          3561 => x"05",
          3562 => x"34",
          3563 => x"43",
          3564 => x"3d",
          3565 => x"53",
          3566 => x"51",
          3567 => x"82",
          3568 => x"80",
          3569 => x"38",
          3570 => x"fc",
          3571 => x"84",
          3572 => x"ce",
          3573 => x"98",
          3574 => x"fc",
          3575 => x"3d",
          3576 => x"53",
          3577 => x"51",
          3578 => x"82",
          3579 => x"80",
          3580 => x"38",
          3581 => x"51",
          3582 => x"3f",
          3583 => x"64",
          3584 => x"62",
          3585 => x"33",
          3586 => x"78",
          3587 => x"38",
          3588 => x"54",
          3589 => x"79",
          3590 => x"94",
          3591 => x"ef",
          3592 => x"63",
          3593 => x"5a",
          3594 => x"51",
          3595 => x"fc",
          3596 => x"3d",
          3597 => x"53",
          3598 => x"51",
          3599 => x"82",
          3600 => x"80",
          3601 => x"de",
          3602 => x"78",
          3603 => x"38",
          3604 => x"08",
          3605 => x"39",
          3606 => x"33",
          3607 => x"2e",
          3608 => x"de",
          3609 => x"bc",
          3610 => x"fe",
          3611 => x"80",
          3612 => x"82",
          3613 => x"45",
          3614 => x"de",
          3615 => x"78",
          3616 => x"38",
          3617 => x"08",
          3618 => x"82",
          3619 => x"59",
          3620 => x"88",
          3621 => x"d4",
          3622 => x"39",
          3623 => x"08",
          3624 => x"45",
          3625 => x"fc",
          3626 => x"84",
          3627 => x"f2",
          3628 => x"98",
          3629 => x"38",
          3630 => x"33",
          3631 => x"2e",
          3632 => x"de",
          3633 => x"80",
          3634 => x"de",
          3635 => x"78",
          3636 => x"38",
          3637 => x"08",
          3638 => x"82",
          3639 => x"59",
          3640 => x"88",
          3641 => x"c8",
          3642 => x"39",
          3643 => x"33",
          3644 => x"2e",
          3645 => x"de",
          3646 => x"99",
          3647 => x"fa",
          3648 => x"80",
          3649 => x"82",
          3650 => x"44",
          3651 => x"de",
          3652 => x"05",
          3653 => x"fe",
          3654 => x"ff",
          3655 => x"e8",
          3656 => x"e0",
          3657 => x"2e",
          3658 => x"63",
          3659 => x"88",
          3660 => x"81",
          3661 => x"32",
          3662 => x"72",
          3663 => x"70",
          3664 => x"51",
          3665 => x"80",
          3666 => x"7a",
          3667 => x"38",
          3668 => x"c5",
          3669 => x"bd",
          3670 => x"55",
          3671 => x"53",
          3672 => x"51",
          3673 => x"82",
          3674 => x"87",
          3675 => x"3d",
          3676 => x"53",
          3677 => x"51",
          3678 => x"82",
          3679 => x"80",
          3680 => x"38",
          3681 => x"fc",
          3682 => x"84",
          3683 => x"92",
          3684 => x"98",
          3685 => x"a4",
          3686 => x"02",
          3687 => x"33",
          3688 => x"81",
          3689 => x"3d",
          3690 => x"53",
          3691 => x"51",
          3692 => x"82",
          3693 => x"e1",
          3694 => x"39",
          3695 => x"54",
          3696 => x"c8",
          3697 => x"c7",
          3698 => x"f8",
          3699 => x"f8",
          3700 => x"ff",
          3701 => x"79",
          3702 => x"59",
          3703 => x"f8",
          3704 => x"79",
          3705 => x"b5",
          3706 => x"11",
          3707 => x"05",
          3708 => x"3f",
          3709 => x"08",
          3710 => x"38",
          3711 => x"80",
          3712 => x"79",
          3713 => x"05",
          3714 => x"39",
          3715 => x"51",
          3716 => x"3f",
          3717 => x"b5",
          3718 => x"11",
          3719 => x"05",
          3720 => x"3f",
          3721 => x"08",
          3722 => x"97",
          3723 => x"fe",
          3724 => x"ff",
          3725 => x"e0",
          3726 => x"e0",
          3727 => x"2e",
          3728 => x"59",
          3729 => x"05",
          3730 => x"82",
          3731 => x"78",
          3732 => x"fe",
          3733 => x"ff",
          3734 => x"df",
          3735 => x"e0",
          3736 => x"38",
          3737 => x"61",
          3738 => x"52",
          3739 => x"51",
          3740 => x"3f",
          3741 => x"08",
          3742 => x"52",
          3743 => x"9f",
          3744 => x"46",
          3745 => x"78",
          3746 => x"b7",
          3747 => x"26",
          3748 => x"82",
          3749 => x"39",
          3750 => x"f0",
          3751 => x"84",
          3752 => x"ad",
          3753 => x"98",
          3754 => x"93",
          3755 => x"02",
          3756 => x"22",
          3757 => x"05",
          3758 => x"42",
          3759 => x"82",
          3760 => x"ff",
          3761 => x"ff",
          3762 => x"3d",
          3763 => x"53",
          3764 => x"51",
          3765 => x"82",
          3766 => x"80",
          3767 => x"38",
          3768 => x"f0",
          3769 => x"84",
          3770 => x"e5",
          3771 => x"98",
          3772 => x"a0",
          3773 => x"71",
          3774 => x"84",
          3775 => x"3d",
          3776 => x"53",
          3777 => x"51",
          3778 => x"82",
          3779 => x"e5",
          3780 => x"39",
          3781 => x"54",
          3782 => x"e4",
          3783 => x"ef",
          3784 => x"f8",
          3785 => x"f8",
          3786 => x"ff",
          3787 => x"79",
          3788 => x"59",
          3789 => x"f6",
          3790 => x"79",
          3791 => x"b5",
          3792 => x"11",
          3793 => x"05",
          3794 => x"3f",
          3795 => x"08",
          3796 => x"38",
          3797 => x"0c",
          3798 => x"05",
          3799 => x"39",
          3800 => x"51",
          3801 => x"3f",
          3802 => x"b5",
          3803 => x"11",
          3804 => x"05",
          3805 => x"3f",
          3806 => x"08",
          3807 => x"c3",
          3808 => x"82",
          3809 => x"ff",
          3810 => x"64",
          3811 => x"b5",
          3812 => x"11",
          3813 => x"05",
          3814 => x"3f",
          3815 => x"08",
          3816 => x"9f",
          3817 => x"82",
          3818 => x"ff",
          3819 => x"64",
          3820 => x"82",
          3821 => x"80",
          3822 => x"38",
          3823 => x"08",
          3824 => x"ac",
          3825 => x"c7",
          3826 => x"39",
          3827 => x"51",
          3828 => x"3f",
          3829 => x"3f",
          3830 => x"82",
          3831 => x"ff",
          3832 => x"80",
          3833 => x"39",
          3834 => x"f4",
          3835 => x"3d",
          3836 => x"80",
          3837 => x"38",
          3838 => x"79",
          3839 => x"3f",
          3840 => x"08",
          3841 => x"98",
          3842 => x"82",
          3843 => x"e0",
          3844 => x"b5",
          3845 => x"05",
          3846 => x"3f",
          3847 => x"08",
          3848 => x"5a",
          3849 => x"2e",
          3850 => x"82",
          3851 => x"51",
          3852 => x"82",
          3853 => x"8f",
          3854 => x"38",
          3855 => x"82",
          3856 => x"7a",
          3857 => x"38",
          3858 => x"8c",
          3859 => x"39",
          3860 => x"ad",
          3861 => x"39",
          3862 => x"56",
          3863 => x"c6",
          3864 => x"53",
          3865 => x"52",
          3866 => x"b0",
          3867 => x"9e",
          3868 => x"39",
          3869 => x"3d",
          3870 => x"51",
          3871 => x"ab",
          3872 => x"82",
          3873 => x"80",
          3874 => x"90",
          3875 => x"ff",
          3876 => x"ff",
          3877 => x"93",
          3878 => x"80",
          3879 => x"9c",
          3880 => x"ff",
          3881 => x"ff",
          3882 => x"82",
          3883 => x"82",
          3884 => x"7c",
          3885 => x"80",
          3886 => x"0a",
          3887 => x"0a",
          3888 => x"ff",
          3889 => x"ea",
          3890 => x"e0",
          3891 => x"e0",
          3892 => x"70",
          3893 => x"07",
          3894 => x"5b",
          3895 => x"5a",
          3896 => x"83",
          3897 => x"78",
          3898 => x"78",
          3899 => x"38",
          3900 => x"81",
          3901 => x"59",
          3902 => x"38",
          3903 => x"7e",
          3904 => x"59",
          3905 => x"7e",
          3906 => x"81",
          3907 => x"82",
          3908 => x"ff",
          3909 => x"7c",
          3910 => x"3f",
          3911 => x"82",
          3912 => x"ff",
          3913 => x"f2",
          3914 => x"3d",
          3915 => x"82",
          3916 => x"87",
          3917 => x"70",
          3918 => x"87",
          3919 => x"72",
          3920 => x"3f",
          3921 => x"08",
          3922 => x"08",
          3923 => x"84",
          3924 => x"51",
          3925 => x"72",
          3926 => x"08",
          3927 => x"87",
          3928 => x"70",
          3929 => x"87",
          3930 => x"72",
          3931 => x"3f",
          3932 => x"08",
          3933 => x"08",
          3934 => x"84",
          3935 => x"51",
          3936 => x"72",
          3937 => x"08",
          3938 => x"8c",
          3939 => x"87",
          3940 => x"0c",
          3941 => x"0b",
          3942 => x"94",
          3943 => x"98",
          3944 => x"84",
          3945 => x"84",
          3946 => x"34",
          3947 => x"fb",
          3948 => x"3d",
          3949 => x"0c",
          3950 => x"82",
          3951 => x"54",
          3952 => x"93",
          3953 => x"c7",
          3954 => x"b4",
          3955 => x"c7",
          3956 => x"b4",
          3957 => x"e8",
          3958 => x"d2",
          3959 => x"ec",
          3960 => x"8c",
          3961 => x"fc",
          3962 => x"70",
          3963 => x"80",
          3964 => x"72",
          3965 => x"8a",
          3966 => x"51",
          3967 => x"09",
          3968 => x"38",
          3969 => x"f1",
          3970 => x"51",
          3971 => x"09",
          3972 => x"38",
          3973 => x"81",
          3974 => x"73",
          3975 => x"81",
          3976 => x"84",
          3977 => x"52",
          3978 => x"52",
          3979 => x"2e",
          3980 => x"54",
          3981 => x"9d",
          3982 => x"38",
          3983 => x"12",
          3984 => x"33",
          3985 => x"a0",
          3986 => x"81",
          3987 => x"2e",
          3988 => x"ea",
          3989 => x"33",
          3990 => x"a0",
          3991 => x"06",
          3992 => x"54",
          3993 => x"70",
          3994 => x"25",
          3995 => x"51",
          3996 => x"2e",
          3997 => x"72",
          3998 => x"54",
          3999 => x"0c",
          4000 => x"82",
          4001 => x"86",
          4002 => x"fc",
          4003 => x"53",
          4004 => x"2e",
          4005 => x"3d",
          4006 => x"72",
          4007 => x"3f",
          4008 => x"08",
          4009 => x"53",
          4010 => x"53",
          4011 => x"98",
          4012 => x"0d",
          4013 => x"0d",
          4014 => x"33",
          4015 => x"53",
          4016 => x"8b",
          4017 => x"38",
          4018 => x"ff",
          4019 => x"52",
          4020 => x"81",
          4021 => x"13",
          4022 => x"52",
          4023 => x"80",
          4024 => x"13",
          4025 => x"52",
          4026 => x"80",
          4027 => x"13",
          4028 => x"52",
          4029 => x"80",
          4030 => x"13",
          4031 => x"52",
          4032 => x"26",
          4033 => x"8a",
          4034 => x"87",
          4035 => x"e7",
          4036 => x"38",
          4037 => x"c0",
          4038 => x"72",
          4039 => x"98",
          4040 => x"13",
          4041 => x"98",
          4042 => x"13",
          4043 => x"98",
          4044 => x"13",
          4045 => x"98",
          4046 => x"13",
          4047 => x"98",
          4048 => x"13",
          4049 => x"98",
          4050 => x"87",
          4051 => x"0c",
          4052 => x"98",
          4053 => x"0b",
          4054 => x"9c",
          4055 => x"71",
          4056 => x"0c",
          4057 => x"04",
          4058 => x"7f",
          4059 => x"98",
          4060 => x"7d",
          4061 => x"98",
          4062 => x"7d",
          4063 => x"c0",
          4064 => x"5a",
          4065 => x"34",
          4066 => x"b4",
          4067 => x"83",
          4068 => x"c0",
          4069 => x"5a",
          4070 => x"34",
          4071 => x"ac",
          4072 => x"85",
          4073 => x"c0",
          4074 => x"5a",
          4075 => x"34",
          4076 => x"a4",
          4077 => x"88",
          4078 => x"c0",
          4079 => x"5a",
          4080 => x"23",
          4081 => x"79",
          4082 => x"06",
          4083 => x"ff",
          4084 => x"86",
          4085 => x"85",
          4086 => x"84",
          4087 => x"83",
          4088 => x"82",
          4089 => x"7d",
          4090 => x"06",
          4091 => x"84",
          4092 => x"9b",
          4093 => x"0d",
          4094 => x"0d",
          4095 => x"33",
          4096 => x"72",
          4097 => x"81",
          4098 => x"72",
          4099 => x"32",
          4100 => x"80",
          4101 => x"51",
          4102 => x"80",
          4103 => x"84",
          4104 => x"39",
          4105 => x"82",
          4106 => x"98",
          4107 => x"2c",
          4108 => x"ff",
          4109 => x"06",
          4110 => x"54",
          4111 => x"09",
          4112 => x"38",
          4113 => x"83",
          4114 => x"70",
          4115 => x"07",
          4116 => x"70",
          4117 => x"71",
          4118 => x"0c",
          4119 => x"04",
          4120 => x"80",
          4121 => x"72",
          4122 => x"81",
          4123 => x"3f",
          4124 => x"08",
          4125 => x"98",
          4126 => x"ff",
          4127 => x"52",
          4128 => x"e3",
          4129 => x"e0",
          4130 => x"3d",
          4131 => x"3d",
          4132 => x"05",
          4133 => x"b0",
          4134 => x"ff",
          4135 => x"55",
          4136 => x"84",
          4137 => x"2e",
          4138 => x"c0",
          4139 => x"70",
          4140 => x"2a",
          4141 => x"53",
          4142 => x"80",
          4143 => x"71",
          4144 => x"81",
          4145 => x"70",
          4146 => x"81",
          4147 => x"06",
          4148 => x"80",
          4149 => x"71",
          4150 => x"81",
          4151 => x"70",
          4152 => x"73",
          4153 => x"51",
          4154 => x"80",
          4155 => x"2e",
          4156 => x"c0",
          4157 => x"74",
          4158 => x"82",
          4159 => x"87",
          4160 => x"ff",
          4161 => x"8f",
          4162 => x"30",
          4163 => x"51",
          4164 => x"82",
          4165 => x"83",
          4166 => x"f9",
          4167 => x"a7",
          4168 => x"77",
          4169 => x"81",
          4170 => x"7a",
          4171 => x"eb",
          4172 => x"b0",
          4173 => x"ff",
          4174 => x"87",
          4175 => x"53",
          4176 => x"86",
          4177 => x"94",
          4178 => x"08",
          4179 => x"70",
          4180 => x"56",
          4181 => x"2e",
          4182 => x"91",
          4183 => x"06",
          4184 => x"d7",
          4185 => x"32",
          4186 => x"51",
          4187 => x"2e",
          4188 => x"93",
          4189 => x"06",
          4190 => x"ff",
          4191 => x"81",
          4192 => x"87",
          4193 => x"54",
          4194 => x"86",
          4195 => x"94",
          4196 => x"74",
          4197 => x"82",
          4198 => x"89",
          4199 => x"f9",
          4200 => x"54",
          4201 => x"70",
          4202 => x"53",
          4203 => x"77",
          4204 => x"38",
          4205 => x"06",
          4206 => x"de",
          4207 => x"81",
          4208 => x"57",
          4209 => x"c0",
          4210 => x"75",
          4211 => x"38",
          4212 => x"94",
          4213 => x"70",
          4214 => x"81",
          4215 => x"52",
          4216 => x"8c",
          4217 => x"2a",
          4218 => x"51",
          4219 => x"38",
          4220 => x"70",
          4221 => x"51",
          4222 => x"8d",
          4223 => x"2a",
          4224 => x"51",
          4225 => x"be",
          4226 => x"ff",
          4227 => x"c0",
          4228 => x"70",
          4229 => x"38",
          4230 => x"90",
          4231 => x"0c",
          4232 => x"33",
          4233 => x"06",
          4234 => x"70",
          4235 => x"76",
          4236 => x"0c",
          4237 => x"04",
          4238 => x"82",
          4239 => x"70",
          4240 => x"54",
          4241 => x"94",
          4242 => x"80",
          4243 => x"87",
          4244 => x"51",
          4245 => x"82",
          4246 => x"06",
          4247 => x"70",
          4248 => x"38",
          4249 => x"06",
          4250 => x"94",
          4251 => x"80",
          4252 => x"87",
          4253 => x"52",
          4254 => x"81",
          4255 => x"e0",
          4256 => x"84",
          4257 => x"ff",
          4258 => x"e0",
          4259 => x"ff",
          4260 => x"98",
          4261 => x"3d",
          4262 => x"b0",
          4263 => x"ff",
          4264 => x"87",
          4265 => x"52",
          4266 => x"86",
          4267 => x"94",
          4268 => x"08",
          4269 => x"70",
          4270 => x"51",
          4271 => x"70",
          4272 => x"38",
          4273 => x"06",
          4274 => x"94",
          4275 => x"80",
          4276 => x"87",
          4277 => x"52",
          4278 => x"98",
          4279 => x"2c",
          4280 => x"71",
          4281 => x"0c",
          4282 => x"04",
          4283 => x"87",
          4284 => x"08",
          4285 => x"8a",
          4286 => x"70",
          4287 => x"b4",
          4288 => x"9e",
          4289 => x"de",
          4290 => x"c0",
          4291 => x"82",
          4292 => x"87",
          4293 => x"08",
          4294 => x"0c",
          4295 => x"98",
          4296 => x"c0",
          4297 => x"9e",
          4298 => x"de",
          4299 => x"c0",
          4300 => x"82",
          4301 => x"87",
          4302 => x"08",
          4303 => x"0c",
          4304 => x"b0",
          4305 => x"d0",
          4306 => x"9e",
          4307 => x"de",
          4308 => x"c0",
          4309 => x"82",
          4310 => x"87",
          4311 => x"08",
          4312 => x"0c",
          4313 => x"c0",
          4314 => x"e0",
          4315 => x"9e",
          4316 => x"de",
          4317 => x"c0",
          4318 => x"51",
          4319 => x"e8",
          4320 => x"9e",
          4321 => x"de",
          4322 => x"c0",
          4323 => x"82",
          4324 => x"87",
          4325 => x"08",
          4326 => x"0c",
          4327 => x"de",
          4328 => x"0b",
          4329 => x"90",
          4330 => x"80",
          4331 => x"52",
          4332 => x"2e",
          4333 => x"52",
          4334 => x"f9",
          4335 => x"87",
          4336 => x"08",
          4337 => x"0a",
          4338 => x"52",
          4339 => x"83",
          4340 => x"71",
          4341 => x"34",
          4342 => x"c0",
          4343 => x"70",
          4344 => x"06",
          4345 => x"70",
          4346 => x"38",
          4347 => x"82",
          4348 => x"80",
          4349 => x"9e",
          4350 => x"88",
          4351 => x"51",
          4352 => x"80",
          4353 => x"81",
          4354 => x"de",
          4355 => x"0b",
          4356 => x"90",
          4357 => x"80",
          4358 => x"52",
          4359 => x"2e",
          4360 => x"52",
          4361 => x"fd",
          4362 => x"87",
          4363 => x"08",
          4364 => x"80",
          4365 => x"52",
          4366 => x"83",
          4367 => x"71",
          4368 => x"34",
          4369 => x"c0",
          4370 => x"70",
          4371 => x"06",
          4372 => x"70",
          4373 => x"38",
          4374 => x"82",
          4375 => x"80",
          4376 => x"9e",
          4377 => x"82",
          4378 => x"51",
          4379 => x"80",
          4380 => x"81",
          4381 => x"df",
          4382 => x"0b",
          4383 => x"90",
          4384 => x"80",
          4385 => x"52",
          4386 => x"2e",
          4387 => x"52",
          4388 => x"81",
          4389 => x"87",
          4390 => x"08",
          4391 => x"80",
          4392 => x"52",
          4393 => x"83",
          4394 => x"71",
          4395 => x"34",
          4396 => x"c0",
          4397 => x"70",
          4398 => x"51",
          4399 => x"80",
          4400 => x"81",
          4401 => x"df",
          4402 => x"c0",
          4403 => x"70",
          4404 => x"70",
          4405 => x"51",
          4406 => x"df",
          4407 => x"0b",
          4408 => x"90",
          4409 => x"80",
          4410 => x"52",
          4411 => x"83",
          4412 => x"71",
          4413 => x"34",
          4414 => x"90",
          4415 => x"f0",
          4416 => x"2a",
          4417 => x"70",
          4418 => x"34",
          4419 => x"c0",
          4420 => x"70",
          4421 => x"52",
          4422 => x"2e",
          4423 => x"52",
          4424 => x"87",
          4425 => x"9e",
          4426 => x"87",
          4427 => x"70",
          4428 => x"34",
          4429 => x"04",
          4430 => x"82",
          4431 => x"ff",
          4432 => x"82",
          4433 => x"54",
          4434 => x"89",
          4435 => x"b0",
          4436 => x"bb",
          4437 => x"c4",
          4438 => x"be",
          4439 => x"fa",
          4440 => x"80",
          4441 => x"82",
          4442 => x"82",
          4443 => x"11",
          4444 => x"c8",
          4445 => x"89",
          4446 => x"de",
          4447 => x"73",
          4448 => x"38",
          4449 => x"08",
          4450 => x"08",
          4451 => x"82",
          4452 => x"ff",
          4453 => x"82",
          4454 => x"54",
          4455 => x"94",
          4456 => x"b4",
          4457 => x"b8",
          4458 => x"52",
          4459 => x"51",
          4460 => x"3f",
          4461 => x"33",
          4462 => x"2e",
          4463 => x"de",
          4464 => x"de",
          4465 => x"54",
          4466 => x"b0",
          4467 => x"bf",
          4468 => x"fe",
          4469 => x"80",
          4470 => x"82",
          4471 => x"82",
          4472 => x"11",
          4473 => x"c9",
          4474 => x"88",
          4475 => x"df",
          4476 => x"73",
          4477 => x"38",
          4478 => x"33",
          4479 => x"e8",
          4480 => x"8b",
          4481 => x"87",
          4482 => x"80",
          4483 => x"82",
          4484 => x"52",
          4485 => x"51",
          4486 => x"3f",
          4487 => x"33",
          4488 => x"2e",
          4489 => x"df",
          4490 => x"82",
          4491 => x"ff",
          4492 => x"82",
          4493 => x"54",
          4494 => x"89",
          4495 => x"c8",
          4496 => x"d6",
          4497 => x"fb",
          4498 => x"80",
          4499 => x"82",
          4500 => x"ff",
          4501 => x"82",
          4502 => x"54",
          4503 => x"89",
          4504 => x"e8",
          4505 => x"b2",
          4506 => x"81",
          4507 => x"80",
          4508 => x"82",
          4509 => x"ff",
          4510 => x"82",
          4511 => x"54",
          4512 => x"89",
          4513 => x"fc",
          4514 => x"8e",
          4515 => x"84",
          4516 => x"86",
          4517 => x"dc",
          4518 => x"cb",
          4519 => x"86",
          4520 => x"de",
          4521 => x"82",
          4522 => x"ff",
          4523 => x"82",
          4524 => x"52",
          4525 => x"51",
          4526 => x"3f",
          4527 => x"51",
          4528 => x"3f",
          4529 => x"22",
          4530 => x"90",
          4531 => x"bf",
          4532 => x"ec",
          4533 => x"84",
          4534 => x"51",
          4535 => x"3f",
          4536 => x"08",
          4537 => x"29",
          4538 => x"54",
          4539 => x"98",
          4540 => x"cc",
          4541 => x"86",
          4542 => x"de",
          4543 => x"73",
          4544 => x"38",
          4545 => x"08",
          4546 => x"c0",
          4547 => x"ff",
          4548 => x"82",
          4549 => x"bd",
          4550 => x"76",
          4551 => x"54",
          4552 => x"08",
          4553 => x"e4",
          4554 => x"e3",
          4555 => x"fa",
          4556 => x"80",
          4557 => x"82",
          4558 => x"56",
          4559 => x"52",
          4560 => x"b7",
          4561 => x"e0",
          4562 => x"84",
          4563 => x"71",
          4564 => x"82",
          4565 => x"52",
          4566 => x"51",
          4567 => x"3f",
          4568 => x"a4",
          4569 => x"3d",
          4570 => x"3d",
          4571 => x"05",
          4572 => x"52",
          4573 => x"aa",
          4574 => x"29",
          4575 => x"05",
          4576 => x"04",
          4577 => x"51",
          4578 => x"cd",
          4579 => x"39",
          4580 => x"51",
          4581 => x"cd",
          4582 => x"39",
          4583 => x"51",
          4584 => x"cd",
          4585 => x"84",
          4586 => x"3d",
          4587 => x"88",
          4588 => x"80",
          4589 => x"96",
          4590 => x"82",
          4591 => x"87",
          4592 => x"0c",
          4593 => x"0d",
          4594 => x"70",
          4595 => x"98",
          4596 => x"2c",
          4597 => x"70",
          4598 => x"53",
          4599 => x"51",
          4600 => x"cd",
          4601 => x"55",
          4602 => x"25",
          4603 => x"cd",
          4604 => x"12",
          4605 => x"97",
          4606 => x"33",
          4607 => x"70",
          4608 => x"81",
          4609 => x"81",
          4610 => x"e0",
          4611 => x"3d",
          4612 => x"3d",
          4613 => x"84",
          4614 => x"33",
          4615 => x"56",
          4616 => x"2e",
          4617 => x"fb",
          4618 => x"88",
          4619 => x"b9",
          4620 => x"fc",
          4621 => x"51",
          4622 => x"3f",
          4623 => x"08",
          4624 => x"ff",
          4625 => x"73",
          4626 => x"53",
          4627 => x"72",
          4628 => x"53",
          4629 => x"51",
          4630 => x"3f",
          4631 => x"87",
          4632 => x"f6",
          4633 => x"02",
          4634 => x"05",
          4635 => x"05",
          4636 => x"82",
          4637 => x"70",
          4638 => x"df",
          4639 => x"08",
          4640 => x"5a",
          4641 => x"80",
          4642 => x"74",
          4643 => x"3f",
          4644 => x"33",
          4645 => x"82",
          4646 => x"81",
          4647 => x"58",
          4648 => x"fe",
          4649 => x"98",
          4650 => x"82",
          4651 => x"70",
          4652 => x"df",
          4653 => x"08",
          4654 => x"74",
          4655 => x"38",
          4656 => x"52",
          4657 => x"ac",
          4658 => x"df",
          4659 => x"05",
          4660 => x"df",
          4661 => x"81",
          4662 => x"93",
          4663 => x"38",
          4664 => x"df",
          4665 => x"80",
          4666 => x"82",
          4667 => x"56",
          4668 => x"ac",
          4669 => x"e0",
          4670 => x"a4",
          4671 => x"fc",
          4672 => x"53",
          4673 => x"51",
          4674 => x"3f",
          4675 => x"08",
          4676 => x"81",
          4677 => x"82",
          4678 => x"51",
          4679 => x"3f",
          4680 => x"04",
          4681 => x"82",
          4682 => x"93",
          4683 => x"52",
          4684 => x"89",
          4685 => x"99",
          4686 => x"73",
          4687 => x"84",
          4688 => x"73",
          4689 => x"38",
          4690 => x"df",
          4691 => x"df",
          4692 => x"71",
          4693 => x"38",
          4694 => x"f0",
          4695 => x"df",
          4696 => x"99",
          4697 => x"0b",
          4698 => x"0c",
          4699 => x"04",
          4700 => x"81",
          4701 => x"82",
          4702 => x"51",
          4703 => x"3f",
          4704 => x"08",
          4705 => x"82",
          4706 => x"53",
          4707 => x"88",
          4708 => x"56",
          4709 => x"3f",
          4710 => x"08",
          4711 => x"38",
          4712 => x"a9",
          4713 => x"e0",
          4714 => x"80",
          4715 => x"98",
          4716 => x"38",
          4717 => x"08",
          4718 => x"17",
          4719 => x"74",
          4720 => x"76",
          4721 => x"82",
          4722 => x"57",
          4723 => x"3f",
          4724 => x"09",
          4725 => x"af",
          4726 => x"0d",
          4727 => x"0d",
          4728 => x"ad",
          4729 => x"5a",
          4730 => x"58",
          4731 => x"df",
          4732 => x"80",
          4733 => x"82",
          4734 => x"81",
          4735 => x"0b",
          4736 => x"08",
          4737 => x"f8",
          4738 => x"70",
          4739 => x"9e",
          4740 => x"e0",
          4741 => x"2e",
          4742 => x"51",
          4743 => x"3f",
          4744 => x"08",
          4745 => x"55",
          4746 => x"e0",
          4747 => x"8e",
          4748 => x"98",
          4749 => x"70",
          4750 => x"80",
          4751 => x"09",
          4752 => x"72",
          4753 => x"51",
          4754 => x"77",
          4755 => x"73",
          4756 => x"82",
          4757 => x"8c",
          4758 => x"51",
          4759 => x"3f",
          4760 => x"08",
          4761 => x"38",
          4762 => x"51",
          4763 => x"3f",
          4764 => x"09",
          4765 => x"38",
          4766 => x"51",
          4767 => x"3f",
          4768 => x"a7",
          4769 => x"3d",
          4770 => x"e0",
          4771 => x"34",
          4772 => x"82",
          4773 => x"a9",
          4774 => x"f6",
          4775 => x"7e",
          4776 => x"72",
          4777 => x"5a",
          4778 => x"2e",
          4779 => x"a2",
          4780 => x"78",
          4781 => x"76",
          4782 => x"81",
          4783 => x"70",
          4784 => x"58",
          4785 => x"2e",
          4786 => x"86",
          4787 => x"26",
          4788 => x"54",
          4789 => x"82",
          4790 => x"70",
          4791 => x"ff",
          4792 => x"82",
          4793 => x"53",
          4794 => x"08",
          4795 => x"d9",
          4796 => x"98",
          4797 => x"38",
          4798 => x"55",
          4799 => x"88",
          4800 => x"2e",
          4801 => x"39",
          4802 => x"ac",
          4803 => x"5a",
          4804 => x"11",
          4805 => x"51",
          4806 => x"82",
          4807 => x"80",
          4808 => x"ff",
          4809 => x"52",
          4810 => x"b1",
          4811 => x"98",
          4812 => x"06",
          4813 => x"38",
          4814 => x"39",
          4815 => x"81",
          4816 => x"54",
          4817 => x"ff",
          4818 => x"54",
          4819 => x"98",
          4820 => x"0d",
          4821 => x"0d",
          4822 => x"b2",
          4823 => x"3d",
          4824 => x"5a",
          4825 => x"3d",
          4826 => x"e8",
          4827 => x"e4",
          4828 => x"73",
          4829 => x"73",
          4830 => x"33",
          4831 => x"83",
          4832 => x"76",
          4833 => x"bc",
          4834 => x"76",
          4835 => x"73",
          4836 => x"ad",
          4837 => x"98",
          4838 => x"e0",
          4839 => x"df",
          4840 => x"e0",
          4841 => x"2e",
          4842 => x"93",
          4843 => x"82",
          4844 => x"51",
          4845 => x"3f",
          4846 => x"08",
          4847 => x"38",
          4848 => x"51",
          4849 => x"3f",
          4850 => x"82",
          4851 => x"5b",
          4852 => x"08",
          4853 => x"52",
          4854 => x"52",
          4855 => x"f8",
          4856 => x"98",
          4857 => x"e0",
          4858 => x"2e",
          4859 => x"80",
          4860 => x"e0",
          4861 => x"ff",
          4862 => x"82",
          4863 => x"55",
          4864 => x"e0",
          4865 => x"a9",
          4866 => x"98",
          4867 => x"70",
          4868 => x"80",
          4869 => x"53",
          4870 => x"06",
          4871 => x"f8",
          4872 => x"1b",
          4873 => x"06",
          4874 => x"7b",
          4875 => x"80",
          4876 => x"2e",
          4877 => x"ff",
          4878 => x"39",
          4879 => x"e0",
          4880 => x"38",
          4881 => x"08",
          4882 => x"38",
          4883 => x"8f",
          4884 => x"51",
          4885 => x"82",
          4886 => x"98",
          4887 => x"2c",
          4888 => x"ff",
          4889 => x"78",
          4890 => x"82",
          4891 => x"70",
          4892 => x"98",
          4893 => x"d0",
          4894 => x"2b",
          4895 => x"71",
          4896 => x"70",
          4897 => x"cd",
          4898 => x"08",
          4899 => x"51",
          4900 => x"59",
          4901 => x"5d",
          4902 => x"73",
          4903 => x"e9",
          4904 => x"27",
          4905 => x"81",
          4906 => x"81",
          4907 => x"70",
          4908 => x"55",
          4909 => x"80",
          4910 => x"53",
          4911 => x"51",
          4912 => x"82",
          4913 => x"81",
          4914 => x"73",
          4915 => x"38",
          4916 => x"d0",
          4917 => x"b1",
          4918 => x"80",
          4919 => x"80",
          4920 => x"98",
          4921 => x"ff",
          4922 => x"55",
          4923 => x"97",
          4924 => x"74",
          4925 => x"f5",
          4926 => x"e0",
          4927 => x"ff",
          4928 => x"cc",
          4929 => x"80",
          4930 => x"2e",
          4931 => x"81",
          4932 => x"82",
          4933 => x"74",
          4934 => x"98",
          4935 => x"d0",
          4936 => x"2b",
          4937 => x"70",
          4938 => x"82",
          4939 => x"ec",
          4940 => x"51",
          4941 => x"58",
          4942 => x"77",
          4943 => x"06",
          4944 => x"82",
          4945 => x"08",
          4946 => x"0b",
          4947 => x"34",
          4948 => x"f7",
          4949 => x"39",
          4950 => x"d4",
          4951 => x"f7",
          4952 => x"af",
          4953 => x"7d",
          4954 => x"73",
          4955 => x"df",
          4956 => x"29",
          4957 => x"05",
          4958 => x"04",
          4959 => x"33",
          4960 => x"2e",
          4961 => x"82",
          4962 => x"55",
          4963 => x"ab",
          4964 => x"2b",
          4965 => x"51",
          4966 => x"24",
          4967 => x"1a",
          4968 => x"81",
          4969 => x"81",
          4970 => x"81",
          4971 => x"70",
          4972 => x"f7",
          4973 => x"51",
          4974 => x"82",
          4975 => x"81",
          4976 => x"74",
          4977 => x"34",
          4978 => x"ae",
          4979 => x"34",
          4980 => x"33",
          4981 => x"25",
          4982 => x"14",
          4983 => x"f7",
          4984 => x"f7",
          4985 => x"81",
          4986 => x"81",
          4987 => x"70",
          4988 => x"f7",
          4989 => x"51",
          4990 => x"77",
          4991 => x"82",
          4992 => x"52",
          4993 => x"33",
          4994 => x"97",
          4995 => x"81",
          4996 => x"81",
          4997 => x"70",
          4998 => x"f7",
          4999 => x"51",
          5000 => x"24",
          5001 => x"f7",
          5002 => x"98",
          5003 => x"2c",
          5004 => x"33",
          5005 => x"56",
          5006 => x"fc",
          5007 => x"fb",
          5008 => x"88",
          5009 => x"a1",
          5010 => x"80",
          5011 => x"80",
          5012 => x"98",
          5013 => x"d8",
          5014 => x"55",
          5015 => x"de",
          5016 => x"39",
          5017 => x"80",
          5018 => x"34",
          5019 => x"53",
          5020 => x"c1",
          5021 => x"9a",
          5022 => x"39",
          5023 => x"33",
          5024 => x"06",
          5025 => x"80",
          5026 => x"38",
          5027 => x"33",
          5028 => x"73",
          5029 => x"34",
          5030 => x"73",
          5031 => x"34",
          5032 => x"08",
          5033 => x"ff",
          5034 => x"82",
          5035 => x"70",
          5036 => x"98",
          5037 => x"d8",
          5038 => x"56",
          5039 => x"25",
          5040 => x"1a",
          5041 => x"33",
          5042 => x"fb",
          5043 => x"73",
          5044 => x"96",
          5045 => x"81",
          5046 => x"81",
          5047 => x"70",
          5048 => x"f7",
          5049 => x"51",
          5050 => x"24",
          5051 => x"fb",
          5052 => x"a0",
          5053 => x"f1",
          5054 => x"dc",
          5055 => x"2b",
          5056 => x"82",
          5057 => x"57",
          5058 => x"74",
          5059 => x"bf",
          5060 => x"fc",
          5061 => x"51",
          5062 => x"3f",
          5063 => x"0a",
          5064 => x"0a",
          5065 => x"2c",
          5066 => x"33",
          5067 => x"75",
          5068 => x"38",
          5069 => x"82",
          5070 => x"7a",
          5071 => x"74",
          5072 => x"fc",
          5073 => x"51",
          5074 => x"3f",
          5075 => x"52",
          5076 => x"c7",
          5077 => x"98",
          5078 => x"06",
          5079 => x"38",
          5080 => x"33",
          5081 => x"2e",
          5082 => x"53",
          5083 => x"51",
          5084 => x"84",
          5085 => x"34",
          5086 => x"f7",
          5087 => x"0b",
          5088 => x"34",
          5089 => x"98",
          5090 => x"0d",
          5091 => x"dc",
          5092 => x"80",
          5093 => x"38",
          5094 => x"08",
          5095 => x"ff",
          5096 => x"82",
          5097 => x"ff",
          5098 => x"82",
          5099 => x"73",
          5100 => x"54",
          5101 => x"f7",
          5102 => x"f7",
          5103 => x"55",
          5104 => x"f9",
          5105 => x"14",
          5106 => x"f7",
          5107 => x"98",
          5108 => x"2c",
          5109 => x"06",
          5110 => x"74",
          5111 => x"38",
          5112 => x"81",
          5113 => x"34",
          5114 => x"08",
          5115 => x"51",
          5116 => x"3f",
          5117 => x"0a",
          5118 => x"0a",
          5119 => x"2c",
          5120 => x"33",
          5121 => x"75",
          5122 => x"38",
          5123 => x"08",
          5124 => x"ff",
          5125 => x"82",
          5126 => x"70",
          5127 => x"98",
          5128 => x"d8",
          5129 => x"56",
          5130 => x"24",
          5131 => x"82",
          5132 => x"52",
          5133 => x"93",
          5134 => x"81",
          5135 => x"81",
          5136 => x"70",
          5137 => x"f7",
          5138 => x"51",
          5139 => x"25",
          5140 => x"fb",
          5141 => x"dc",
          5142 => x"ff",
          5143 => x"d8",
          5144 => x"54",
          5145 => x"f7",
          5146 => x"fb",
          5147 => x"81",
          5148 => x"82",
          5149 => x"74",
          5150 => x"52",
          5151 => x"e9",
          5152 => x"dc",
          5153 => x"ff",
          5154 => x"d8",
          5155 => x"54",
          5156 => x"d6",
          5157 => x"39",
          5158 => x"53",
          5159 => x"c1",
          5160 => x"ee",
          5161 => x"82",
          5162 => x"80",
          5163 => x"d8",
          5164 => x"39",
          5165 => x"82",
          5166 => x"55",
          5167 => x"a6",
          5168 => x"ff",
          5169 => x"82",
          5170 => x"82",
          5171 => x"82",
          5172 => x"81",
          5173 => x"05",
          5174 => x"79",
          5175 => x"bc",
          5176 => x"81",
          5177 => x"84",
          5178 => x"90",
          5179 => x"08",
          5180 => x"80",
          5181 => x"74",
          5182 => x"c0",
          5183 => x"98",
          5184 => x"d8",
          5185 => x"98",
          5186 => x"06",
          5187 => x"74",
          5188 => x"ff",
          5189 => x"ff",
          5190 => x"fa",
          5191 => x"55",
          5192 => x"f6",
          5193 => x"51",
          5194 => x"3f",
          5195 => x"93",
          5196 => x"06",
          5197 => x"df",
          5198 => x"74",
          5199 => x"38",
          5200 => x"99",
          5201 => x"e0",
          5202 => x"f7",
          5203 => x"e0",
          5204 => x"ff",
          5205 => x"53",
          5206 => x"51",
          5207 => x"3f",
          5208 => x"7a",
          5209 => x"df",
          5210 => x"08",
          5211 => x"80",
          5212 => x"74",
          5213 => x"c4",
          5214 => x"98",
          5215 => x"d8",
          5216 => x"98",
          5217 => x"06",
          5218 => x"74",
          5219 => x"ff",
          5220 => x"81",
          5221 => x"81",
          5222 => x"89",
          5223 => x"f7",
          5224 => x"7a",
          5225 => x"dc",
          5226 => x"d8",
          5227 => x"51",
          5228 => x"f5",
          5229 => x"f7",
          5230 => x"81",
          5231 => x"f7",
          5232 => x"56",
          5233 => x"27",
          5234 => x"82",
          5235 => x"52",
          5236 => x"73",
          5237 => x"34",
          5238 => x"33",
          5239 => x"90",
          5240 => x"eb",
          5241 => x"dc",
          5242 => x"80",
          5243 => x"38",
          5244 => x"08",
          5245 => x"ff",
          5246 => x"82",
          5247 => x"ff",
          5248 => x"82",
          5249 => x"f4",
          5250 => x"3d",
          5251 => x"f4",
          5252 => x"88",
          5253 => x"0b",
          5254 => x"23",
          5255 => x"53",
          5256 => x"fa",
          5257 => x"a0",
          5258 => x"e0",
          5259 => x"80",
          5260 => x"34",
          5261 => x"81",
          5262 => x"e0",
          5263 => x"77",
          5264 => x"76",
          5265 => x"82",
          5266 => x"54",
          5267 => x"34",
          5268 => x"34",
          5269 => x"08",
          5270 => x"22",
          5271 => x"80",
          5272 => x"83",
          5273 => x"70",
          5274 => x"51",
          5275 => x"88",
          5276 => x"89",
          5277 => x"e0",
          5278 => x"88",
          5279 => x"88",
          5280 => x"11",
          5281 => x"77",
          5282 => x"76",
          5283 => x"89",
          5284 => x"ff",
          5285 => x"52",
          5286 => x"72",
          5287 => x"fb",
          5288 => x"82",
          5289 => x"ff",
          5290 => x"51",
          5291 => x"e0",
          5292 => x"3d",
          5293 => x"3d",
          5294 => x"05",
          5295 => x"05",
          5296 => x"71",
          5297 => x"88",
          5298 => x"2b",
          5299 => x"83",
          5300 => x"70",
          5301 => x"33",
          5302 => x"07",
          5303 => x"ae",
          5304 => x"81",
          5305 => x"07",
          5306 => x"53",
          5307 => x"54",
          5308 => x"53",
          5309 => x"77",
          5310 => x"18",
          5311 => x"88",
          5312 => x"88",
          5313 => x"70",
          5314 => x"74",
          5315 => x"82",
          5316 => x"70",
          5317 => x"81",
          5318 => x"88",
          5319 => x"83",
          5320 => x"f8",
          5321 => x"56",
          5322 => x"73",
          5323 => x"06",
          5324 => x"54",
          5325 => x"82",
          5326 => x"81",
          5327 => x"72",
          5328 => x"82",
          5329 => x"16",
          5330 => x"34",
          5331 => x"34",
          5332 => x"04",
          5333 => x"82",
          5334 => x"02",
          5335 => x"05",
          5336 => x"2b",
          5337 => x"11",
          5338 => x"33",
          5339 => x"71",
          5340 => x"58",
          5341 => x"55",
          5342 => x"84",
          5343 => x"13",
          5344 => x"2b",
          5345 => x"2a",
          5346 => x"52",
          5347 => x"34",
          5348 => x"34",
          5349 => x"08",
          5350 => x"11",
          5351 => x"33",
          5352 => x"71",
          5353 => x"56",
          5354 => x"72",
          5355 => x"33",
          5356 => x"71",
          5357 => x"70",
          5358 => x"56",
          5359 => x"86",
          5360 => x"87",
          5361 => x"e0",
          5362 => x"70",
          5363 => x"33",
          5364 => x"07",
          5365 => x"ff",
          5366 => x"2a",
          5367 => x"53",
          5368 => x"34",
          5369 => x"34",
          5370 => x"04",
          5371 => x"02",
          5372 => x"82",
          5373 => x"71",
          5374 => x"11",
          5375 => x"12",
          5376 => x"2b",
          5377 => x"29",
          5378 => x"81",
          5379 => x"98",
          5380 => x"2b",
          5381 => x"53",
          5382 => x"56",
          5383 => x"71",
          5384 => x"f6",
          5385 => x"fe",
          5386 => x"e0",
          5387 => x"16",
          5388 => x"12",
          5389 => x"2b",
          5390 => x"07",
          5391 => x"33",
          5392 => x"71",
          5393 => x"70",
          5394 => x"ff",
          5395 => x"52",
          5396 => x"5a",
          5397 => x"05",
          5398 => x"54",
          5399 => x"13",
          5400 => x"13",
          5401 => x"88",
          5402 => x"70",
          5403 => x"33",
          5404 => x"71",
          5405 => x"56",
          5406 => x"72",
          5407 => x"81",
          5408 => x"88",
          5409 => x"81",
          5410 => x"70",
          5411 => x"51",
          5412 => x"72",
          5413 => x"81",
          5414 => x"3d",
          5415 => x"3d",
          5416 => x"88",
          5417 => x"05",
          5418 => x"70",
          5419 => x"11",
          5420 => x"83",
          5421 => x"8b",
          5422 => x"2b",
          5423 => x"59",
          5424 => x"73",
          5425 => x"81",
          5426 => x"88",
          5427 => x"8c",
          5428 => x"22",
          5429 => x"88",
          5430 => x"53",
          5431 => x"73",
          5432 => x"14",
          5433 => x"88",
          5434 => x"70",
          5435 => x"33",
          5436 => x"71",
          5437 => x"56",
          5438 => x"72",
          5439 => x"33",
          5440 => x"71",
          5441 => x"70",
          5442 => x"55",
          5443 => x"82",
          5444 => x"83",
          5445 => x"e0",
          5446 => x"82",
          5447 => x"12",
          5448 => x"2b",
          5449 => x"98",
          5450 => x"87",
          5451 => x"f7",
          5452 => x"82",
          5453 => x"31",
          5454 => x"83",
          5455 => x"70",
          5456 => x"fd",
          5457 => x"e0",
          5458 => x"83",
          5459 => x"82",
          5460 => x"12",
          5461 => x"2b",
          5462 => x"07",
          5463 => x"33",
          5464 => x"71",
          5465 => x"90",
          5466 => x"42",
          5467 => x"5b",
          5468 => x"54",
          5469 => x"8d",
          5470 => x"80",
          5471 => x"fe",
          5472 => x"84",
          5473 => x"33",
          5474 => x"71",
          5475 => x"83",
          5476 => x"11",
          5477 => x"53",
          5478 => x"55",
          5479 => x"34",
          5480 => x"06",
          5481 => x"14",
          5482 => x"88",
          5483 => x"84",
          5484 => x"13",
          5485 => x"2b",
          5486 => x"2a",
          5487 => x"56",
          5488 => x"16",
          5489 => x"16",
          5490 => x"88",
          5491 => x"80",
          5492 => x"34",
          5493 => x"14",
          5494 => x"88",
          5495 => x"84",
          5496 => x"85",
          5497 => x"e0",
          5498 => x"70",
          5499 => x"33",
          5500 => x"07",
          5501 => x"80",
          5502 => x"2a",
          5503 => x"56",
          5504 => x"34",
          5505 => x"34",
          5506 => x"04",
          5507 => x"73",
          5508 => x"88",
          5509 => x"f7",
          5510 => x"80",
          5511 => x"71",
          5512 => x"3f",
          5513 => x"04",
          5514 => x"80",
          5515 => x"f8",
          5516 => x"e0",
          5517 => x"ff",
          5518 => x"e0",
          5519 => x"11",
          5520 => x"33",
          5521 => x"07",
          5522 => x"56",
          5523 => x"ff",
          5524 => x"78",
          5525 => x"38",
          5526 => x"17",
          5527 => x"12",
          5528 => x"2b",
          5529 => x"ff",
          5530 => x"31",
          5531 => x"ff",
          5532 => x"27",
          5533 => x"56",
          5534 => x"79",
          5535 => x"73",
          5536 => x"38",
          5537 => x"5b",
          5538 => x"85",
          5539 => x"88",
          5540 => x"54",
          5541 => x"78",
          5542 => x"2e",
          5543 => x"79",
          5544 => x"76",
          5545 => x"e0",
          5546 => x"70",
          5547 => x"33",
          5548 => x"07",
          5549 => x"ff",
          5550 => x"5a",
          5551 => x"73",
          5552 => x"38",
          5553 => x"54",
          5554 => x"81",
          5555 => x"54",
          5556 => x"81",
          5557 => x"7a",
          5558 => x"06",
          5559 => x"51",
          5560 => x"81",
          5561 => x"80",
          5562 => x"52",
          5563 => x"c6",
          5564 => x"88",
          5565 => x"86",
          5566 => x"12",
          5567 => x"2b",
          5568 => x"07",
          5569 => x"55",
          5570 => x"17",
          5571 => x"ff",
          5572 => x"2a",
          5573 => x"54",
          5574 => x"34",
          5575 => x"06",
          5576 => x"15",
          5577 => x"88",
          5578 => x"2b",
          5579 => x"1e",
          5580 => x"87",
          5581 => x"88",
          5582 => x"88",
          5583 => x"5e",
          5584 => x"54",
          5585 => x"34",
          5586 => x"34",
          5587 => x"08",
          5588 => x"11",
          5589 => x"33",
          5590 => x"71",
          5591 => x"53",
          5592 => x"74",
          5593 => x"86",
          5594 => x"87",
          5595 => x"e0",
          5596 => x"16",
          5597 => x"11",
          5598 => x"33",
          5599 => x"07",
          5600 => x"53",
          5601 => x"56",
          5602 => x"16",
          5603 => x"16",
          5604 => x"88",
          5605 => x"05",
          5606 => x"e0",
          5607 => x"3d",
          5608 => x"3d",
          5609 => x"82",
          5610 => x"84",
          5611 => x"3f",
          5612 => x"80",
          5613 => x"71",
          5614 => x"3f",
          5615 => x"08",
          5616 => x"e0",
          5617 => x"3d",
          5618 => x"3d",
          5619 => x"40",
          5620 => x"42",
          5621 => x"88",
          5622 => x"09",
          5623 => x"38",
          5624 => x"7b",
          5625 => x"51",
          5626 => x"82",
          5627 => x"54",
          5628 => x"7e",
          5629 => x"51",
          5630 => x"7e",
          5631 => x"39",
          5632 => x"8f",
          5633 => x"98",
          5634 => x"ff",
          5635 => x"88",
          5636 => x"31",
          5637 => x"83",
          5638 => x"70",
          5639 => x"11",
          5640 => x"12",
          5641 => x"2b",
          5642 => x"31",
          5643 => x"ff",
          5644 => x"29",
          5645 => x"88",
          5646 => x"33",
          5647 => x"71",
          5648 => x"70",
          5649 => x"44",
          5650 => x"41",
          5651 => x"5b",
          5652 => x"5b",
          5653 => x"25",
          5654 => x"81",
          5655 => x"75",
          5656 => x"ff",
          5657 => x"54",
          5658 => x"83",
          5659 => x"88",
          5660 => x"88",
          5661 => x"33",
          5662 => x"71",
          5663 => x"90",
          5664 => x"47",
          5665 => x"54",
          5666 => x"8b",
          5667 => x"31",
          5668 => x"ff",
          5669 => x"77",
          5670 => x"fe",
          5671 => x"54",
          5672 => x"09",
          5673 => x"38",
          5674 => x"c0",
          5675 => x"ff",
          5676 => x"81",
          5677 => x"8e",
          5678 => x"24",
          5679 => x"51",
          5680 => x"81",
          5681 => x"18",
          5682 => x"24",
          5683 => x"79",
          5684 => x"33",
          5685 => x"71",
          5686 => x"53",
          5687 => x"f4",
          5688 => x"78",
          5689 => x"3f",
          5690 => x"08",
          5691 => x"06",
          5692 => x"53",
          5693 => x"82",
          5694 => x"11",
          5695 => x"55",
          5696 => x"ce",
          5697 => x"88",
          5698 => x"05",
          5699 => x"ff",
          5700 => x"81",
          5701 => x"15",
          5702 => x"24",
          5703 => x"78",
          5704 => x"3f",
          5705 => x"08",
          5706 => x"33",
          5707 => x"71",
          5708 => x"53",
          5709 => x"9c",
          5710 => x"78",
          5711 => x"3f",
          5712 => x"08",
          5713 => x"06",
          5714 => x"53",
          5715 => x"82",
          5716 => x"11",
          5717 => x"55",
          5718 => x"f6",
          5719 => x"88",
          5720 => x"05",
          5721 => x"19",
          5722 => x"83",
          5723 => x"58",
          5724 => x"7f",
          5725 => x"b0",
          5726 => x"98",
          5727 => x"e0",
          5728 => x"2e",
          5729 => x"53",
          5730 => x"e0",
          5731 => x"ff",
          5732 => x"73",
          5733 => x"3f",
          5734 => x"78",
          5735 => x"80",
          5736 => x"78",
          5737 => x"3f",
          5738 => x"2b",
          5739 => x"08",
          5740 => x"51",
          5741 => x"7b",
          5742 => x"e0",
          5743 => x"3d",
          5744 => x"3d",
          5745 => x"29",
          5746 => x"fb",
          5747 => x"e0",
          5748 => x"82",
          5749 => x"80",
          5750 => x"73",
          5751 => x"82",
          5752 => x"51",
          5753 => x"3f",
          5754 => x"98",
          5755 => x"0d",
          5756 => x"0d",
          5757 => x"33",
          5758 => x"70",
          5759 => x"38",
          5760 => x"11",
          5761 => x"82",
          5762 => x"83",
          5763 => x"fc",
          5764 => x"9b",
          5765 => x"84",
          5766 => x"33",
          5767 => x"51",
          5768 => x"80",
          5769 => x"84",
          5770 => x"92",
          5771 => x"51",
          5772 => x"80",
          5773 => x"81",
          5774 => x"72",
          5775 => x"92",
          5776 => x"81",
          5777 => x"0b",
          5778 => x"8c",
          5779 => x"71",
          5780 => x"06",
          5781 => x"80",
          5782 => x"87",
          5783 => x"08",
          5784 => x"38",
          5785 => x"80",
          5786 => x"71",
          5787 => x"c0",
          5788 => x"51",
          5789 => x"87",
          5790 => x"e0",
          5791 => x"82",
          5792 => x"33",
          5793 => x"e0",
          5794 => x"3d",
          5795 => x"3d",
          5796 => x"64",
          5797 => x"bf",
          5798 => x"40",
          5799 => x"74",
          5800 => x"cd",
          5801 => x"98",
          5802 => x"7a",
          5803 => x"81",
          5804 => x"72",
          5805 => x"87",
          5806 => x"11",
          5807 => x"8c",
          5808 => x"92",
          5809 => x"5a",
          5810 => x"58",
          5811 => x"c0",
          5812 => x"76",
          5813 => x"76",
          5814 => x"70",
          5815 => x"81",
          5816 => x"54",
          5817 => x"8e",
          5818 => x"52",
          5819 => x"81",
          5820 => x"81",
          5821 => x"74",
          5822 => x"53",
          5823 => x"83",
          5824 => x"78",
          5825 => x"8f",
          5826 => x"2e",
          5827 => x"c0",
          5828 => x"52",
          5829 => x"87",
          5830 => x"08",
          5831 => x"2e",
          5832 => x"84",
          5833 => x"38",
          5834 => x"87",
          5835 => x"15",
          5836 => x"70",
          5837 => x"52",
          5838 => x"ff",
          5839 => x"39",
          5840 => x"81",
          5841 => x"ff",
          5842 => x"57",
          5843 => x"90",
          5844 => x"80",
          5845 => x"71",
          5846 => x"78",
          5847 => x"38",
          5848 => x"80",
          5849 => x"80",
          5850 => x"81",
          5851 => x"72",
          5852 => x"0c",
          5853 => x"04",
          5854 => x"60",
          5855 => x"8c",
          5856 => x"33",
          5857 => x"5b",
          5858 => x"74",
          5859 => x"e1",
          5860 => x"98",
          5861 => x"79",
          5862 => x"78",
          5863 => x"06",
          5864 => x"77",
          5865 => x"87",
          5866 => x"11",
          5867 => x"8c",
          5868 => x"92",
          5869 => x"59",
          5870 => x"85",
          5871 => x"98",
          5872 => x"7d",
          5873 => x"0c",
          5874 => x"08",
          5875 => x"70",
          5876 => x"53",
          5877 => x"2e",
          5878 => x"70",
          5879 => x"33",
          5880 => x"18",
          5881 => x"2a",
          5882 => x"51",
          5883 => x"2e",
          5884 => x"c0",
          5885 => x"52",
          5886 => x"87",
          5887 => x"08",
          5888 => x"2e",
          5889 => x"84",
          5890 => x"38",
          5891 => x"87",
          5892 => x"15",
          5893 => x"70",
          5894 => x"52",
          5895 => x"ff",
          5896 => x"39",
          5897 => x"81",
          5898 => x"80",
          5899 => x"52",
          5900 => x"90",
          5901 => x"80",
          5902 => x"71",
          5903 => x"7a",
          5904 => x"38",
          5905 => x"80",
          5906 => x"80",
          5907 => x"81",
          5908 => x"72",
          5909 => x"0c",
          5910 => x"04",
          5911 => x"7a",
          5912 => x"a3",
          5913 => x"88",
          5914 => x"33",
          5915 => x"56",
          5916 => x"3f",
          5917 => x"08",
          5918 => x"83",
          5919 => x"fe",
          5920 => x"87",
          5921 => x"0c",
          5922 => x"76",
          5923 => x"38",
          5924 => x"93",
          5925 => x"2b",
          5926 => x"8c",
          5927 => x"71",
          5928 => x"38",
          5929 => x"71",
          5930 => x"c6",
          5931 => x"39",
          5932 => x"81",
          5933 => x"06",
          5934 => x"71",
          5935 => x"38",
          5936 => x"8c",
          5937 => x"e8",
          5938 => x"98",
          5939 => x"71",
          5940 => x"73",
          5941 => x"92",
          5942 => x"72",
          5943 => x"06",
          5944 => x"f7",
          5945 => x"80",
          5946 => x"88",
          5947 => x"0c",
          5948 => x"80",
          5949 => x"56",
          5950 => x"56",
          5951 => x"82",
          5952 => x"88",
          5953 => x"fe",
          5954 => x"81",
          5955 => x"33",
          5956 => x"07",
          5957 => x"0c",
          5958 => x"3d",
          5959 => x"3d",
          5960 => x"11",
          5961 => x"33",
          5962 => x"71",
          5963 => x"81",
          5964 => x"72",
          5965 => x"75",
          5966 => x"82",
          5967 => x"52",
          5968 => x"54",
          5969 => x"0d",
          5970 => x"0d",
          5971 => x"05",
          5972 => x"52",
          5973 => x"70",
          5974 => x"34",
          5975 => x"51",
          5976 => x"83",
          5977 => x"ff",
          5978 => x"75",
          5979 => x"72",
          5980 => x"54",
          5981 => x"2a",
          5982 => x"70",
          5983 => x"34",
          5984 => x"51",
          5985 => x"81",
          5986 => x"70",
          5987 => x"70",
          5988 => x"3d",
          5989 => x"3d",
          5990 => x"77",
          5991 => x"70",
          5992 => x"38",
          5993 => x"05",
          5994 => x"70",
          5995 => x"34",
          5996 => x"eb",
          5997 => x"0d",
          5998 => x"0d",
          5999 => x"54",
          6000 => x"72",
          6001 => x"54",
          6002 => x"51",
          6003 => x"84",
          6004 => x"fc",
          6005 => x"77",
          6006 => x"53",
          6007 => x"05",
          6008 => x"70",
          6009 => x"33",
          6010 => x"ff",
          6011 => x"52",
          6012 => x"2e",
          6013 => x"80",
          6014 => x"71",
          6015 => x"0c",
          6016 => x"04",
          6017 => x"74",
          6018 => x"89",
          6019 => x"2e",
          6020 => x"11",
          6021 => x"52",
          6022 => x"70",
          6023 => x"98",
          6024 => x"0d",
          6025 => x"82",
          6026 => x"04",
          6027 => x"77",
          6028 => x"70",
          6029 => x"33",
          6030 => x"55",
          6031 => x"ff",
          6032 => x"98",
          6033 => x"72",
          6034 => x"38",
          6035 => x"72",
          6036 => x"a2",
          6037 => x"98",
          6038 => x"ff",
          6039 => x"80",
          6040 => x"73",
          6041 => x"55",
          6042 => x"98",
          6043 => x"0d",
          6044 => x"0d",
          6045 => x"0b",
          6046 => x"56",
          6047 => x"2e",
          6048 => x"81",
          6049 => x"08",
          6050 => x"70",
          6051 => x"33",
          6052 => x"e4",
          6053 => x"98",
          6054 => x"09",
          6055 => x"38",
          6056 => x"08",
          6057 => x"b4",
          6058 => x"a8",
          6059 => x"a0",
          6060 => x"56",
          6061 => x"27",
          6062 => x"16",
          6063 => x"82",
          6064 => x"06",
          6065 => x"54",
          6066 => x"78",
          6067 => x"33",
          6068 => x"3f",
          6069 => x"5a",
          6070 => x"98",
          6071 => x"0d",
          6072 => x"0d",
          6073 => x"56",
          6074 => x"b4",
          6075 => x"af",
          6076 => x"fe",
          6077 => x"e0",
          6078 => x"82",
          6079 => x"9f",
          6080 => x"74",
          6081 => x"52",
          6082 => x"51",
          6083 => x"82",
          6084 => x"80",
          6085 => x"ff",
          6086 => x"74",
          6087 => x"76",
          6088 => x"0c",
          6089 => x"04",
          6090 => x"7a",
          6091 => x"fe",
          6092 => x"e0",
          6093 => x"82",
          6094 => x"81",
          6095 => x"33",
          6096 => x"2e",
          6097 => x"80",
          6098 => x"17",
          6099 => x"81",
          6100 => x"06",
          6101 => x"84",
          6102 => x"e0",
          6103 => x"b8",
          6104 => x"56",
          6105 => x"82",
          6106 => x"84",
          6107 => x"fb",
          6108 => x"8b",
          6109 => x"52",
          6110 => x"eb",
          6111 => x"85",
          6112 => x"84",
          6113 => x"fb",
          6114 => x"17",
          6115 => x"a0",
          6116 => x"d3",
          6117 => x"08",
          6118 => x"17",
          6119 => x"3f",
          6120 => x"81",
          6121 => x"19",
          6122 => x"53",
          6123 => x"17",
          6124 => x"c4",
          6125 => x"18",
          6126 => x"80",
          6127 => x"33",
          6128 => x"3f",
          6129 => x"08",
          6130 => x"38",
          6131 => x"82",
          6132 => x"8a",
          6133 => x"fb",
          6134 => x"fe",
          6135 => x"08",
          6136 => x"56",
          6137 => x"74",
          6138 => x"38",
          6139 => x"75",
          6140 => x"16",
          6141 => x"53",
          6142 => x"98",
          6143 => x"0d",
          6144 => x"0d",
          6145 => x"08",
          6146 => x"81",
          6147 => x"df",
          6148 => x"15",
          6149 => x"d7",
          6150 => x"33",
          6151 => x"82",
          6152 => x"38",
          6153 => x"89",
          6154 => x"2e",
          6155 => x"bf",
          6156 => x"2e",
          6157 => x"81",
          6158 => x"81",
          6159 => x"89",
          6160 => x"08",
          6161 => x"52",
          6162 => x"3f",
          6163 => x"08",
          6164 => x"74",
          6165 => x"14",
          6166 => x"81",
          6167 => x"2a",
          6168 => x"05",
          6169 => x"57",
          6170 => x"f5",
          6171 => x"98",
          6172 => x"38",
          6173 => x"06",
          6174 => x"33",
          6175 => x"78",
          6176 => x"06",
          6177 => x"5c",
          6178 => x"53",
          6179 => x"38",
          6180 => x"06",
          6181 => x"39",
          6182 => x"a8",
          6183 => x"52",
          6184 => x"bd",
          6185 => x"98",
          6186 => x"38",
          6187 => x"fe",
          6188 => x"b8",
          6189 => x"cf",
          6190 => x"98",
          6191 => x"ff",
          6192 => x"39",
          6193 => x"a8",
          6194 => x"52",
          6195 => x"91",
          6196 => x"98",
          6197 => x"76",
          6198 => x"fc",
          6199 => x"b8",
          6200 => x"ba",
          6201 => x"98",
          6202 => x"06",
          6203 => x"81",
          6204 => x"e0",
          6205 => x"3d",
          6206 => x"3d",
          6207 => x"7e",
          6208 => x"82",
          6209 => x"27",
          6210 => x"76",
          6211 => x"27",
          6212 => x"75",
          6213 => x"79",
          6214 => x"38",
          6215 => x"89",
          6216 => x"2e",
          6217 => x"80",
          6218 => x"2e",
          6219 => x"81",
          6220 => x"81",
          6221 => x"89",
          6222 => x"08",
          6223 => x"52",
          6224 => x"3f",
          6225 => x"08",
          6226 => x"98",
          6227 => x"38",
          6228 => x"06",
          6229 => x"81",
          6230 => x"06",
          6231 => x"77",
          6232 => x"2e",
          6233 => x"84",
          6234 => x"06",
          6235 => x"06",
          6236 => x"53",
          6237 => x"81",
          6238 => x"34",
          6239 => x"a8",
          6240 => x"52",
          6241 => x"d9",
          6242 => x"98",
          6243 => x"e0",
          6244 => x"94",
          6245 => x"ff",
          6246 => x"05",
          6247 => x"54",
          6248 => x"38",
          6249 => x"74",
          6250 => x"06",
          6251 => x"07",
          6252 => x"74",
          6253 => x"39",
          6254 => x"a8",
          6255 => x"52",
          6256 => x"9d",
          6257 => x"98",
          6258 => x"e0",
          6259 => x"d8",
          6260 => x"ff",
          6261 => x"76",
          6262 => x"06",
          6263 => x"05",
          6264 => x"3f",
          6265 => x"87",
          6266 => x"08",
          6267 => x"51",
          6268 => x"82",
          6269 => x"59",
          6270 => x"08",
          6271 => x"f0",
          6272 => x"82",
          6273 => x"06",
          6274 => x"05",
          6275 => x"54",
          6276 => x"3f",
          6277 => x"08",
          6278 => x"74",
          6279 => x"51",
          6280 => x"81",
          6281 => x"34",
          6282 => x"98",
          6283 => x"0d",
          6284 => x"0d",
          6285 => x"72",
          6286 => x"56",
          6287 => x"27",
          6288 => x"9c",
          6289 => x"9d",
          6290 => x"2e",
          6291 => x"53",
          6292 => x"51",
          6293 => x"82",
          6294 => x"54",
          6295 => x"08",
          6296 => x"93",
          6297 => x"80",
          6298 => x"54",
          6299 => x"82",
          6300 => x"54",
          6301 => x"74",
          6302 => x"fb",
          6303 => x"e0",
          6304 => x"82",
          6305 => x"80",
          6306 => x"38",
          6307 => x"08",
          6308 => x"38",
          6309 => x"08",
          6310 => x"38",
          6311 => x"52",
          6312 => x"d6",
          6313 => x"98",
          6314 => x"9c",
          6315 => x"11",
          6316 => x"57",
          6317 => x"74",
          6318 => x"81",
          6319 => x"0c",
          6320 => x"81",
          6321 => x"84",
          6322 => x"55",
          6323 => x"ff",
          6324 => x"54",
          6325 => x"98",
          6326 => x"0d",
          6327 => x"0d",
          6328 => x"08",
          6329 => x"79",
          6330 => x"17",
          6331 => x"80",
          6332 => x"9c",
          6333 => x"26",
          6334 => x"58",
          6335 => x"52",
          6336 => x"fd",
          6337 => x"74",
          6338 => x"08",
          6339 => x"38",
          6340 => x"08",
          6341 => x"98",
          6342 => x"82",
          6343 => x"17",
          6344 => x"98",
          6345 => x"c7",
          6346 => x"94",
          6347 => x"56",
          6348 => x"2e",
          6349 => x"77",
          6350 => x"81",
          6351 => x"38",
          6352 => x"9c",
          6353 => x"26",
          6354 => x"56",
          6355 => x"51",
          6356 => x"80",
          6357 => x"98",
          6358 => x"09",
          6359 => x"38",
          6360 => x"08",
          6361 => x"98",
          6362 => x"30",
          6363 => x"80",
          6364 => x"07",
          6365 => x"08",
          6366 => x"55",
          6367 => x"ef",
          6368 => x"98",
          6369 => x"95",
          6370 => x"08",
          6371 => x"27",
          6372 => x"9c",
          6373 => x"89",
          6374 => x"85",
          6375 => x"db",
          6376 => x"81",
          6377 => x"17",
          6378 => x"89",
          6379 => x"75",
          6380 => x"ac",
          6381 => x"7a",
          6382 => x"3f",
          6383 => x"08",
          6384 => x"38",
          6385 => x"e0",
          6386 => x"2e",
          6387 => x"86",
          6388 => x"98",
          6389 => x"e0",
          6390 => x"70",
          6391 => x"07",
          6392 => x"7c",
          6393 => x"55",
          6394 => x"f8",
          6395 => x"2e",
          6396 => x"ff",
          6397 => x"55",
          6398 => x"ff",
          6399 => x"76",
          6400 => x"3f",
          6401 => x"08",
          6402 => x"08",
          6403 => x"e0",
          6404 => x"80",
          6405 => x"55",
          6406 => x"94",
          6407 => x"2e",
          6408 => x"53",
          6409 => x"51",
          6410 => x"82",
          6411 => x"55",
          6412 => x"75",
          6413 => x"9c",
          6414 => x"05",
          6415 => x"56",
          6416 => x"26",
          6417 => x"15",
          6418 => x"84",
          6419 => x"07",
          6420 => x"18",
          6421 => x"ff",
          6422 => x"2e",
          6423 => x"39",
          6424 => x"39",
          6425 => x"08",
          6426 => x"81",
          6427 => x"74",
          6428 => x"0c",
          6429 => x"04",
          6430 => x"7a",
          6431 => x"f3",
          6432 => x"e0",
          6433 => x"81",
          6434 => x"98",
          6435 => x"38",
          6436 => x"51",
          6437 => x"82",
          6438 => x"82",
          6439 => x"b4",
          6440 => x"84",
          6441 => x"52",
          6442 => x"52",
          6443 => x"3f",
          6444 => x"39",
          6445 => x"8a",
          6446 => x"75",
          6447 => x"38",
          6448 => x"19",
          6449 => x"81",
          6450 => x"ed",
          6451 => x"e0",
          6452 => x"2e",
          6453 => x"15",
          6454 => x"70",
          6455 => x"07",
          6456 => x"53",
          6457 => x"75",
          6458 => x"0c",
          6459 => x"04",
          6460 => x"7a",
          6461 => x"58",
          6462 => x"f0",
          6463 => x"80",
          6464 => x"9f",
          6465 => x"80",
          6466 => x"90",
          6467 => x"17",
          6468 => x"aa",
          6469 => x"53",
          6470 => x"88",
          6471 => x"08",
          6472 => x"38",
          6473 => x"53",
          6474 => x"17",
          6475 => x"72",
          6476 => x"fe",
          6477 => x"08",
          6478 => x"80",
          6479 => x"16",
          6480 => x"2b",
          6481 => x"75",
          6482 => x"73",
          6483 => x"f5",
          6484 => x"e0",
          6485 => x"82",
          6486 => x"ff",
          6487 => x"81",
          6488 => x"98",
          6489 => x"38",
          6490 => x"82",
          6491 => x"26",
          6492 => x"58",
          6493 => x"73",
          6494 => x"39",
          6495 => x"51",
          6496 => x"82",
          6497 => x"98",
          6498 => x"94",
          6499 => x"17",
          6500 => x"58",
          6501 => x"9a",
          6502 => x"81",
          6503 => x"74",
          6504 => x"98",
          6505 => x"83",
          6506 => x"b8",
          6507 => x"0c",
          6508 => x"82",
          6509 => x"8a",
          6510 => x"f8",
          6511 => x"70",
          6512 => x"08",
          6513 => x"57",
          6514 => x"0a",
          6515 => x"38",
          6516 => x"15",
          6517 => x"08",
          6518 => x"72",
          6519 => x"cb",
          6520 => x"ff",
          6521 => x"81",
          6522 => x"13",
          6523 => x"94",
          6524 => x"74",
          6525 => x"85",
          6526 => x"22",
          6527 => x"73",
          6528 => x"38",
          6529 => x"8a",
          6530 => x"05",
          6531 => x"06",
          6532 => x"8a",
          6533 => x"73",
          6534 => x"3f",
          6535 => x"08",
          6536 => x"81",
          6537 => x"98",
          6538 => x"ff",
          6539 => x"82",
          6540 => x"ff",
          6541 => x"38",
          6542 => x"82",
          6543 => x"26",
          6544 => x"7b",
          6545 => x"98",
          6546 => x"55",
          6547 => x"94",
          6548 => x"73",
          6549 => x"3f",
          6550 => x"08",
          6551 => x"82",
          6552 => x"80",
          6553 => x"38",
          6554 => x"e0",
          6555 => x"2e",
          6556 => x"55",
          6557 => x"08",
          6558 => x"38",
          6559 => x"08",
          6560 => x"fb",
          6561 => x"e0",
          6562 => x"38",
          6563 => x"0c",
          6564 => x"51",
          6565 => x"82",
          6566 => x"98",
          6567 => x"90",
          6568 => x"16",
          6569 => x"15",
          6570 => x"74",
          6571 => x"0c",
          6572 => x"04",
          6573 => x"7b",
          6574 => x"5b",
          6575 => x"52",
          6576 => x"ac",
          6577 => x"98",
          6578 => x"e0",
          6579 => x"ec",
          6580 => x"98",
          6581 => x"17",
          6582 => x"51",
          6583 => x"82",
          6584 => x"54",
          6585 => x"08",
          6586 => x"82",
          6587 => x"9c",
          6588 => x"33",
          6589 => x"72",
          6590 => x"09",
          6591 => x"38",
          6592 => x"e0",
          6593 => x"72",
          6594 => x"55",
          6595 => x"53",
          6596 => x"8e",
          6597 => x"56",
          6598 => x"09",
          6599 => x"38",
          6600 => x"e0",
          6601 => x"81",
          6602 => x"fd",
          6603 => x"e0",
          6604 => x"82",
          6605 => x"80",
          6606 => x"38",
          6607 => x"09",
          6608 => x"38",
          6609 => x"82",
          6610 => x"8b",
          6611 => x"fd",
          6612 => x"9a",
          6613 => x"eb",
          6614 => x"e0",
          6615 => x"ff",
          6616 => x"70",
          6617 => x"53",
          6618 => x"09",
          6619 => x"38",
          6620 => x"eb",
          6621 => x"e0",
          6622 => x"2b",
          6623 => x"72",
          6624 => x"0c",
          6625 => x"04",
          6626 => x"77",
          6627 => x"ff",
          6628 => x"9a",
          6629 => x"55",
          6630 => x"76",
          6631 => x"53",
          6632 => x"09",
          6633 => x"38",
          6634 => x"52",
          6635 => x"eb",
          6636 => x"3d",
          6637 => x"3d",
          6638 => x"80",
          6639 => x"70",
          6640 => x"81",
          6641 => x"74",
          6642 => x"56",
          6643 => x"70",
          6644 => x"ff",
          6645 => x"51",
          6646 => x"38",
          6647 => x"98",
          6648 => x"0d",
          6649 => x"0d",
          6650 => x"59",
          6651 => x"5f",
          6652 => x"70",
          6653 => x"19",
          6654 => x"83",
          6655 => x"19",
          6656 => x"51",
          6657 => x"82",
          6658 => x"5b",
          6659 => x"08",
          6660 => x"9c",
          6661 => x"33",
          6662 => x"86",
          6663 => x"82",
          6664 => x"15",
          6665 => x"70",
          6666 => x"58",
          6667 => x"1a",
          6668 => x"98",
          6669 => x"81",
          6670 => x"81",
          6671 => x"81",
          6672 => x"98",
          6673 => x"ae",
          6674 => x"06",
          6675 => x"53",
          6676 => x"53",
          6677 => x"82",
          6678 => x"77",
          6679 => x"56",
          6680 => x"09",
          6681 => x"38",
          6682 => x"7f",
          6683 => x"81",
          6684 => x"ef",
          6685 => x"2e",
          6686 => x"81",
          6687 => x"86",
          6688 => x"06",
          6689 => x"80",
          6690 => x"8d",
          6691 => x"81",
          6692 => x"90",
          6693 => x"1d",
          6694 => x"5d",
          6695 => x"09",
          6696 => x"9c",
          6697 => x"33",
          6698 => x"2e",
          6699 => x"81",
          6700 => x"1e",
          6701 => x"52",
          6702 => x"3f",
          6703 => x"08",
          6704 => x"06",
          6705 => x"f8",
          6706 => x"70",
          6707 => x"8d",
          6708 => x"51",
          6709 => x"58",
          6710 => x"a8",
          6711 => x"05",
          6712 => x"3f",
          6713 => x"08",
          6714 => x"06",
          6715 => x"2e",
          6716 => x"81",
          6717 => x"c8",
          6718 => x"1a",
          6719 => x"75",
          6720 => x"14",
          6721 => x"75",
          6722 => x"2e",
          6723 => x"b0",
          6724 => x"57",
          6725 => x"c1",
          6726 => x"70",
          6727 => x"81",
          6728 => x"55",
          6729 => x"8e",
          6730 => x"fe",
          6731 => x"73",
          6732 => x"80",
          6733 => x"1c",
          6734 => x"06",
          6735 => x"39",
          6736 => x"72",
          6737 => x"7b",
          6738 => x"51",
          6739 => x"82",
          6740 => x"81",
          6741 => x"72",
          6742 => x"38",
          6743 => x"1a",
          6744 => x"80",
          6745 => x"f8",
          6746 => x"e0",
          6747 => x"82",
          6748 => x"89",
          6749 => x"08",
          6750 => x"86",
          6751 => x"98",
          6752 => x"82",
          6753 => x"90",
          6754 => x"f2",
          6755 => x"70",
          6756 => x"80",
          6757 => x"f6",
          6758 => x"e0",
          6759 => x"82",
          6760 => x"83",
          6761 => x"ff",
          6762 => x"ff",
          6763 => x"0c",
          6764 => x"52",
          6765 => x"a9",
          6766 => x"98",
          6767 => x"e0",
          6768 => x"85",
          6769 => x"08",
          6770 => x"57",
          6771 => x"84",
          6772 => x"39",
          6773 => x"bf",
          6774 => x"ff",
          6775 => x"73",
          6776 => x"75",
          6777 => x"82",
          6778 => x"83",
          6779 => x"06",
          6780 => x"8f",
          6781 => x"73",
          6782 => x"74",
          6783 => x"81",
          6784 => x"38",
          6785 => x"70",
          6786 => x"81",
          6787 => x"55",
          6788 => x"38",
          6789 => x"70",
          6790 => x"54",
          6791 => x"92",
          6792 => x"33",
          6793 => x"06",
          6794 => x"08",
          6795 => x"58",
          6796 => x"7c",
          6797 => x"06",
          6798 => x"8d",
          6799 => x"7d",
          6800 => x"81",
          6801 => x"38",
          6802 => x"9a",
          6803 => x"e5",
          6804 => x"e0",
          6805 => x"ff",
          6806 => x"74",
          6807 => x"76",
          6808 => x"06",
          6809 => x"05",
          6810 => x"75",
          6811 => x"d2",
          6812 => x"77",
          6813 => x"8f",
          6814 => x"98",
          6815 => x"ff",
          6816 => x"80",
          6817 => x"77",
          6818 => x"80",
          6819 => x"51",
          6820 => x"3f",
          6821 => x"08",
          6822 => x"70",
          6823 => x"81",
          6824 => x"80",
          6825 => x"74",
          6826 => x"08",
          6827 => x"06",
          6828 => x"75",
          6829 => x"75",
          6830 => x"2e",
          6831 => x"b3",
          6832 => x"5b",
          6833 => x"ff",
          6834 => x"33",
          6835 => x"70",
          6836 => x"55",
          6837 => x"2e",
          6838 => x"80",
          6839 => x"77",
          6840 => x"22",
          6841 => x"8b",
          6842 => x"70",
          6843 => x"51",
          6844 => x"81",
          6845 => x"5c",
          6846 => x"93",
          6847 => x"f9",
          6848 => x"e0",
          6849 => x"ff",
          6850 => x"7e",
          6851 => x"ab",
          6852 => x"06",
          6853 => x"38",
          6854 => x"19",
          6855 => x"08",
          6856 => x"3f",
          6857 => x"08",
          6858 => x"38",
          6859 => x"ff",
          6860 => x"0c",
          6861 => x"51",
          6862 => x"82",
          6863 => x"58",
          6864 => x"08",
          6865 => x"e8",
          6866 => x"e0",
          6867 => x"3d",
          6868 => x"3d",
          6869 => x"08",
          6870 => x"81",
          6871 => x"5d",
          6872 => x"73",
          6873 => x"73",
          6874 => x"70",
          6875 => x"5d",
          6876 => x"8d",
          6877 => x"70",
          6878 => x"22",
          6879 => x"f0",
          6880 => x"a0",
          6881 => x"92",
          6882 => x"5f",
          6883 => x"3f",
          6884 => x"05",
          6885 => x"54",
          6886 => x"82",
          6887 => x"c0",
          6888 => x"34",
          6889 => x"1c",
          6890 => x"58",
          6891 => x"52",
          6892 => x"e2",
          6893 => x"27",
          6894 => x"7a",
          6895 => x"70",
          6896 => x"06",
          6897 => x"80",
          6898 => x"74",
          6899 => x"06",
          6900 => x"55",
          6901 => x"81",
          6902 => x"07",
          6903 => x"71",
          6904 => x"81",
          6905 => x"56",
          6906 => x"2e",
          6907 => x"84",
          6908 => x"56",
          6909 => x"76",
          6910 => x"38",
          6911 => x"55",
          6912 => x"05",
          6913 => x"57",
          6914 => x"bf",
          6915 => x"74",
          6916 => x"87",
          6917 => x"76",
          6918 => x"ff",
          6919 => x"2a",
          6920 => x"74",
          6921 => x"3d",
          6922 => x"54",
          6923 => x"34",
          6924 => x"b5",
          6925 => x"54",
          6926 => x"ad",
          6927 => x"70",
          6928 => x"e3",
          6929 => x"e0",
          6930 => x"2e",
          6931 => x"17",
          6932 => x"2e",
          6933 => x"15",
          6934 => x"55",
          6935 => x"89",
          6936 => x"70",
          6937 => x"d0",
          6938 => x"77",
          6939 => x"54",
          6940 => x"16",
          6941 => x"56",
          6942 => x"8a",
          6943 => x"81",
          6944 => x"58",
          6945 => x"78",
          6946 => x"27",
          6947 => x"51",
          6948 => x"82",
          6949 => x"8b",
          6950 => x"5b",
          6951 => x"27",
          6952 => x"87",
          6953 => x"e4",
          6954 => x"38",
          6955 => x"08",
          6956 => x"98",
          6957 => x"09",
          6958 => x"df",
          6959 => x"cb",
          6960 => x"1b",
          6961 => x"cb",
          6962 => x"81",
          6963 => x"06",
          6964 => x"81",
          6965 => x"2e",
          6966 => x"52",
          6967 => x"fe",
          6968 => x"82",
          6969 => x"19",
          6970 => x"79",
          6971 => x"3f",
          6972 => x"08",
          6973 => x"98",
          6974 => x"38",
          6975 => x"78",
          6976 => x"d4",
          6977 => x"2b",
          6978 => x"71",
          6979 => x"79",
          6980 => x"3f",
          6981 => x"08",
          6982 => x"98",
          6983 => x"38",
          6984 => x"f5",
          6985 => x"e0",
          6986 => x"ff",
          6987 => x"1a",
          6988 => x"51",
          6989 => x"82",
          6990 => x"57",
          6991 => x"08",
          6992 => x"8c",
          6993 => x"1b",
          6994 => x"ff",
          6995 => x"5b",
          6996 => x"34",
          6997 => x"17",
          6998 => x"98",
          6999 => x"34",
          7000 => x"08",
          7001 => x"51",
          7002 => x"77",
          7003 => x"05",
          7004 => x"73",
          7005 => x"2e",
          7006 => x"10",
          7007 => x"81",
          7008 => x"54",
          7009 => x"d2",
          7010 => x"76",
          7011 => x"b9",
          7012 => x"38",
          7013 => x"54",
          7014 => x"8c",
          7015 => x"38",
          7016 => x"ff",
          7017 => x"74",
          7018 => x"22",
          7019 => x"86",
          7020 => x"c0",
          7021 => x"76",
          7022 => x"83",
          7023 => x"52",
          7024 => x"f7",
          7025 => x"98",
          7026 => x"e0",
          7027 => x"c9",
          7028 => x"59",
          7029 => x"38",
          7030 => x"52",
          7031 => x"81",
          7032 => x"98",
          7033 => x"e0",
          7034 => x"38",
          7035 => x"e0",
          7036 => x"9c",
          7037 => x"df",
          7038 => x"53",
          7039 => x"9c",
          7040 => x"df",
          7041 => x"1a",
          7042 => x"33",
          7043 => x"55",
          7044 => x"34",
          7045 => x"1d",
          7046 => x"74",
          7047 => x"0c",
          7048 => x"04",
          7049 => x"78",
          7050 => x"12",
          7051 => x"08",
          7052 => x"55",
          7053 => x"94",
          7054 => x"74",
          7055 => x"3f",
          7056 => x"08",
          7057 => x"98",
          7058 => x"38",
          7059 => x"52",
          7060 => x"8d",
          7061 => x"98",
          7062 => x"e0",
          7063 => x"38",
          7064 => x"53",
          7065 => x"81",
          7066 => x"34",
          7067 => x"77",
          7068 => x"82",
          7069 => x"52",
          7070 => x"bf",
          7071 => x"98",
          7072 => x"e0",
          7073 => x"2e",
          7074 => x"84",
          7075 => x"06",
          7076 => x"54",
          7077 => x"98",
          7078 => x"0d",
          7079 => x"0d",
          7080 => x"08",
          7081 => x"80",
          7082 => x"34",
          7083 => x"80",
          7084 => x"38",
          7085 => x"ff",
          7086 => x"38",
          7087 => x"7f",
          7088 => x"70",
          7089 => x"5b",
          7090 => x"77",
          7091 => x"38",
          7092 => x"70",
          7093 => x"5b",
          7094 => x"97",
          7095 => x"80",
          7096 => x"ff",
          7097 => x"53",
          7098 => x"26",
          7099 => x"5b",
          7100 => x"76",
          7101 => x"81",
          7102 => x"58",
          7103 => x"b5",
          7104 => x"2b",
          7105 => x"80",
          7106 => x"82",
          7107 => x"83",
          7108 => x"55",
          7109 => x"27",
          7110 => x"76",
          7111 => x"74",
          7112 => x"72",
          7113 => x"97",
          7114 => x"55",
          7115 => x"30",
          7116 => x"78",
          7117 => x"72",
          7118 => x"52",
          7119 => x"80",
          7120 => x"80",
          7121 => x"74",
          7122 => x"55",
          7123 => x"80",
          7124 => x"08",
          7125 => x"70",
          7126 => x"54",
          7127 => x"38",
          7128 => x"80",
          7129 => x"79",
          7130 => x"53",
          7131 => x"05",
          7132 => x"82",
          7133 => x"70",
          7134 => x"5a",
          7135 => x"08",
          7136 => x"81",
          7137 => x"53",
          7138 => x"b7",
          7139 => x"2e",
          7140 => x"84",
          7141 => x"55",
          7142 => x"70",
          7143 => x"07",
          7144 => x"54",
          7145 => x"26",
          7146 => x"80",
          7147 => x"ae",
          7148 => x"05",
          7149 => x"17",
          7150 => x"70",
          7151 => x"34",
          7152 => x"8a",
          7153 => x"b5",
          7154 => x"88",
          7155 => x"0b",
          7156 => x"96",
          7157 => x"72",
          7158 => x"76",
          7159 => x"0b",
          7160 => x"81",
          7161 => x"39",
          7162 => x"1a",
          7163 => x"57",
          7164 => x"80",
          7165 => x"18",
          7166 => x"56",
          7167 => x"bf",
          7168 => x"72",
          7169 => x"38",
          7170 => x"8c",
          7171 => x"53",
          7172 => x"87",
          7173 => x"2a",
          7174 => x"72",
          7175 => x"72",
          7176 => x"72",
          7177 => x"38",
          7178 => x"83",
          7179 => x"56",
          7180 => x"70",
          7181 => x"34",
          7182 => x"15",
          7183 => x"33",
          7184 => x"59",
          7185 => x"38",
          7186 => x"05",
          7187 => x"82",
          7188 => x"1c",
          7189 => x"33",
          7190 => x"85",
          7191 => x"19",
          7192 => x"08",
          7193 => x"33",
          7194 => x"9c",
          7195 => x"11",
          7196 => x"aa",
          7197 => x"98",
          7198 => x"96",
          7199 => x"87",
          7200 => x"98",
          7201 => x"23",
          7202 => x"d8",
          7203 => x"e0",
          7204 => x"19",
          7205 => x"0d",
          7206 => x"0d",
          7207 => x"41",
          7208 => x"70",
          7209 => x"55",
          7210 => x"83",
          7211 => x"73",
          7212 => x"92",
          7213 => x"2e",
          7214 => x"98",
          7215 => x"1f",
          7216 => x"81",
          7217 => x"64",
          7218 => x"56",
          7219 => x"2e",
          7220 => x"83",
          7221 => x"73",
          7222 => x"70",
          7223 => x"25",
          7224 => x"51",
          7225 => x"38",
          7226 => x"0c",
          7227 => x"51",
          7228 => x"26",
          7229 => x"80",
          7230 => x"34",
          7231 => x"51",
          7232 => x"82",
          7233 => x"56",
          7234 => x"63",
          7235 => x"8c",
          7236 => x"54",
          7237 => x"3d",
          7238 => x"da",
          7239 => x"e0",
          7240 => x"2e",
          7241 => x"83",
          7242 => x"82",
          7243 => x"27",
          7244 => x"10",
          7245 => x"98",
          7246 => x"55",
          7247 => x"23",
          7248 => x"82",
          7249 => x"83",
          7250 => x"70",
          7251 => x"30",
          7252 => x"71",
          7253 => x"51",
          7254 => x"73",
          7255 => x"80",
          7256 => x"38",
          7257 => x"26",
          7258 => x"52",
          7259 => x"51",
          7260 => x"82",
          7261 => x"81",
          7262 => x"81",
          7263 => x"d7",
          7264 => x"1a",
          7265 => x"23",
          7266 => x"ff",
          7267 => x"15",
          7268 => x"70",
          7269 => x"57",
          7270 => x"09",
          7271 => x"38",
          7272 => x"80",
          7273 => x"30",
          7274 => x"79",
          7275 => x"54",
          7276 => x"74",
          7277 => x"27",
          7278 => x"78",
          7279 => x"81",
          7280 => x"79",
          7281 => x"ae",
          7282 => x"80",
          7283 => x"82",
          7284 => x"06",
          7285 => x"82",
          7286 => x"73",
          7287 => x"81",
          7288 => x"38",
          7289 => x"73",
          7290 => x"81",
          7291 => x"78",
          7292 => x"80",
          7293 => x"0b",
          7294 => x"58",
          7295 => x"78",
          7296 => x"a0",
          7297 => x"70",
          7298 => x"34",
          7299 => x"8a",
          7300 => x"38",
          7301 => x"54",
          7302 => x"34",
          7303 => x"78",
          7304 => x"38",
          7305 => x"fe",
          7306 => x"22",
          7307 => x"72",
          7308 => x"30",
          7309 => x"51",
          7310 => x"56",
          7311 => x"2e",
          7312 => x"87",
          7313 => x"59",
          7314 => x"78",
          7315 => x"55",
          7316 => x"23",
          7317 => x"86",
          7318 => x"39",
          7319 => x"57",
          7320 => x"80",
          7321 => x"83",
          7322 => x"56",
          7323 => x"a0",
          7324 => x"06",
          7325 => x"1d",
          7326 => x"70",
          7327 => x"5d",
          7328 => x"f2",
          7329 => x"38",
          7330 => x"ff",
          7331 => x"ae",
          7332 => x"06",
          7333 => x"83",
          7334 => x"80",
          7335 => x"79",
          7336 => x"70",
          7337 => x"73",
          7338 => x"38",
          7339 => x"fe",
          7340 => x"19",
          7341 => x"2e",
          7342 => x"15",
          7343 => x"55",
          7344 => x"09",
          7345 => x"38",
          7346 => x"52",
          7347 => x"d5",
          7348 => x"70",
          7349 => x"5f",
          7350 => x"70",
          7351 => x"5f",
          7352 => x"80",
          7353 => x"38",
          7354 => x"96",
          7355 => x"32",
          7356 => x"80",
          7357 => x"54",
          7358 => x"8c",
          7359 => x"2e",
          7360 => x"83",
          7361 => x"39",
          7362 => x"5b",
          7363 => x"83",
          7364 => x"7c",
          7365 => x"30",
          7366 => x"80",
          7367 => x"07",
          7368 => x"55",
          7369 => x"a6",
          7370 => x"2e",
          7371 => x"7c",
          7372 => x"38",
          7373 => x"57",
          7374 => x"81",
          7375 => x"5d",
          7376 => x"7c",
          7377 => x"fc",
          7378 => x"ff",
          7379 => x"ff",
          7380 => x"38",
          7381 => x"57",
          7382 => x"75",
          7383 => x"ae",
          7384 => x"98",
          7385 => x"ff",
          7386 => x"2a",
          7387 => x"51",
          7388 => x"80",
          7389 => x"75",
          7390 => x"82",
          7391 => x"33",
          7392 => x"ff",
          7393 => x"38",
          7394 => x"73",
          7395 => x"38",
          7396 => x"7f",
          7397 => x"c0",
          7398 => x"a0",
          7399 => x"2a",
          7400 => x"75",
          7401 => x"58",
          7402 => x"75",
          7403 => x"38",
          7404 => x"d1",
          7405 => x"cc",
          7406 => x"98",
          7407 => x"8a",
          7408 => x"77",
          7409 => x"56",
          7410 => x"bf",
          7411 => x"99",
          7412 => x"7b",
          7413 => x"ff",
          7414 => x"73",
          7415 => x"38",
          7416 => x"e0",
          7417 => x"ff",
          7418 => x"55",
          7419 => x"a0",
          7420 => x"74",
          7421 => x"58",
          7422 => x"a0",
          7423 => x"73",
          7424 => x"09",
          7425 => x"38",
          7426 => x"1f",
          7427 => x"2e",
          7428 => x"88",
          7429 => x"2b",
          7430 => x"5c",
          7431 => x"54",
          7432 => x"8d",
          7433 => x"06",
          7434 => x"2e",
          7435 => x"85",
          7436 => x"07",
          7437 => x"2a",
          7438 => x"51",
          7439 => x"38",
          7440 => x"54",
          7441 => x"85",
          7442 => x"07",
          7443 => x"2a",
          7444 => x"51",
          7445 => x"2e",
          7446 => x"88",
          7447 => x"ab",
          7448 => x"51",
          7449 => x"82",
          7450 => x"ab",
          7451 => x"56",
          7452 => x"08",
          7453 => x"38",
          7454 => x"08",
          7455 => x"81",
          7456 => x"38",
          7457 => x"70",
          7458 => x"82",
          7459 => x"54",
          7460 => x"96",
          7461 => x"06",
          7462 => x"2e",
          7463 => x"ff",
          7464 => x"1f",
          7465 => x"80",
          7466 => x"81",
          7467 => x"bb",
          7468 => x"b7",
          7469 => x"2a",
          7470 => x"51",
          7471 => x"38",
          7472 => x"70",
          7473 => x"81",
          7474 => x"55",
          7475 => x"e1",
          7476 => x"08",
          7477 => x"60",
          7478 => x"52",
          7479 => x"ef",
          7480 => x"98",
          7481 => x"0c",
          7482 => x"75",
          7483 => x"0c",
          7484 => x"04",
          7485 => x"7c",
          7486 => x"08",
          7487 => x"55",
          7488 => x"59",
          7489 => x"81",
          7490 => x"70",
          7491 => x"33",
          7492 => x"52",
          7493 => x"2e",
          7494 => x"ee",
          7495 => x"2e",
          7496 => x"81",
          7497 => x"33",
          7498 => x"81",
          7499 => x"52",
          7500 => x"26",
          7501 => x"14",
          7502 => x"06",
          7503 => x"52",
          7504 => x"80",
          7505 => x"0b",
          7506 => x"59",
          7507 => x"7a",
          7508 => x"70",
          7509 => x"33",
          7510 => x"05",
          7511 => x"9f",
          7512 => x"53",
          7513 => x"89",
          7514 => x"70",
          7515 => x"54",
          7516 => x"12",
          7517 => x"26",
          7518 => x"12",
          7519 => x"06",
          7520 => x"30",
          7521 => x"51",
          7522 => x"2e",
          7523 => x"85",
          7524 => x"be",
          7525 => x"74",
          7526 => x"30",
          7527 => x"9f",
          7528 => x"2a",
          7529 => x"54",
          7530 => x"2e",
          7531 => x"15",
          7532 => x"55",
          7533 => x"ff",
          7534 => x"39",
          7535 => x"86",
          7536 => x"7c",
          7537 => x"51",
          7538 => x"f7",
          7539 => x"70",
          7540 => x"0c",
          7541 => x"04",
          7542 => x"78",
          7543 => x"83",
          7544 => x"0b",
          7545 => x"79",
          7546 => x"d1",
          7547 => x"55",
          7548 => x"08",
          7549 => x"84",
          7550 => x"ce",
          7551 => x"e0",
          7552 => x"ff",
          7553 => x"83",
          7554 => x"d4",
          7555 => x"81",
          7556 => x"38",
          7557 => x"17",
          7558 => x"74",
          7559 => x"09",
          7560 => x"38",
          7561 => x"81",
          7562 => x"30",
          7563 => x"79",
          7564 => x"54",
          7565 => x"74",
          7566 => x"09",
          7567 => x"38",
          7568 => x"d1",
          7569 => x"ee",
          7570 => x"87",
          7571 => x"98",
          7572 => x"e0",
          7573 => x"2e",
          7574 => x"53",
          7575 => x"52",
          7576 => x"51",
          7577 => x"82",
          7578 => x"55",
          7579 => x"08",
          7580 => x"38",
          7581 => x"82",
          7582 => x"88",
          7583 => x"f2",
          7584 => x"02",
          7585 => x"cb",
          7586 => x"55",
          7587 => x"60",
          7588 => x"3f",
          7589 => x"08",
          7590 => x"80",
          7591 => x"98",
          7592 => x"c7",
          7593 => x"98",
          7594 => x"82",
          7595 => x"70",
          7596 => x"8c",
          7597 => x"2e",
          7598 => x"73",
          7599 => x"81",
          7600 => x"33",
          7601 => x"80",
          7602 => x"81",
          7603 => x"c6",
          7604 => x"e0",
          7605 => x"ff",
          7606 => x"06",
          7607 => x"98",
          7608 => x"2e",
          7609 => x"74",
          7610 => x"81",
          7611 => x"8a",
          7612 => x"f7",
          7613 => x"39",
          7614 => x"77",
          7615 => x"e0",
          7616 => x"81",
          7617 => x"52",
          7618 => x"51",
          7619 => x"82",
          7620 => x"81",
          7621 => x"81",
          7622 => x"83",
          7623 => x"cb",
          7624 => x"2e",
          7625 => x"82",
          7626 => x"06",
          7627 => x"56",
          7628 => x"38",
          7629 => x"74",
          7630 => x"9c",
          7631 => x"98",
          7632 => x"06",
          7633 => x"2e",
          7634 => x"81",
          7635 => x"38",
          7636 => x"19",
          7637 => x"7b",
          7638 => x"38",
          7639 => x"56",
          7640 => x"83",
          7641 => x"70",
          7642 => x"80",
          7643 => x"83",
          7644 => x"cb",
          7645 => x"e0",
          7646 => x"76",
          7647 => x"05",
          7648 => x"16",
          7649 => x"56",
          7650 => x"d7",
          7651 => x"82",
          7652 => x"33",
          7653 => x"9f",
          7654 => x"31",
          7655 => x"84",
          7656 => x"05",
          7657 => x"55",
          7658 => x"08",
          7659 => x"7a",
          7660 => x"38",
          7661 => x"51",
          7662 => x"82",
          7663 => x"81",
          7664 => x"80",
          7665 => x"8d",
          7666 => x"58",
          7667 => x"09",
          7668 => x"38",
          7669 => x"77",
          7670 => x"77",
          7671 => x"38",
          7672 => x"16",
          7673 => x"76",
          7674 => x"81",
          7675 => x"2e",
          7676 => x"8d",
          7677 => x"26",
          7678 => x"80",
          7679 => x"ca",
          7680 => x"e0",
          7681 => x"ff",
          7682 => x"72",
          7683 => x"09",
          7684 => x"d7",
          7685 => x"14",
          7686 => x"3f",
          7687 => x"08",
          7688 => x"06",
          7689 => x"38",
          7690 => x"51",
          7691 => x"82",
          7692 => x"58",
          7693 => x"0c",
          7694 => x"33",
          7695 => x"80",
          7696 => x"ff",
          7697 => x"ff",
          7698 => x"55",
          7699 => x"81",
          7700 => x"38",
          7701 => x"06",
          7702 => x"80",
          7703 => x"52",
          7704 => x"8a",
          7705 => x"80",
          7706 => x"ff",
          7707 => x"53",
          7708 => x"86",
          7709 => x"83",
          7710 => x"c9",
          7711 => x"87",
          7712 => x"98",
          7713 => x"e0",
          7714 => x"15",
          7715 => x"06",
          7716 => x"76",
          7717 => x"80",
          7718 => x"c8",
          7719 => x"e0",
          7720 => x"ff",
          7721 => x"74",
          7722 => x"d8",
          7723 => x"ee",
          7724 => x"98",
          7725 => x"c6",
          7726 => x"cb",
          7727 => x"98",
          7728 => x"ff",
          7729 => x"56",
          7730 => x"83",
          7731 => x"14",
          7732 => x"71",
          7733 => x"5a",
          7734 => x"26",
          7735 => x"8a",
          7736 => x"74",
          7737 => x"fe",
          7738 => x"82",
          7739 => x"55",
          7740 => x"08",
          7741 => x"f3",
          7742 => x"98",
          7743 => x"ff",
          7744 => x"83",
          7745 => x"74",
          7746 => x"26",
          7747 => x"57",
          7748 => x"26",
          7749 => x"57",
          7750 => x"56",
          7751 => x"82",
          7752 => x"15",
          7753 => x"0c",
          7754 => x"0c",
          7755 => x"a8",
          7756 => x"1d",
          7757 => x"54",
          7758 => x"2e",
          7759 => x"af",
          7760 => x"14",
          7761 => x"3f",
          7762 => x"08",
          7763 => x"06",
          7764 => x"72",
          7765 => x"79",
          7766 => x"80",
          7767 => x"c7",
          7768 => x"e0",
          7769 => x"15",
          7770 => x"2b",
          7771 => x"8d",
          7772 => x"2e",
          7773 => x"77",
          7774 => x"0c",
          7775 => x"76",
          7776 => x"38",
          7777 => x"70",
          7778 => x"81",
          7779 => x"53",
          7780 => x"89",
          7781 => x"56",
          7782 => x"08",
          7783 => x"38",
          7784 => x"15",
          7785 => x"90",
          7786 => x"80",
          7787 => x"34",
          7788 => x"09",
          7789 => x"92",
          7790 => x"14",
          7791 => x"3f",
          7792 => x"08",
          7793 => x"06",
          7794 => x"2e",
          7795 => x"80",
          7796 => x"1b",
          7797 => x"ca",
          7798 => x"e0",
          7799 => x"ea",
          7800 => x"98",
          7801 => x"34",
          7802 => x"51",
          7803 => x"82",
          7804 => x"83",
          7805 => x"53",
          7806 => x"d5",
          7807 => x"06",
          7808 => x"b8",
          7809 => x"96",
          7810 => x"98",
          7811 => x"85",
          7812 => x"09",
          7813 => x"38",
          7814 => x"51",
          7815 => x"82",
          7816 => x"86",
          7817 => x"f2",
          7818 => x"06",
          7819 => x"a0",
          7820 => x"ea",
          7821 => x"98",
          7822 => x"0c",
          7823 => x"51",
          7824 => x"82",
          7825 => x"90",
          7826 => x"74",
          7827 => x"f0",
          7828 => x"53",
          7829 => x"f0",
          7830 => x"15",
          7831 => x"f8",
          7832 => x"0c",
          7833 => x"15",
          7834 => x"75",
          7835 => x"0c",
          7836 => x"04",
          7837 => x"77",
          7838 => x"73",
          7839 => x"38",
          7840 => x"72",
          7841 => x"38",
          7842 => x"71",
          7843 => x"38",
          7844 => x"84",
          7845 => x"52",
          7846 => x"09",
          7847 => x"38",
          7848 => x"51",
          7849 => x"3f",
          7850 => x"08",
          7851 => x"71",
          7852 => x"74",
          7853 => x"83",
          7854 => x"78",
          7855 => x"52",
          7856 => x"98",
          7857 => x"0d",
          7858 => x"0d",
          7859 => x"33",
          7860 => x"3d",
          7861 => x"56",
          7862 => x"8b",
          7863 => x"82",
          7864 => x"24",
          7865 => x"e0",
          7866 => x"29",
          7867 => x"05",
          7868 => x"55",
          7869 => x"84",
          7870 => x"34",
          7871 => x"80",
          7872 => x"80",
          7873 => x"75",
          7874 => x"75",
          7875 => x"38",
          7876 => x"3d",
          7877 => x"05",
          7878 => x"3f",
          7879 => x"08",
          7880 => x"e0",
          7881 => x"3d",
          7882 => x"3d",
          7883 => x"84",
          7884 => x"05",
          7885 => x"89",
          7886 => x"2e",
          7887 => x"77",
          7888 => x"54",
          7889 => x"05",
          7890 => x"84",
          7891 => x"f6",
          7892 => x"e0",
          7893 => x"82",
          7894 => x"84",
          7895 => x"5c",
          7896 => x"3d",
          7897 => x"ea",
          7898 => x"e0",
          7899 => x"82",
          7900 => x"92",
          7901 => x"d7",
          7902 => x"98",
          7903 => x"73",
          7904 => x"38",
          7905 => x"9c",
          7906 => x"80",
          7907 => x"38",
          7908 => x"95",
          7909 => x"2e",
          7910 => x"aa",
          7911 => x"df",
          7912 => x"e0",
          7913 => x"9e",
          7914 => x"05",
          7915 => x"54",
          7916 => x"38",
          7917 => x"70",
          7918 => x"54",
          7919 => x"8e",
          7920 => x"83",
          7921 => x"88",
          7922 => x"83",
          7923 => x"83",
          7924 => x"06",
          7925 => x"80",
          7926 => x"38",
          7927 => x"51",
          7928 => x"82",
          7929 => x"56",
          7930 => x"0a",
          7931 => x"05",
          7932 => x"3f",
          7933 => x"0b",
          7934 => x"80",
          7935 => x"7a",
          7936 => x"3f",
          7937 => x"9c",
          7938 => x"db",
          7939 => x"81",
          7940 => x"34",
          7941 => x"80",
          7942 => x"b4",
          7943 => x"54",
          7944 => x"52",
          7945 => x"05",
          7946 => x"3f",
          7947 => x"08",
          7948 => x"98",
          7949 => x"38",
          7950 => x"82",
          7951 => x"b2",
          7952 => x"84",
          7953 => x"06",
          7954 => x"73",
          7955 => x"38",
          7956 => x"ad",
          7957 => x"2a",
          7958 => x"51",
          7959 => x"2e",
          7960 => x"81",
          7961 => x"80",
          7962 => x"87",
          7963 => x"39",
          7964 => x"51",
          7965 => x"82",
          7966 => x"7b",
          7967 => x"12",
          7968 => x"82",
          7969 => x"81",
          7970 => x"83",
          7971 => x"06",
          7972 => x"80",
          7973 => x"77",
          7974 => x"58",
          7975 => x"08",
          7976 => x"63",
          7977 => x"63",
          7978 => x"57",
          7979 => x"82",
          7980 => x"82",
          7981 => x"88",
          7982 => x"9c",
          7983 => x"c0",
          7984 => x"e0",
          7985 => x"e0",
          7986 => x"1b",
          7987 => x"0c",
          7988 => x"22",
          7989 => x"77",
          7990 => x"80",
          7991 => x"34",
          7992 => x"1a",
          7993 => x"94",
          7994 => x"85",
          7995 => x"06",
          7996 => x"80",
          7997 => x"38",
          7998 => x"08",
          7999 => x"84",
          8000 => x"98",
          8001 => x"0c",
          8002 => x"70",
          8003 => x"52",
          8004 => x"39",
          8005 => x"51",
          8006 => x"82",
          8007 => x"57",
          8008 => x"08",
          8009 => x"38",
          8010 => x"e0",
          8011 => x"2e",
          8012 => x"83",
          8013 => x"75",
          8014 => x"74",
          8015 => x"07",
          8016 => x"54",
          8017 => x"8a",
          8018 => x"75",
          8019 => x"73",
          8020 => x"98",
          8021 => x"a9",
          8022 => x"ff",
          8023 => x"80",
          8024 => x"76",
          8025 => x"c4",
          8026 => x"e0",
          8027 => x"38",
          8028 => x"39",
          8029 => x"82",
          8030 => x"05",
          8031 => x"84",
          8032 => x"0c",
          8033 => x"82",
          8034 => x"98",
          8035 => x"f2",
          8036 => x"63",
          8037 => x"40",
          8038 => x"7e",
          8039 => x"fc",
          8040 => x"51",
          8041 => x"82",
          8042 => x"55",
          8043 => x"08",
          8044 => x"19",
          8045 => x"80",
          8046 => x"74",
          8047 => x"39",
          8048 => x"81",
          8049 => x"56",
          8050 => x"82",
          8051 => x"39",
          8052 => x"1a",
          8053 => x"82",
          8054 => x"0b",
          8055 => x"81",
          8056 => x"39",
          8057 => x"94",
          8058 => x"55",
          8059 => x"83",
          8060 => x"7b",
          8061 => x"8c",
          8062 => x"08",
          8063 => x"06",
          8064 => x"81",
          8065 => x"8a",
          8066 => x"05",
          8067 => x"06",
          8068 => x"a8",
          8069 => x"38",
          8070 => x"55",
          8071 => x"19",
          8072 => x"51",
          8073 => x"82",
          8074 => x"55",
          8075 => x"ff",
          8076 => x"ff",
          8077 => x"38",
          8078 => x"0c",
          8079 => x"52",
          8080 => x"93",
          8081 => x"98",
          8082 => x"ff",
          8083 => x"e0",
          8084 => x"7c",
          8085 => x"57",
          8086 => x"80",
          8087 => x"1a",
          8088 => x"22",
          8089 => x"75",
          8090 => x"38",
          8091 => x"58",
          8092 => x"53",
          8093 => x"1b",
          8094 => x"b8",
          8095 => x"e0",
          8096 => x"d6",
          8097 => x"11",
          8098 => x"74",
          8099 => x"38",
          8100 => x"77",
          8101 => x"78",
          8102 => x"84",
          8103 => x"16",
          8104 => x"08",
          8105 => x"2b",
          8106 => x"ff",
          8107 => x"77",
          8108 => x"ba",
          8109 => x"1a",
          8110 => x"08",
          8111 => x"84",
          8112 => x"57",
          8113 => x"27",
          8114 => x"56",
          8115 => x"52",
          8116 => x"8d",
          8117 => x"98",
          8118 => x"38",
          8119 => x"19",
          8120 => x"06",
          8121 => x"52",
          8122 => x"bd",
          8123 => x"76",
          8124 => x"17",
          8125 => x"1e",
          8126 => x"18",
          8127 => x"5e",
          8128 => x"39",
          8129 => x"82",
          8130 => x"90",
          8131 => x"f2",
          8132 => x"63",
          8133 => x"40",
          8134 => x"7e",
          8135 => x"fc",
          8136 => x"51",
          8137 => x"82",
          8138 => x"55",
          8139 => x"08",
          8140 => x"18",
          8141 => x"80",
          8142 => x"74",
          8143 => x"39",
          8144 => x"70",
          8145 => x"81",
          8146 => x"56",
          8147 => x"80",
          8148 => x"38",
          8149 => x"0b",
          8150 => x"82",
          8151 => x"39",
          8152 => x"19",
          8153 => x"83",
          8154 => x"18",
          8155 => x"56",
          8156 => x"27",
          8157 => x"09",
          8158 => x"2e",
          8159 => x"94",
          8160 => x"83",
          8161 => x"56",
          8162 => x"38",
          8163 => x"22",
          8164 => x"89",
          8165 => x"55",
          8166 => x"75",
          8167 => x"18",
          8168 => x"9c",
          8169 => x"85",
          8170 => x"08",
          8171 => x"c6",
          8172 => x"e0",
          8173 => x"82",
          8174 => x"80",
          8175 => x"38",
          8176 => x"ff",
          8177 => x"ff",
          8178 => x"38",
          8179 => x"0c",
          8180 => x"85",
          8181 => x"19",
          8182 => x"b4",
          8183 => x"19",
          8184 => x"81",
          8185 => x"74",
          8186 => x"85",
          8187 => x"98",
          8188 => x"38",
          8189 => x"52",
          8190 => x"bf",
          8191 => x"e0",
          8192 => x"2e",
          8193 => x"82",
          8194 => x"1b",
          8195 => x"5a",
          8196 => x"2e",
          8197 => x"78",
          8198 => x"11",
          8199 => x"55",
          8200 => x"85",
          8201 => x"31",
          8202 => x"76",
          8203 => x"81",
          8204 => x"ff",
          8205 => x"82",
          8206 => x"fe",
          8207 => x"b4",
          8208 => x"31",
          8209 => x"79",
          8210 => x"84",
          8211 => x"16",
          8212 => x"89",
          8213 => x"52",
          8214 => x"ff",
          8215 => x"7e",
          8216 => x"83",
          8217 => x"89",
          8218 => x"de",
          8219 => x"08",
          8220 => x"26",
          8221 => x"51",
          8222 => x"3f",
          8223 => x"08",
          8224 => x"7e",
          8225 => x"0c",
          8226 => x"19",
          8227 => x"08",
          8228 => x"84",
          8229 => x"57",
          8230 => x"27",
          8231 => x"56",
          8232 => x"52",
          8233 => x"bc",
          8234 => x"e0",
          8235 => x"b0",
          8236 => x"7c",
          8237 => x"08",
          8238 => x"1f",
          8239 => x"ff",
          8240 => x"7e",
          8241 => x"83",
          8242 => x"76",
          8243 => x"17",
          8244 => x"1e",
          8245 => x"18",
          8246 => x"0c",
          8247 => x"58",
          8248 => x"74",
          8249 => x"38",
          8250 => x"8c",
          8251 => x"89",
          8252 => x"33",
          8253 => x"55",
          8254 => x"34",
          8255 => x"82",
          8256 => x"90",
          8257 => x"f8",
          8258 => x"8b",
          8259 => x"53",
          8260 => x"f2",
          8261 => x"e0",
          8262 => x"82",
          8263 => x"81",
          8264 => x"16",
          8265 => x"2a",
          8266 => x"51",
          8267 => x"80",
          8268 => x"38",
          8269 => x"52",
          8270 => x"bb",
          8271 => x"e0",
          8272 => x"82",
          8273 => x"80",
          8274 => x"16",
          8275 => x"33",
          8276 => x"55",
          8277 => x"34",
          8278 => x"53",
          8279 => x"08",
          8280 => x"3f",
          8281 => x"52",
          8282 => x"ff",
          8283 => x"82",
          8284 => x"52",
          8285 => x"ff",
          8286 => x"76",
          8287 => x"51",
          8288 => x"3f",
          8289 => x"0b",
          8290 => x"78",
          8291 => x"98",
          8292 => x"98",
          8293 => x"33",
          8294 => x"55",
          8295 => x"17",
          8296 => x"e0",
          8297 => x"3d",
          8298 => x"3d",
          8299 => x"52",
          8300 => x"3f",
          8301 => x"08",
          8302 => x"98",
          8303 => x"86",
          8304 => x"52",
          8305 => x"ac",
          8306 => x"98",
          8307 => x"e0",
          8308 => x"38",
          8309 => x"08",
          8310 => x"82",
          8311 => x"86",
          8312 => x"ff",
          8313 => x"3d",
          8314 => x"3f",
          8315 => x"0b",
          8316 => x"08",
          8317 => x"82",
          8318 => x"82",
          8319 => x"80",
          8320 => x"e0",
          8321 => x"3d",
          8322 => x"3d",
          8323 => x"94",
          8324 => x"52",
          8325 => x"e8",
          8326 => x"e0",
          8327 => x"82",
          8328 => x"80",
          8329 => x"58",
          8330 => x"3d",
          8331 => x"dc",
          8332 => x"e0",
          8333 => x"82",
          8334 => x"bc",
          8335 => x"c7",
          8336 => x"98",
          8337 => x"73",
          8338 => x"38",
          8339 => x"12",
          8340 => x"39",
          8341 => x"33",
          8342 => x"70",
          8343 => x"55",
          8344 => x"2e",
          8345 => x"7f",
          8346 => x"54",
          8347 => x"82",
          8348 => x"98",
          8349 => x"39",
          8350 => x"08",
          8351 => x"81",
          8352 => x"85",
          8353 => x"e0",
          8354 => x"3d",
          8355 => x"a3",
          8356 => x"e1",
          8357 => x"e1",
          8358 => x"5b",
          8359 => x"80",
          8360 => x"3d",
          8361 => x"52",
          8362 => x"51",
          8363 => x"82",
          8364 => x"57",
          8365 => x"08",
          8366 => x"7b",
          8367 => x"0c",
          8368 => x"11",
          8369 => x"3d",
          8370 => x"80",
          8371 => x"54",
          8372 => x"82",
          8373 => x"52",
          8374 => x"70",
          8375 => x"90",
          8376 => x"98",
          8377 => x"e0",
          8378 => x"ef",
          8379 => x"3d",
          8380 => x"51",
          8381 => x"3f",
          8382 => x"08",
          8383 => x"98",
          8384 => x"38",
          8385 => x"08",
          8386 => x"c8",
          8387 => x"e0",
          8388 => x"d6",
          8389 => x"52",
          8390 => x"d4",
          8391 => x"98",
          8392 => x"e0",
          8393 => x"b3",
          8394 => x"74",
          8395 => x"3f",
          8396 => x"08",
          8397 => x"98",
          8398 => x"80",
          8399 => x"52",
          8400 => x"8b",
          8401 => x"e0",
          8402 => x"a6",
          8403 => x"74",
          8404 => x"3f",
          8405 => x"08",
          8406 => x"98",
          8407 => x"c9",
          8408 => x"2e",
          8409 => x"86",
          8410 => x"81",
          8411 => x"81",
          8412 => x"df",
          8413 => x"05",
          8414 => x"d6",
          8415 => x"93",
          8416 => x"82",
          8417 => x"56",
          8418 => x"80",
          8419 => x"02",
          8420 => x"55",
          8421 => x"16",
          8422 => x"56",
          8423 => x"38",
          8424 => x"73",
          8425 => x"99",
          8426 => x"2e",
          8427 => x"16",
          8428 => x"ff",
          8429 => x"3d",
          8430 => x"18",
          8431 => x"58",
          8432 => x"33",
          8433 => x"eb",
          8434 => x"80",
          8435 => x"11",
          8436 => x"74",
          8437 => x"39",
          8438 => x"09",
          8439 => x"38",
          8440 => x"e1",
          8441 => x"55",
          8442 => x"34",
          8443 => x"f7",
          8444 => x"84",
          8445 => x"98",
          8446 => x"70",
          8447 => x"56",
          8448 => x"76",
          8449 => x"81",
          8450 => x"70",
          8451 => x"56",
          8452 => x"82",
          8453 => x"78",
          8454 => x"80",
          8455 => x"27",
          8456 => x"19",
          8457 => x"7a",
          8458 => x"5c",
          8459 => x"55",
          8460 => x"7a",
          8461 => x"5c",
          8462 => x"2e",
          8463 => x"85",
          8464 => x"97",
          8465 => x"3d",
          8466 => x"19",
          8467 => x"33",
          8468 => x"05",
          8469 => x"78",
          8470 => x"80",
          8471 => x"82",
          8472 => x"80",
          8473 => x"04",
          8474 => x"7b",
          8475 => x"fc",
          8476 => x"53",
          8477 => x"fc",
          8478 => x"98",
          8479 => x"e0",
          8480 => x"fe",
          8481 => x"33",
          8482 => x"f6",
          8483 => x"08",
          8484 => x"27",
          8485 => x"15",
          8486 => x"2a",
          8487 => x"51",
          8488 => x"83",
          8489 => x"94",
          8490 => x"80",
          8491 => x"0c",
          8492 => x"2e",
          8493 => x"79",
          8494 => x"70",
          8495 => x"51",
          8496 => x"2e",
          8497 => x"52",
          8498 => x"fe",
          8499 => x"82",
          8500 => x"ff",
          8501 => x"70",
          8502 => x"fe",
          8503 => x"82",
          8504 => x"73",
          8505 => x"76",
          8506 => x"06",
          8507 => x"0c",
          8508 => x"98",
          8509 => x"58",
          8510 => x"39",
          8511 => x"54",
          8512 => x"73",
          8513 => x"ff",
          8514 => x"82",
          8515 => x"54",
          8516 => x"08",
          8517 => x"9d",
          8518 => x"98",
          8519 => x"81",
          8520 => x"e0",
          8521 => x"16",
          8522 => x"16",
          8523 => x"2e",
          8524 => x"76",
          8525 => x"de",
          8526 => x"31",
          8527 => x"18",
          8528 => x"90",
          8529 => x"81",
          8530 => x"06",
          8531 => x"56",
          8532 => x"9b",
          8533 => x"74",
          8534 => x"81",
          8535 => x"98",
          8536 => x"e0",
          8537 => x"38",
          8538 => x"08",
          8539 => x"73",
          8540 => x"ff",
          8541 => x"82",
          8542 => x"54",
          8543 => x"bf",
          8544 => x"27",
          8545 => x"53",
          8546 => x"08",
          8547 => x"73",
          8548 => x"ff",
          8549 => x"15",
          8550 => x"16",
          8551 => x"ff",
          8552 => x"80",
          8553 => x"73",
          8554 => x"ff",
          8555 => x"82",
          8556 => x"94",
          8557 => x"91",
          8558 => x"53",
          8559 => x"81",
          8560 => x"34",
          8561 => x"39",
          8562 => x"82",
          8563 => x"05",
          8564 => x"08",
          8565 => x"08",
          8566 => x"38",
          8567 => x"0c",
          8568 => x"80",
          8569 => x"72",
          8570 => x"73",
          8571 => x"53",
          8572 => x"8c",
          8573 => x"16",
          8574 => x"38",
          8575 => x"0c",
          8576 => x"82",
          8577 => x"8b",
          8578 => x"f9",
          8579 => x"56",
          8580 => x"80",
          8581 => x"38",
          8582 => x"3d",
          8583 => x"8a",
          8584 => x"51",
          8585 => x"82",
          8586 => x"55",
          8587 => x"08",
          8588 => x"77",
          8589 => x"52",
          8590 => x"dd",
          8591 => x"98",
          8592 => x"e0",
          8593 => x"c4",
          8594 => x"33",
          8595 => x"55",
          8596 => x"24",
          8597 => x"16",
          8598 => x"2a",
          8599 => x"51",
          8600 => x"80",
          8601 => x"9c",
          8602 => x"77",
          8603 => x"3f",
          8604 => x"08",
          8605 => x"77",
          8606 => x"22",
          8607 => x"74",
          8608 => x"ff",
          8609 => x"82",
          8610 => x"55",
          8611 => x"09",
          8612 => x"38",
          8613 => x"39",
          8614 => x"84",
          8615 => x"0c",
          8616 => x"82",
          8617 => x"89",
          8618 => x"fc",
          8619 => x"87",
          8620 => x"53",
          8621 => x"e7",
          8622 => x"e0",
          8623 => x"38",
          8624 => x"08",
          8625 => x"3d",
          8626 => x"3d",
          8627 => x"89",
          8628 => x"54",
          8629 => x"54",
          8630 => x"82",
          8631 => x"53",
          8632 => x"08",
          8633 => x"74",
          8634 => x"e0",
          8635 => x"73",
          8636 => x"fc",
          8637 => x"98",
          8638 => x"cb",
          8639 => x"98",
          8640 => x"51",
          8641 => x"82",
          8642 => x"53",
          8643 => x"08",
          8644 => x"81",
          8645 => x"80",
          8646 => x"82",
          8647 => x"a7",
          8648 => x"73",
          8649 => x"3f",
          8650 => x"51",
          8651 => x"3f",
          8652 => x"08",
          8653 => x"30",
          8654 => x"9f",
          8655 => x"e0",
          8656 => x"51",
          8657 => x"72",
          8658 => x"0c",
          8659 => x"04",
          8660 => x"66",
          8661 => x"89",
          8662 => x"97",
          8663 => x"de",
          8664 => x"e0",
          8665 => x"82",
          8666 => x"b2",
          8667 => x"75",
          8668 => x"3f",
          8669 => x"08",
          8670 => x"98",
          8671 => x"02",
          8672 => x"33",
          8673 => x"55",
          8674 => x"25",
          8675 => x"55",
          8676 => x"80",
          8677 => x"76",
          8678 => x"ce",
          8679 => x"82",
          8680 => x"95",
          8681 => x"f0",
          8682 => x"65",
          8683 => x"53",
          8684 => x"05",
          8685 => x"51",
          8686 => x"82",
          8687 => x"5b",
          8688 => x"08",
          8689 => x"7c",
          8690 => x"08",
          8691 => x"fe",
          8692 => x"08",
          8693 => x"55",
          8694 => x"91",
          8695 => x"0c",
          8696 => x"81",
          8697 => x"39",
          8698 => x"c9",
          8699 => x"98",
          8700 => x"55",
          8701 => x"2e",
          8702 => x"80",
          8703 => x"75",
          8704 => x"52",
          8705 => x"05",
          8706 => x"f5",
          8707 => x"98",
          8708 => x"cf",
          8709 => x"98",
          8710 => x"cc",
          8711 => x"98",
          8712 => x"82",
          8713 => x"07",
          8714 => x"05",
          8715 => x"53",
          8716 => x"9c",
          8717 => x"26",
          8718 => x"f9",
          8719 => x"08",
          8720 => x"08",
          8721 => x"98",
          8722 => x"81",
          8723 => x"58",
          8724 => x"3f",
          8725 => x"08",
          8726 => x"98",
          8727 => x"38",
          8728 => x"77",
          8729 => x"5d",
          8730 => x"74",
          8731 => x"81",
          8732 => x"b8",
          8733 => x"a9",
          8734 => x"e0",
          8735 => x"ff",
          8736 => x"30",
          8737 => x"1b",
          8738 => x"5b",
          8739 => x"39",
          8740 => x"ff",
          8741 => x"82",
          8742 => x"f0",
          8743 => x"30",
          8744 => x"1b",
          8745 => x"5b",
          8746 => x"83",
          8747 => x"58",
          8748 => x"92",
          8749 => x"0c",
          8750 => x"12",
          8751 => x"33",
          8752 => x"54",
          8753 => x"34",
          8754 => x"98",
          8755 => x"0d",
          8756 => x"0d",
          8757 => x"fc",
          8758 => x"52",
          8759 => x"3f",
          8760 => x"08",
          8761 => x"98",
          8762 => x"38",
          8763 => x"56",
          8764 => x"38",
          8765 => x"70",
          8766 => x"81",
          8767 => x"55",
          8768 => x"80",
          8769 => x"38",
          8770 => x"54",
          8771 => x"08",
          8772 => x"38",
          8773 => x"82",
          8774 => x"53",
          8775 => x"52",
          8776 => x"b2",
          8777 => x"e0",
          8778 => x"88",
          8779 => x"80",
          8780 => x"17",
          8781 => x"51",
          8782 => x"3f",
          8783 => x"08",
          8784 => x"81",
          8785 => x"81",
          8786 => x"98",
          8787 => x"09",
          8788 => x"38",
          8789 => x"39",
          8790 => x"77",
          8791 => x"98",
          8792 => x"08",
          8793 => x"98",
          8794 => x"82",
          8795 => x"52",
          8796 => x"b1",
          8797 => x"e0",
          8798 => x"94",
          8799 => x"18",
          8800 => x"33",
          8801 => x"54",
          8802 => x"34",
          8803 => x"85",
          8804 => x"18",
          8805 => x"74",
          8806 => x"0c",
          8807 => x"04",
          8808 => x"82",
          8809 => x"ff",
          8810 => x"a3",
          8811 => x"cf",
          8812 => x"98",
          8813 => x"e0",
          8814 => x"f9",
          8815 => x"a3",
          8816 => x"96",
          8817 => x"58",
          8818 => x"82",
          8819 => x"55",
          8820 => x"08",
          8821 => x"02",
          8822 => x"33",
          8823 => x"70",
          8824 => x"55",
          8825 => x"73",
          8826 => x"75",
          8827 => x"80",
          8828 => x"c1",
          8829 => x"da",
          8830 => x"81",
          8831 => x"87",
          8832 => x"b1",
          8833 => x"78",
          8834 => x"c3",
          8835 => x"98",
          8836 => x"2a",
          8837 => x"51",
          8838 => x"80",
          8839 => x"38",
          8840 => x"e0",
          8841 => x"15",
          8842 => x"89",
          8843 => x"82",
          8844 => x"5c",
          8845 => x"3d",
          8846 => x"ff",
          8847 => x"82",
          8848 => x"55",
          8849 => x"08",
          8850 => x"82",
          8851 => x"52",
          8852 => x"bb",
          8853 => x"e0",
          8854 => x"82",
          8855 => x"86",
          8856 => x"80",
          8857 => x"e0",
          8858 => x"2e",
          8859 => x"e0",
          8860 => x"c1",
          8861 => x"c7",
          8862 => x"e0",
          8863 => x"e0",
          8864 => x"70",
          8865 => x"08",
          8866 => x"51",
          8867 => x"80",
          8868 => x"73",
          8869 => x"38",
          8870 => x"52",
          8871 => x"af",
          8872 => x"e0",
          8873 => x"74",
          8874 => x"51",
          8875 => x"3f",
          8876 => x"08",
          8877 => x"e0",
          8878 => x"3d",
          8879 => x"3d",
          8880 => x"9a",
          8881 => x"05",
          8882 => x"51",
          8883 => x"82",
          8884 => x"54",
          8885 => x"08",
          8886 => x"78",
          8887 => x"8e",
          8888 => x"58",
          8889 => x"82",
          8890 => x"54",
          8891 => x"08",
          8892 => x"54",
          8893 => x"82",
          8894 => x"84",
          8895 => x"06",
          8896 => x"02",
          8897 => x"33",
          8898 => x"81",
          8899 => x"86",
          8900 => x"fd",
          8901 => x"74",
          8902 => x"70",
          8903 => x"af",
          8904 => x"e0",
          8905 => x"55",
          8906 => x"98",
          8907 => x"87",
          8908 => x"98",
          8909 => x"09",
          8910 => x"38",
          8911 => x"e0",
          8912 => x"2e",
          8913 => x"86",
          8914 => x"81",
          8915 => x"81",
          8916 => x"e0",
          8917 => x"78",
          8918 => x"9c",
          8919 => x"98",
          8920 => x"e0",
          8921 => x"9f",
          8922 => x"a0",
          8923 => x"51",
          8924 => x"3f",
          8925 => x"0b",
          8926 => x"78",
          8927 => x"80",
          8928 => x"82",
          8929 => x"52",
          8930 => x"51",
          8931 => x"3f",
          8932 => x"b8",
          8933 => x"ff",
          8934 => x"a0",
          8935 => x"11",
          8936 => x"05",
          8937 => x"ee",
          8938 => x"ae",
          8939 => x"15",
          8940 => x"78",
          8941 => x"53",
          8942 => x"cc",
          8943 => x"81",
          8944 => x"34",
          8945 => x"bf",
          8946 => x"e0",
          8947 => x"82",
          8948 => x"b3",
          8949 => x"b2",
          8950 => x"96",
          8951 => x"a3",
          8952 => x"53",
          8953 => x"51",
          8954 => x"3f",
          8955 => x"0b",
          8956 => x"78",
          8957 => x"83",
          8958 => x"51",
          8959 => x"3f",
          8960 => x"08",
          8961 => x"80",
          8962 => x"76",
          8963 => x"a1",
          8964 => x"e0",
          8965 => x"3d",
          8966 => x"3d",
          8967 => x"84",
          8968 => x"d0",
          8969 => x"aa",
          8970 => x"05",
          8971 => x"51",
          8972 => x"82",
          8973 => x"55",
          8974 => x"08",
          8975 => x"78",
          8976 => x"08",
          8977 => x"70",
          8978 => x"cd",
          8979 => x"98",
          8980 => x"e0",
          8981 => x"be",
          8982 => x"9f",
          8983 => x"a0",
          8984 => x"55",
          8985 => x"38",
          8986 => x"3d",
          8987 => x"3d",
          8988 => x"51",
          8989 => x"3f",
          8990 => x"52",
          8991 => x"52",
          8992 => x"92",
          8993 => x"08",
          8994 => x"c8",
          8995 => x"e0",
          8996 => x"82",
          8997 => x"97",
          8998 => x"3d",
          8999 => x"81",
          9000 => x"65",
          9001 => x"2e",
          9002 => x"55",
          9003 => x"82",
          9004 => x"84",
          9005 => x"06",
          9006 => x"73",
          9007 => x"92",
          9008 => x"98",
          9009 => x"e0",
          9010 => x"ca",
          9011 => x"93",
          9012 => x"ff",
          9013 => x"8d",
          9014 => x"a1",
          9015 => x"af",
          9016 => x"17",
          9017 => x"33",
          9018 => x"70",
          9019 => x"55",
          9020 => x"38",
          9021 => x"54",
          9022 => x"34",
          9023 => x"0b",
          9024 => x"8b",
          9025 => x"84",
          9026 => x"06",
          9027 => x"73",
          9028 => x"e7",
          9029 => x"2e",
          9030 => x"75",
          9031 => x"ff",
          9032 => x"82",
          9033 => x"52",
          9034 => x"a5",
          9035 => x"55",
          9036 => x"08",
          9037 => x"de",
          9038 => x"98",
          9039 => x"51",
          9040 => x"3f",
          9041 => x"08",
          9042 => x"11",
          9043 => x"82",
          9044 => x"80",
          9045 => x"16",
          9046 => x"ae",
          9047 => x"06",
          9048 => x"53",
          9049 => x"51",
          9050 => x"3f",
          9051 => x"0b",
          9052 => x"87",
          9053 => x"98",
          9054 => x"77",
          9055 => x"3f",
          9056 => x"08",
          9057 => x"98",
          9058 => x"78",
          9059 => x"98",
          9060 => x"98",
          9061 => x"82",
          9062 => x"aa",
          9063 => x"ec",
          9064 => x"80",
          9065 => x"02",
          9066 => x"e3",
          9067 => x"57",
          9068 => x"3d",
          9069 => x"97",
          9070 => x"c3",
          9071 => x"98",
          9072 => x"e0",
          9073 => x"cf",
          9074 => x"66",
          9075 => x"d0",
          9076 => x"c5",
          9077 => x"98",
          9078 => x"e0",
          9079 => x"38",
          9080 => x"05",
          9081 => x"06",
          9082 => x"73",
          9083 => x"a7",
          9084 => x"09",
          9085 => x"71",
          9086 => x"06",
          9087 => x"55",
          9088 => x"15",
          9089 => x"81",
          9090 => x"34",
          9091 => x"a2",
          9092 => x"e0",
          9093 => x"74",
          9094 => x"0c",
          9095 => x"04",
          9096 => x"65",
          9097 => x"94",
          9098 => x"52",
          9099 => x"d0",
          9100 => x"e0",
          9101 => x"82",
          9102 => x"80",
          9103 => x"58",
          9104 => x"3d",
          9105 => x"c4",
          9106 => x"e0",
          9107 => x"82",
          9108 => x"b4",
          9109 => x"c7",
          9110 => x"a0",
          9111 => x"55",
          9112 => x"84",
          9113 => x"17",
          9114 => x"2b",
          9115 => x"96",
          9116 => x"9d",
          9117 => x"54",
          9118 => x"15",
          9119 => x"ff",
          9120 => x"82",
          9121 => x"55",
          9122 => x"98",
          9123 => x"0d",
          9124 => x"0d",
          9125 => x"5a",
          9126 => x"3d",
          9127 => x"9a",
          9128 => x"db",
          9129 => x"98",
          9130 => x"98",
          9131 => x"82",
          9132 => x"07",
          9133 => x"55",
          9134 => x"2e",
          9135 => x"81",
          9136 => x"55",
          9137 => x"2e",
          9138 => x"7b",
          9139 => x"80",
          9140 => x"70",
          9141 => x"ac",
          9142 => x"e0",
          9143 => x"82",
          9144 => x"80",
          9145 => x"52",
          9146 => x"b1",
          9147 => x"e0",
          9148 => x"82",
          9149 => x"bf",
          9150 => x"98",
          9151 => x"98",
          9152 => x"59",
          9153 => x"81",
          9154 => x"56",
          9155 => x"33",
          9156 => x"16",
          9157 => x"27",
          9158 => x"56",
          9159 => x"80",
          9160 => x"80",
          9161 => x"ff",
          9162 => x"70",
          9163 => x"56",
          9164 => x"e8",
          9165 => x"76",
          9166 => x"81",
          9167 => x"80",
          9168 => x"57",
          9169 => x"78",
          9170 => x"51",
          9171 => x"2e",
          9172 => x"73",
          9173 => x"38",
          9174 => x"08",
          9175 => x"9f",
          9176 => x"e0",
          9177 => x"82",
          9178 => x"a7",
          9179 => x"33",
          9180 => x"c3",
          9181 => x"2e",
          9182 => x"e4",
          9183 => x"2e",
          9184 => x"56",
          9185 => x"05",
          9186 => x"92",
          9187 => x"98",
          9188 => x"76",
          9189 => x"0c",
          9190 => x"04",
          9191 => x"82",
          9192 => x"ff",
          9193 => x"9d",
          9194 => x"d3",
          9195 => x"98",
          9196 => x"98",
          9197 => x"82",
          9198 => x"82",
          9199 => x"53",
          9200 => x"3d",
          9201 => x"ff",
          9202 => x"73",
          9203 => x"51",
          9204 => x"74",
          9205 => x"38",
          9206 => x"3d",
          9207 => x"cc",
          9208 => x"98",
          9209 => x"ff",
          9210 => x"38",
          9211 => x"08",
          9212 => x"3f",
          9213 => x"82",
          9214 => x"51",
          9215 => x"82",
          9216 => x"83",
          9217 => x"55",
          9218 => x"a3",
          9219 => x"82",
          9220 => x"ff",
          9221 => x"82",
          9222 => x"93",
          9223 => x"75",
          9224 => x"75",
          9225 => x"38",
          9226 => x"76",
          9227 => x"86",
          9228 => x"39",
          9229 => x"27",
          9230 => x"88",
          9231 => x"77",
          9232 => x"59",
          9233 => x"56",
          9234 => x"81",
          9235 => x"81",
          9236 => x"33",
          9237 => x"73",
          9238 => x"fe",
          9239 => x"33",
          9240 => x"73",
          9241 => x"81",
          9242 => x"80",
          9243 => x"02",
          9244 => x"75",
          9245 => x"51",
          9246 => x"2e",
          9247 => x"87",
          9248 => x"56",
          9249 => x"78",
          9250 => x"80",
          9251 => x"70",
          9252 => x"a8",
          9253 => x"e0",
          9254 => x"82",
          9255 => x"80",
          9256 => x"52",
          9257 => x"ae",
          9258 => x"e0",
          9259 => x"82",
          9260 => x"8d",
          9261 => x"c4",
          9262 => x"e5",
          9263 => x"c6",
          9264 => x"98",
          9265 => x"09",
          9266 => x"cc",
          9267 => x"75",
          9268 => x"c4",
          9269 => x"74",
          9270 => x"d8",
          9271 => x"98",
          9272 => x"e0",
          9273 => x"38",
          9274 => x"e0",
          9275 => x"66",
          9276 => x"c5",
          9277 => x"88",
          9278 => x"34",
          9279 => x"52",
          9280 => x"99",
          9281 => x"54",
          9282 => x"15",
          9283 => x"ff",
          9284 => x"82",
          9285 => x"54",
          9286 => x"82",
          9287 => x"9c",
          9288 => x"f2",
          9289 => x"62",
          9290 => x"80",
          9291 => x"93",
          9292 => x"55",
          9293 => x"5e",
          9294 => x"3f",
          9295 => x"08",
          9296 => x"98",
          9297 => x"38",
          9298 => x"58",
          9299 => x"38",
          9300 => x"97",
          9301 => x"08",
          9302 => x"38",
          9303 => x"70",
          9304 => x"81",
          9305 => x"55",
          9306 => x"87",
          9307 => x"39",
          9308 => x"90",
          9309 => x"82",
          9310 => x"8a",
          9311 => x"89",
          9312 => x"7f",
          9313 => x"56",
          9314 => x"3f",
          9315 => x"06",
          9316 => x"72",
          9317 => x"82",
          9318 => x"05",
          9319 => x"7c",
          9320 => x"55",
          9321 => x"27",
          9322 => x"16",
          9323 => x"83",
          9324 => x"76",
          9325 => x"80",
          9326 => x"79",
          9327 => x"c1",
          9328 => x"7f",
          9329 => x"14",
          9330 => x"83",
          9331 => x"82",
          9332 => x"81",
          9333 => x"38",
          9334 => x"08",
          9335 => x"95",
          9336 => x"98",
          9337 => x"81",
          9338 => x"7b",
          9339 => x"06",
          9340 => x"39",
          9341 => x"56",
          9342 => x"09",
          9343 => x"b9",
          9344 => x"80",
          9345 => x"80",
          9346 => x"78",
          9347 => x"7a",
          9348 => x"38",
          9349 => x"73",
          9350 => x"81",
          9351 => x"ff",
          9352 => x"74",
          9353 => x"ff",
          9354 => x"82",
          9355 => x"58",
          9356 => x"08",
          9357 => x"74",
          9358 => x"16",
          9359 => x"73",
          9360 => x"39",
          9361 => x"7e",
          9362 => x"0c",
          9363 => x"2e",
          9364 => x"88",
          9365 => x"8c",
          9366 => x"1a",
          9367 => x"07",
          9368 => x"1b",
          9369 => x"08",
          9370 => x"16",
          9371 => x"75",
          9372 => x"38",
          9373 => x"94",
          9374 => x"15",
          9375 => x"54",
          9376 => x"34",
          9377 => x"82",
          9378 => x"90",
          9379 => x"e8",
          9380 => x"6e",
          9381 => x"80",
          9382 => x"9e",
          9383 => x"5c",
          9384 => x"3f",
          9385 => x"0b",
          9386 => x"08",
          9387 => x"38",
          9388 => x"08",
          9389 => x"f7",
          9390 => x"08",
          9391 => x"80",
          9392 => x"80",
          9393 => x"e0",
          9394 => x"e0",
          9395 => x"82",
          9396 => x"33",
          9397 => x"12",
          9398 => x"55",
          9399 => x"51",
          9400 => x"3f",
          9401 => x"08",
          9402 => x"70",
          9403 => x"57",
          9404 => x"8c",
          9405 => x"82",
          9406 => x"06",
          9407 => x"56",
          9408 => x"38",
          9409 => x"05",
          9410 => x"7f",
          9411 => x"cc",
          9412 => x"98",
          9413 => x"68",
          9414 => x"2e",
          9415 => x"82",
          9416 => x"8b",
          9417 => x"75",
          9418 => x"80",
          9419 => x"81",
          9420 => x"2e",
          9421 => x"80",
          9422 => x"38",
          9423 => x"0a",
          9424 => x"ff",
          9425 => x"55",
          9426 => x"86",
          9427 => x"8b",
          9428 => x"89",
          9429 => x"2a",
          9430 => x"77",
          9431 => x"59",
          9432 => x"81",
          9433 => x"70",
          9434 => x"07",
          9435 => x"56",
          9436 => x"38",
          9437 => x"80",
          9438 => x"54",
          9439 => x"52",
          9440 => x"8e",
          9441 => x"56",
          9442 => x"08",
          9443 => x"83",
          9444 => x"ff",
          9445 => x"82",
          9446 => x"83",
          9447 => x"55",
          9448 => x"82",
          9449 => x"09",
          9450 => x"a3",
          9451 => x"29",
          9452 => x"11",
          9453 => x"74",
          9454 => x"93",
          9455 => x"17",
          9456 => x"da",
          9457 => x"98",
          9458 => x"18",
          9459 => x"92",
          9460 => x"e0",
          9461 => x"b7",
          9462 => x"f8",
          9463 => x"52",
          9464 => x"90",
          9465 => x"56",
          9466 => x"08",
          9467 => x"62",
          9468 => x"77",
          9469 => x"98",
          9470 => x"55",
          9471 => x"bf",
          9472 => x"8e",
          9473 => x"26",
          9474 => x"74",
          9475 => x"8e",
          9476 => x"68",
          9477 => x"38",
          9478 => x"81",
          9479 => x"af",
          9480 => x"2a",
          9481 => x"56",
          9482 => x"2e",
          9483 => x"87",
          9484 => x"82",
          9485 => x"38",
          9486 => x"55",
          9487 => x"83",
          9488 => x"81",
          9489 => x"56",
          9490 => x"80",
          9491 => x"38",
          9492 => x"83",
          9493 => x"06",
          9494 => x"78",
          9495 => x"91",
          9496 => x"0b",
          9497 => x"22",
          9498 => x"80",
          9499 => x"74",
          9500 => x"38",
          9501 => x"56",
          9502 => x"17",
          9503 => x"57",
          9504 => x"2e",
          9505 => x"75",
          9506 => x"79",
          9507 => x"fe",
          9508 => x"82",
          9509 => x"84",
          9510 => x"05",
          9511 => x"5e",
          9512 => x"80",
          9513 => x"98",
          9514 => x"8a",
          9515 => x"fd",
          9516 => x"75",
          9517 => x"38",
          9518 => x"78",
          9519 => x"8c",
          9520 => x"0b",
          9521 => x"22",
          9522 => x"80",
          9523 => x"74",
          9524 => x"38",
          9525 => x"56",
          9526 => x"17",
          9527 => x"57",
          9528 => x"2e",
          9529 => x"75",
          9530 => x"79",
          9531 => x"fe",
          9532 => x"82",
          9533 => x"10",
          9534 => x"82",
          9535 => x"9f",
          9536 => x"38",
          9537 => x"e0",
          9538 => x"82",
          9539 => x"05",
          9540 => x"2a",
          9541 => x"56",
          9542 => x"17",
          9543 => x"81",
          9544 => x"7b",
          9545 => x"67",
          9546 => x"12",
          9547 => x"30",
          9548 => x"74",
          9549 => x"59",
          9550 => x"7d",
          9551 => x"81",
          9552 => x"76",
          9553 => x"42",
          9554 => x"76",
          9555 => x"90",
          9556 => x"60",
          9557 => x"51",
          9558 => x"26",
          9559 => x"75",
          9560 => x"31",
          9561 => x"67",
          9562 => x"fe",
          9563 => x"82",
          9564 => x"58",
          9565 => x"09",
          9566 => x"38",
          9567 => x"08",
          9568 => x"26",
          9569 => x"78",
          9570 => x"79",
          9571 => x"78",
          9572 => x"87",
          9573 => x"82",
          9574 => x"06",
          9575 => x"83",
          9576 => x"82",
          9577 => x"27",
          9578 => x"8f",
          9579 => x"55",
          9580 => x"26",
          9581 => x"59",
          9582 => x"63",
          9583 => x"74",
          9584 => x"38",
          9585 => x"88",
          9586 => x"98",
          9587 => x"26",
          9588 => x"86",
          9589 => x"1a",
          9590 => x"79",
          9591 => x"38",
          9592 => x"80",
          9593 => x"2e",
          9594 => x"83",
          9595 => x"9f",
          9596 => x"8b",
          9597 => x"06",
          9598 => x"74",
          9599 => x"84",
          9600 => x"52",
          9601 => x"8f",
          9602 => x"53",
          9603 => x"52",
          9604 => x"8f",
          9605 => x"80",
          9606 => x"51",
          9607 => x"3f",
          9608 => x"34",
          9609 => x"ff",
          9610 => x"1b",
          9611 => x"99",
          9612 => x"90",
          9613 => x"83",
          9614 => x"70",
          9615 => x"80",
          9616 => x"55",
          9617 => x"ff",
          9618 => x"67",
          9619 => x"ff",
          9620 => x"38",
          9621 => x"ff",
          9622 => x"1b",
          9623 => x"e9",
          9624 => x"74",
          9625 => x"51",
          9626 => x"3f",
          9627 => x"1c",
          9628 => x"98",
          9629 => x"8d",
          9630 => x"ff",
          9631 => x"51",
          9632 => x"3f",
          9633 => x"1b",
          9634 => x"db",
          9635 => x"2e",
          9636 => x"80",
          9637 => x"88",
          9638 => x"80",
          9639 => x"ff",
          9640 => x"7c",
          9641 => x"51",
          9642 => x"3f",
          9643 => x"1b",
          9644 => x"b3",
          9645 => x"b0",
          9646 => x"8d",
          9647 => x"52",
          9648 => x"ff",
          9649 => x"ff",
          9650 => x"c0",
          9651 => x"0b",
          9652 => x"34",
          9653 => x"d1",
          9654 => x"c7",
          9655 => x"39",
          9656 => x"0a",
          9657 => x"51",
          9658 => x"3f",
          9659 => x"ff",
          9660 => x"1b",
          9661 => x"d1",
          9662 => x"0b",
          9663 => x"a9",
          9664 => x"34",
          9665 => x"d2",
          9666 => x"1b",
          9667 => x"86",
          9668 => x"d5",
          9669 => x"1b",
          9670 => x"ff",
          9671 => x"81",
          9672 => x"7a",
          9673 => x"ff",
          9674 => x"81",
          9675 => x"98",
          9676 => x"38",
          9677 => x"09",
          9678 => x"ec",
          9679 => x"86",
          9680 => x"52",
          9681 => x"88",
          9682 => x"80",
          9683 => x"7a",
          9684 => x"e5",
          9685 => x"85",
          9686 => x"7a",
          9687 => x"87",
          9688 => x"85",
          9689 => x"83",
          9690 => x"ff",
          9691 => x"ff",
          9692 => x"e8",
          9693 => x"8b",
          9694 => x"52",
          9695 => x"51",
          9696 => x"3f",
          9697 => x"52",
          9698 => x"8b",
          9699 => x"54",
          9700 => x"7a",
          9701 => x"ff",
          9702 => x"75",
          9703 => x"53",
          9704 => x"51",
          9705 => x"3f",
          9706 => x"52",
          9707 => x"8c",
          9708 => x"56",
          9709 => x"83",
          9710 => x"06",
          9711 => x"52",
          9712 => x"8b",
          9713 => x"52",
          9714 => x"ff",
          9715 => x"f0",
          9716 => x"1b",
          9717 => x"87",
          9718 => x"55",
          9719 => x"83",
          9720 => x"74",
          9721 => x"ff",
          9722 => x"7c",
          9723 => x"74",
          9724 => x"38",
          9725 => x"54",
          9726 => x"52",
          9727 => x"86",
          9728 => x"e0",
          9729 => x"be",
          9730 => x"53",
          9731 => x"08",
          9732 => x"ff",
          9733 => x"76",
          9734 => x"31",
          9735 => x"cd",
          9736 => x"58",
          9737 => x"ff",
          9738 => x"55",
          9739 => x"83",
          9740 => x"61",
          9741 => x"26",
          9742 => x"57",
          9743 => x"53",
          9744 => x"51",
          9745 => x"3f",
          9746 => x"08",
          9747 => x"76",
          9748 => x"31",
          9749 => x"db",
          9750 => x"7d",
          9751 => x"38",
          9752 => x"83",
          9753 => x"8a",
          9754 => x"7d",
          9755 => x"38",
          9756 => x"80",
          9757 => x"81",
          9758 => x"7a",
          9759 => x"ff",
          9760 => x"81",
          9761 => x"98",
          9762 => x"38",
          9763 => x"1b",
          9764 => x"b2",
          9765 => x"54",
          9766 => x"08",
          9767 => x"7f",
          9768 => x"d4",
          9769 => x"39",
          9770 => x"81",
          9771 => x"80",
          9772 => x"80",
          9773 => x"7a",
          9774 => x"fd",
          9775 => x"d5",
          9776 => x"ff",
          9777 => x"83",
          9778 => x"77",
          9779 => x"0b",
          9780 => x"81",
          9781 => x"34",
          9782 => x"34",
          9783 => x"34",
          9784 => x"80",
          9785 => x"75",
          9786 => x"ea",
          9787 => x"85",
          9788 => x"e0",
          9789 => x"2a",
          9790 => x"75",
          9791 => x"82",
          9792 => x"87",
          9793 => x"52",
          9794 => x"51",
          9795 => x"3f",
          9796 => x"ca",
          9797 => x"88",
          9798 => x"54",
          9799 => x"52",
          9800 => x"84",
          9801 => x"56",
          9802 => x"08",
          9803 => x"53",
          9804 => x"51",
          9805 => x"3f",
          9806 => x"e0",
          9807 => x"38",
          9808 => x"56",
          9809 => x"56",
          9810 => x"e0",
          9811 => x"75",
          9812 => x"0c",
          9813 => x"04",
          9814 => x"7d",
          9815 => x"80",
          9816 => x"05",
          9817 => x"76",
          9818 => x"38",
          9819 => x"11",
          9820 => x"53",
          9821 => x"79",
          9822 => x"3f",
          9823 => x"09",
          9824 => x"38",
          9825 => x"55",
          9826 => x"db",
          9827 => x"70",
          9828 => x"34",
          9829 => x"74",
          9830 => x"81",
          9831 => x"80",
          9832 => x"55",
          9833 => x"76",
          9834 => x"e0",
          9835 => x"3d",
          9836 => x"3d",
          9837 => x"84",
          9838 => x"33",
          9839 => x"8a",
          9840 => x"06",
          9841 => x"52",
          9842 => x"3f",
          9843 => x"56",
          9844 => x"be",
          9845 => x"08",
          9846 => x"05",
          9847 => x"75",
          9848 => x"56",
          9849 => x"a1",
          9850 => x"fc",
          9851 => x"53",
          9852 => x"76",
          9853 => x"97",
          9854 => x"32",
          9855 => x"72",
          9856 => x"70",
          9857 => x"56",
          9858 => x"18",
          9859 => x"88",
          9860 => x"3d",
          9861 => x"3d",
          9862 => x"11",
          9863 => x"80",
          9864 => x"38",
          9865 => x"05",
          9866 => x"8c",
          9867 => x"08",
          9868 => x"3f",
          9869 => x"08",
          9870 => x"16",
          9871 => x"09",
          9872 => x"38",
          9873 => x"55",
          9874 => x"55",
          9875 => x"98",
          9876 => x"0d",
          9877 => x"0d",
          9878 => x"cc",
          9879 => x"73",
          9880 => x"d5",
          9881 => x"0c",
          9882 => x"04",
          9883 => x"02",
          9884 => x"33",
          9885 => x"3d",
          9886 => x"54",
          9887 => x"52",
          9888 => x"ae",
          9889 => x"ff",
          9890 => x"3d",
          9891 => x"3d",
          9892 => x"84",
          9893 => x"22",
          9894 => x"52",
          9895 => x"26",
          9896 => x"83",
          9897 => x"52",
          9898 => x"83",
          9899 => x"27",
          9900 => x"b5",
          9901 => x"06",
          9902 => x"80",
          9903 => x"82",
          9904 => x"51",
          9905 => x"9c",
          9906 => x"70",
          9907 => x"06",
          9908 => x"80",
          9909 => x"38",
          9910 => x"d3",
          9911 => x"22",
          9912 => x"39",
          9913 => x"70",
          9914 => x"53",
          9915 => x"e0",
          9916 => x"3d",
          9917 => x"3d",
          9918 => x"05",
          9919 => x"05",
          9920 => x"53",
          9921 => x"70",
          9922 => x"85",
          9923 => x"9a",
          9924 => x"b5",
          9925 => x"06",
          9926 => x"81",
          9927 => x"38",
          9928 => x"d1",
          9929 => x"22",
          9930 => x"82",
          9931 => x"84",
          9932 => x"fb",
          9933 => x"51",
          9934 => x"ff",
          9935 => x"38",
          9936 => x"ff",
          9937 => x"ec",
          9938 => x"ff",
          9939 => x"38",
          9940 => x"56",
          9941 => x"05",
          9942 => x"30",
          9943 => x"72",
          9944 => x"51",
          9945 => x"80",
          9946 => x"70",
          9947 => x"22",
          9948 => x"71",
          9949 => x"70",
          9950 => x"55",
          9951 => x"25",
          9952 => x"73",
          9953 => x"dc",
          9954 => x"29",
          9955 => x"05",
          9956 => x"04",
          9957 => x"10",
          9958 => x"22",
          9959 => x"80",
          9960 => x"75",
          9961 => x"72",
          9962 => x"51",
          9963 => x"12",
          9964 => x"e0",
          9965 => x"39",
          9966 => x"95",
          9967 => x"51",
          9968 => x"12",
          9969 => x"ff",
          9970 => x"85",
          9971 => x"12",
          9972 => x"ff",
          9973 => x"8c",
          9974 => x"f8",
          9975 => x"16",
          9976 => x"39",
          9977 => x"82",
          9978 => x"87",
          9979 => x"00",
          9980 => x"ff",
          9981 => x"ff",
          9982 => x"ff",
          9983 => x"00",
          9984 => x"00",
          9985 => x"00",
          9986 => x"00",
          9987 => x"00",
          9988 => x"00",
          9989 => x"00",
          9990 => x"00",
          9991 => x"00",
          9992 => x"00",
          9993 => x"00",
          9994 => x"00",
          9995 => x"00",
          9996 => x"00",
          9997 => x"00",
          9998 => x"00",
          9999 => x"00",
         10000 => x"00",
         10001 => x"00",
         10002 => x"00",
         10003 => x"00",
         10004 => x"00",
         10005 => x"00",
         10006 => x"00",
         10007 => x"00",
         10008 => x"00",
         10009 => x"00",
         10010 => x"00",
         10011 => x"00",
         10012 => x"00",
         10013 => x"00",
         10014 => x"00",
         10015 => x"00",
         10016 => x"00",
         10017 => x"00",
         10018 => x"00",
         10019 => x"00",
         10020 => x"00",
         10021 => x"00",
         10022 => x"00",
         10023 => x"00",
         10024 => x"00",
         10025 => x"00",
         10026 => x"00",
         10027 => x"00",
         10028 => x"00",
         10029 => x"00",
         10030 => x"00",
         10031 => x"00",
         10032 => x"00",
         10033 => x"00",
         10034 => x"00",
         10035 => x"00",
         10036 => x"00",
         10037 => x"00",
         10038 => x"00",
         10039 => x"00",
         10040 => x"00",
         10041 => x"00",
         10042 => x"00",
         10043 => x"00",
         10044 => x"00",
         10045 => x"00",
         10046 => x"00",
         10047 => x"00",
         10048 => x"00",
         10049 => x"00",
         10050 => x"00",
         10051 => x"00",
         10052 => x"00",
         10053 => x"00",
         10054 => x"00",
         10055 => x"00",
         10056 => x"00",
         10057 => x"00",
         10058 => x"00",
         10059 => x"00",
         10060 => x"00",
         10061 => x"00",
         10062 => x"00",
         10063 => x"00",
         10064 => x"00",
         10065 => x"00",
         10066 => x"00",
         10067 => x"00",
         10068 => x"00",
         10069 => x"00",
         10070 => x"00",
         10071 => x"00",
         10072 => x"00",
         10073 => x"00",
         10074 => x"00",
         10075 => x"00",
         10076 => x"00",
         10077 => x"00",
         10078 => x"00",
         10079 => x"00",
         10080 => x"00",
         10081 => x"00",
         10082 => x"00",
         10083 => x"00",
         10084 => x"00",
         10085 => x"00",
         10086 => x"00",
         10087 => x"00",
         10088 => x"00",
         10089 => x"00",
         10090 => x"00",
         10091 => x"00",
         10092 => x"00",
         10093 => x"00",
         10094 => x"00",
         10095 => x"00",
         10096 => x"00",
         10097 => x"00",
         10098 => x"00",
         10099 => x"00",
         10100 => x"00",
         10101 => x"00",
         10102 => x"00",
         10103 => x"00",
         10104 => x"00",
         10105 => x"00",
         10106 => x"00",
         10107 => x"00",
         10108 => x"00",
         10109 => x"00",
         10110 => x"00",
         10111 => x"00",
         10112 => x"00",
         10113 => x"00",
         10114 => x"00",
         10115 => x"00",
         10116 => x"00",
         10117 => x"00",
         10118 => x"00",
         10119 => x"00",
         10120 => x"00",
         10121 => x"00",
         10122 => x"00",
         10123 => x"00",
         10124 => x"00",
         10125 => x"00",
         10126 => x"00",
         10127 => x"00",
         10128 => x"64",
         10129 => x"74",
         10130 => x"64",
         10131 => x"74",
         10132 => x"66",
         10133 => x"74",
         10134 => x"66",
         10135 => x"64",
         10136 => x"66",
         10137 => x"63",
         10138 => x"6d",
         10139 => x"61",
         10140 => x"6d",
         10141 => x"79",
         10142 => x"6d",
         10143 => x"66",
         10144 => x"6d",
         10145 => x"70",
         10146 => x"6d",
         10147 => x"6d",
         10148 => x"6d",
         10149 => x"68",
         10150 => x"68",
         10151 => x"68",
         10152 => x"68",
         10153 => x"63",
         10154 => x"00",
         10155 => x"6a",
         10156 => x"72",
         10157 => x"61",
         10158 => x"72",
         10159 => x"74",
         10160 => x"69",
         10161 => x"00",
         10162 => x"74",
         10163 => x"69",
         10164 => x"6d",
         10165 => x"69",
         10166 => x"6b",
         10167 => x"00",
         10168 => x"65",
         10169 => x"44",
         10170 => x"20",
         10171 => x"6f",
         10172 => x"49",
         10173 => x"72",
         10174 => x"20",
         10175 => x"6f",
         10176 => x"44",
         10177 => x"20",
         10178 => x"20",
         10179 => x"64",
         10180 => x"4e",
         10181 => x"69",
         10182 => x"66",
         10183 => x"64",
         10184 => x"4e",
         10185 => x"61",
         10186 => x"66",
         10187 => x"64",
         10188 => x"49",
         10189 => x"6c",
         10190 => x"66",
         10191 => x"6e",
         10192 => x"2e",
         10193 => x"41",
         10194 => x"73",
         10195 => x"65",
         10196 => x"64",
         10197 => x"46",
         10198 => x"20",
         10199 => x"65",
         10200 => x"20",
         10201 => x"73",
         10202 => x"00",
         10203 => x"46",
         10204 => x"20",
         10205 => x"64",
         10206 => x"69",
         10207 => x"6c",
         10208 => x"00",
         10209 => x"53",
         10210 => x"73",
         10211 => x"69",
         10212 => x"70",
         10213 => x"65",
         10214 => x"64",
         10215 => x"44",
         10216 => x"65",
         10217 => x"6d",
         10218 => x"20",
         10219 => x"69",
         10220 => x"6c",
         10221 => x"00",
         10222 => x"44",
         10223 => x"20",
         10224 => x"20",
         10225 => x"62",
         10226 => x"2e",
         10227 => x"4e",
         10228 => x"6f",
         10229 => x"74",
         10230 => x"65",
         10231 => x"6c",
         10232 => x"73",
         10233 => x"20",
         10234 => x"6e",
         10235 => x"6e",
         10236 => x"73",
         10237 => x"46",
         10238 => x"61",
         10239 => x"62",
         10240 => x"65",
         10241 => x"54",
         10242 => x"6f",
         10243 => x"20",
         10244 => x"72",
         10245 => x"6f",
         10246 => x"61",
         10247 => x"6c",
         10248 => x"2e",
         10249 => x"46",
         10250 => x"20",
         10251 => x"6c",
         10252 => x"65",
         10253 => x"49",
         10254 => x"66",
         10255 => x"69",
         10256 => x"20",
         10257 => x"6f",
         10258 => x"00",
         10259 => x"54",
         10260 => x"6d",
         10261 => x"20",
         10262 => x"6e",
         10263 => x"6c",
         10264 => x"00",
         10265 => x"50",
         10266 => x"6d",
         10267 => x"72",
         10268 => x"6e",
         10269 => x"72",
         10270 => x"2e",
         10271 => x"53",
         10272 => x"65",
         10273 => x"00",
         10274 => x"55",
         10275 => x"6f",
         10276 => x"65",
         10277 => x"72",
         10278 => x"0a",
         10279 => x"20",
         10280 => x"65",
         10281 => x"73",
         10282 => x"20",
         10283 => x"20",
         10284 => x"65",
         10285 => x"65",
         10286 => x"00",
         10287 => x"72",
         10288 => x"00",
         10289 => x"25",
         10290 => x"58",
         10291 => x"3a",
         10292 => x"25",
         10293 => x"00",
         10294 => x"20",
         10295 => x"20",
         10296 => x"00",
         10297 => x"25",
         10298 => x"00",
         10299 => x"20",
         10300 => x"20",
         10301 => x"7c",
         10302 => x"7a",
         10303 => x"2a",
         10304 => x"73",
         10305 => x"31",
         10306 => x"32",
         10307 => x"32",
         10308 => x"76",
         10309 => x"63",
         10310 => x"20",
         10311 => x"2c",
         10312 => x"76",
         10313 => x"32",
         10314 => x"25",
         10315 => x"73",
         10316 => x"0a",
         10317 => x"5a",
         10318 => x"49",
         10319 => x"72",
         10320 => x"74",
         10321 => x"6e",
         10322 => x"72",
         10323 => x"54",
         10324 => x"72",
         10325 => x"74",
         10326 => x"75",
         10327 => x"50",
         10328 => x"69",
         10329 => x"72",
         10330 => x"74",
         10331 => x"49",
         10332 => x"4c",
         10333 => x"20",
         10334 => x"65",
         10335 => x"70",
         10336 => x"49",
         10337 => x"4c",
         10338 => x"20",
         10339 => x"65",
         10340 => x"70",
         10341 => x"55",
         10342 => x"30",
         10343 => x"20",
         10344 => x"65",
         10345 => x"70",
         10346 => x"55",
         10347 => x"30",
         10348 => x"20",
         10349 => x"65",
         10350 => x"70",
         10351 => x"55",
         10352 => x"31",
         10353 => x"20",
         10354 => x"65",
         10355 => x"70",
         10356 => x"55",
         10357 => x"31",
         10358 => x"20",
         10359 => x"65",
         10360 => x"70",
         10361 => x"53",
         10362 => x"69",
         10363 => x"75",
         10364 => x"69",
         10365 => x"2e",
         10366 => x"45",
         10367 => x"6c",
         10368 => x"20",
         10369 => x"65",
         10370 => x"2e",
         10371 => x"61",
         10372 => x"65",
         10373 => x"2e",
         10374 => x"00",
         10375 => x"7a",
         10376 => x"7a",
         10377 => x"68",
         10378 => x"30",
         10379 => x"46",
         10380 => x"65",
         10381 => x"6f",
         10382 => x"69",
         10383 => x"6c",
         10384 => x"20",
         10385 => x"63",
         10386 => x"20",
         10387 => x"70",
         10388 => x"73",
         10389 => x"6e",
         10390 => x"6d",
         10391 => x"61",
         10392 => x"2e",
         10393 => x"2a",
         10394 => x"43",
         10395 => x"72",
         10396 => x"2e",
         10397 => x"00",
         10398 => x"43",
         10399 => x"69",
         10400 => x"2e",
         10401 => x"43",
         10402 => x"61",
         10403 => x"67",
         10404 => x"00",
         10405 => x"25",
         10406 => x"78",
         10407 => x"38",
         10408 => x"3e",
         10409 => x"6c",
         10410 => x"30",
         10411 => x"0a",
         10412 => x"44",
         10413 => x"20",
         10414 => x"6f",
         10415 => x"0a",
         10416 => x"70",
         10417 => x"65",
         10418 => x"25",
         10419 => x"58",
         10420 => x"32",
         10421 => x"3f",
         10422 => x"25",
         10423 => x"58",
         10424 => x"34",
         10425 => x"25",
         10426 => x"58",
         10427 => x"38",
         10428 => x"00",
         10429 => x"45",
         10430 => x"75",
         10431 => x"67",
         10432 => x"64",
         10433 => x"20",
         10434 => x"6c",
         10435 => x"2e",
         10436 => x"43",
         10437 => x"69",
         10438 => x"63",
         10439 => x"20",
         10440 => x"30",
         10441 => x"20",
         10442 => x"0a",
         10443 => x"43",
         10444 => x"20",
         10445 => x"75",
         10446 => x"64",
         10447 => x"64",
         10448 => x"25",
         10449 => x"0a",
         10450 => x"52",
         10451 => x"61",
         10452 => x"6e",
         10453 => x"70",
         10454 => x"63",
         10455 => x"6f",
         10456 => x"2e",
         10457 => x"43",
         10458 => x"20",
         10459 => x"6f",
         10460 => x"6e",
         10461 => x"2e",
         10462 => x"5a",
         10463 => x"62",
         10464 => x"25",
         10465 => x"25",
         10466 => x"73",
         10467 => x"00",
         10468 => x"25",
         10469 => x"25",
         10470 => x"73",
         10471 => x"25",
         10472 => x"25",
         10473 => x"42",
         10474 => x"63",
         10475 => x"61",
         10476 => x"00",
         10477 => x"4d",
         10478 => x"72",
         10479 => x"78",
         10480 => x"73",
         10481 => x"2c",
         10482 => x"6e",
         10483 => x"20",
         10484 => x"63",
         10485 => x"20",
         10486 => x"6d",
         10487 => x"2e",
         10488 => x"52",
         10489 => x"69",
         10490 => x"2e",
         10491 => x"45",
         10492 => x"6c",
         10493 => x"20",
         10494 => x"65",
         10495 => x"70",
         10496 => x"2e",
         10497 => x"25",
         10498 => x"64",
         10499 => x"20",
         10500 => x"25",
         10501 => x"64",
         10502 => x"25",
         10503 => x"53",
         10504 => x"43",
         10505 => x"69",
         10506 => x"61",
         10507 => x"6e",
         10508 => x"20",
         10509 => x"6f",
         10510 => x"6f",
         10511 => x"6f",
         10512 => x"67",
         10513 => x"3a",
         10514 => x"76",
         10515 => x"73",
         10516 => x"70",
         10517 => x"65",
         10518 => x"64",
         10519 => x"20",
         10520 => x"57",
         10521 => x"44",
         10522 => x"20",
         10523 => x"30",
         10524 => x"25",
         10525 => x"29",
         10526 => x"20",
         10527 => x"53",
         10528 => x"4d",
         10529 => x"20",
         10530 => x"30",
         10531 => x"25",
         10532 => x"29",
         10533 => x"20",
         10534 => x"49",
         10535 => x"20",
         10536 => x"4d",
         10537 => x"30",
         10538 => x"25",
         10539 => x"29",
         10540 => x"20",
         10541 => x"42",
         10542 => x"20",
         10543 => x"20",
         10544 => x"30",
         10545 => x"25",
         10546 => x"29",
         10547 => x"20",
         10548 => x"52",
         10549 => x"20",
         10550 => x"20",
         10551 => x"30",
         10552 => x"25",
         10553 => x"29",
         10554 => x"20",
         10555 => x"53",
         10556 => x"41",
         10557 => x"20",
         10558 => x"65",
         10559 => x"65",
         10560 => x"25",
         10561 => x"29",
         10562 => x"20",
         10563 => x"54",
         10564 => x"52",
         10565 => x"20",
         10566 => x"69",
         10567 => x"73",
         10568 => x"25",
         10569 => x"29",
         10570 => x"20",
         10571 => x"49",
         10572 => x"20",
         10573 => x"4c",
         10574 => x"68",
         10575 => x"65",
         10576 => x"25",
         10577 => x"29",
         10578 => x"20",
         10579 => x"57",
         10580 => x"42",
         10581 => x"20",
         10582 => x"00",
         10583 => x"20",
         10584 => x"57",
         10585 => x"32",
         10586 => x"20",
         10587 => x"49",
         10588 => x"4c",
         10589 => x"20",
         10590 => x"50",
         10591 => x"20",
         10592 => x"53",
         10593 => x"41",
         10594 => x"65",
         10595 => x"73",
         10596 => x"20",
         10597 => x"43",
         10598 => x"52",
         10599 => x"74",
         10600 => x"63",
         10601 => x"20",
         10602 => x"72",
         10603 => x"20",
         10604 => x"30",
         10605 => x"00",
         10606 => x"20",
         10607 => x"43",
         10608 => x"4d",
         10609 => x"72",
         10610 => x"74",
         10611 => x"20",
         10612 => x"72",
         10613 => x"20",
         10614 => x"30",
         10615 => x"00",
         10616 => x"20",
         10617 => x"53",
         10618 => x"6b",
         10619 => x"61",
         10620 => x"41",
         10621 => x"65",
         10622 => x"20",
         10623 => x"20",
         10624 => x"30",
         10625 => x"00",
         10626 => x"4d",
         10627 => x"3a",
         10628 => x"20",
         10629 => x"5a",
         10630 => x"49",
         10631 => x"20",
         10632 => x"20",
         10633 => x"20",
         10634 => x"20",
         10635 => x"20",
         10636 => x"30",
         10637 => x"00",
         10638 => x"20",
         10639 => x"53",
         10640 => x"65",
         10641 => x"6c",
         10642 => x"20",
         10643 => x"71",
         10644 => x"20",
         10645 => x"20",
         10646 => x"64",
         10647 => x"34",
         10648 => x"7a",
         10649 => x"20",
         10650 => x"53",
         10651 => x"4d",
         10652 => x"6f",
         10653 => x"46",
         10654 => x"20",
         10655 => x"20",
         10656 => x"20",
         10657 => x"64",
         10658 => x"34",
         10659 => x"7a",
         10660 => x"20",
         10661 => x"57",
         10662 => x"62",
         10663 => x"20",
         10664 => x"41",
         10665 => x"6c",
         10666 => x"20",
         10667 => x"71",
         10668 => x"64",
         10669 => x"34",
         10670 => x"7a",
         10671 => x"53",
         10672 => x"6c",
         10673 => x"4d",
         10674 => x"75",
         10675 => x"46",
         10676 => x"00",
         10677 => x"45",
         10678 => x"45",
         10679 => x"00",
         10680 => x"55",
         10681 => x"6f",
         10682 => x"00",
         10683 => x"01",
         10684 => x"00",
         10685 => x"00",
         10686 => x"01",
         10687 => x"00",
         10688 => x"00",
         10689 => x"01",
         10690 => x"00",
         10691 => x"00",
         10692 => x"01",
         10693 => x"00",
         10694 => x"00",
         10695 => x"01",
         10696 => x"00",
         10697 => x"00",
         10698 => x"01",
         10699 => x"00",
         10700 => x"00",
         10701 => x"01",
         10702 => x"00",
         10703 => x"00",
         10704 => x"01",
         10705 => x"00",
         10706 => x"00",
         10707 => x"01",
         10708 => x"00",
         10709 => x"00",
         10710 => x"01",
         10711 => x"00",
         10712 => x"00",
         10713 => x"01",
         10714 => x"00",
         10715 => x"00",
         10716 => x"04",
         10717 => x"00",
         10718 => x"00",
         10719 => x"04",
         10720 => x"00",
         10721 => x"00",
         10722 => x"04",
         10723 => x"00",
         10724 => x"00",
         10725 => x"03",
         10726 => x"00",
         10727 => x"00",
         10728 => x"04",
         10729 => x"00",
         10730 => x"00",
         10731 => x"04",
         10732 => x"00",
         10733 => x"00",
         10734 => x"04",
         10735 => x"00",
         10736 => x"00",
         10737 => x"03",
         10738 => x"00",
         10739 => x"00",
         10740 => x"03",
         10741 => x"00",
         10742 => x"00",
         10743 => x"03",
         10744 => x"00",
         10745 => x"00",
         10746 => x"03",
         10747 => x"00",
         10748 => x"1b",
         10749 => x"1b",
         10750 => x"1b",
         10751 => x"1b",
         10752 => x"1b",
         10753 => x"1b",
         10754 => x"1b",
         10755 => x"1b",
         10756 => x"1b",
         10757 => x"1b",
         10758 => x"1b",
         10759 => x"10",
         10760 => x"0e",
         10761 => x"0d",
         10762 => x"0b",
         10763 => x"08",
         10764 => x"06",
         10765 => x"05",
         10766 => x"04",
         10767 => x"03",
         10768 => x"02",
         10769 => x"01",
         10770 => x"68",
         10771 => x"6f",
         10772 => x"68",
         10773 => x"00",
         10774 => x"21",
         10775 => x"25",
         10776 => x"75",
         10777 => x"73",
         10778 => x"46",
         10779 => x"65",
         10780 => x"6f",
         10781 => x"73",
         10782 => x"74",
         10783 => x"68",
         10784 => x"6f",
         10785 => x"66",
         10786 => x"20",
         10787 => x"45",
         10788 => x"00",
         10789 => x"43",
         10790 => x"6f",
         10791 => x"70",
         10792 => x"63",
         10793 => x"74",
         10794 => x"69",
         10795 => x"72",
         10796 => x"69",
         10797 => x"20",
         10798 => x"61",
         10799 => x"6e",
         10800 => x"53",
         10801 => x"22",
         10802 => x"3e",
         10803 => x"00",
         10804 => x"2b",
         10805 => x"5b",
         10806 => x"46",
         10807 => x"46",
         10808 => x"32",
         10809 => x"eb",
         10810 => x"53",
         10811 => x"35",
         10812 => x"4e",
         10813 => x"41",
         10814 => x"20",
         10815 => x"41",
         10816 => x"20",
         10817 => x"4e",
         10818 => x"41",
         10819 => x"20",
         10820 => x"41",
         10821 => x"20",
         10822 => x"00",
         10823 => x"00",
         10824 => x"00",
         10825 => x"00",
         10826 => x"01",
         10827 => x"09",
         10828 => x"14",
         10829 => x"1e",
         10830 => x"80",
         10831 => x"8e",
         10832 => x"45",
         10833 => x"49",
         10834 => x"90",
         10835 => x"99",
         10836 => x"59",
         10837 => x"9c",
         10838 => x"41",
         10839 => x"a5",
         10840 => x"a8",
         10841 => x"ac",
         10842 => x"b0",
         10843 => x"b4",
         10844 => x"b8",
         10845 => x"bc",
         10846 => x"c0",
         10847 => x"c4",
         10848 => x"c8",
         10849 => x"cc",
         10850 => x"d0",
         10851 => x"d4",
         10852 => x"d8",
         10853 => x"dc",
         10854 => x"e0",
         10855 => x"e4",
         10856 => x"e8",
         10857 => x"ec",
         10858 => x"f0",
         10859 => x"f4",
         10860 => x"f8",
         10861 => x"fc",
         10862 => x"2b",
         10863 => x"3d",
         10864 => x"5c",
         10865 => x"3c",
         10866 => x"7f",
         10867 => x"00",
         10868 => x"00",
         10869 => x"01",
         10870 => x"00",
         10871 => x"00",
         10872 => x"00",
         10873 => x"00",
         10874 => x"00",
         10875 => x"00",
         10876 => x"00",
         10877 => x"00",
         10878 => x"00",
         10879 => x"00",
         10880 => x"00",
         10881 => x"00",
         10882 => x"00",
         10883 => x"00",
         10884 => x"00",
         10885 => x"00",
         10886 => x"00",
         10887 => x"00",
         10888 => x"00",
         10889 => x"00",
         10890 => x"20",
         10891 => x"00",
         10892 => x"00",
         10893 => x"00",
         10894 => x"00",
         10895 => x"00",
         10896 => x"00",
         10897 => x"00",
         10898 => x"00",
         10899 => x"25",
         10900 => x"25",
         10901 => x"25",
         10902 => x"25",
         10903 => x"25",
         10904 => x"25",
         10905 => x"25",
         10906 => x"25",
         10907 => x"25",
         10908 => x"25",
         10909 => x"25",
         10910 => x"25",
         10911 => x"25",
         10912 => x"25",
         10913 => x"25",
         10914 => x"25",
         10915 => x"25",
         10916 => x"25",
         10917 => x"25",
         10918 => x"25",
         10919 => x"25",
         10920 => x"25",
         10921 => x"25",
         10922 => x"25",
         10923 => x"03",
         10924 => x"03",
         10925 => x"03",
         10926 => x"00",
         10927 => x"03",
         10928 => x"03",
         10929 => x"22",
         10930 => x"03",
         10931 => x"22",
         10932 => x"22",
         10933 => x"23",
         10934 => x"00",
         10935 => x"00",
         10936 => x"00",
         10937 => x"20",
         10938 => x"25",
         10939 => x"00",
         10940 => x"00",
         10941 => x"00",
         10942 => x"00",
         10943 => x"01",
         10944 => x"01",
         10945 => x"01",
         10946 => x"01",
         10947 => x"01",
         10948 => x"01",
         10949 => x"00",
         10950 => x"01",
         10951 => x"01",
         10952 => x"01",
         10953 => x"01",
         10954 => x"01",
         10955 => x"01",
         10956 => x"01",
         10957 => x"01",
         10958 => x"01",
         10959 => x"01",
         10960 => x"01",
         10961 => x"01",
         10962 => x"01",
         10963 => x"01",
         10964 => x"01",
         10965 => x"01",
         10966 => x"01",
         10967 => x"01",
         10968 => x"01",
         10969 => x"01",
         10970 => x"01",
         10971 => x"01",
         10972 => x"01",
         10973 => x"01",
         10974 => x"01",
         10975 => x"01",
         10976 => x"01",
         10977 => x"01",
         10978 => x"01",
         10979 => x"01",
         10980 => x"01",
         10981 => x"01",
         10982 => x"01",
         10983 => x"01",
         10984 => x"01",
         10985 => x"01",
         10986 => x"01",
         10987 => x"01",
         10988 => x"01",
         10989 => x"01",
         10990 => x"01",
         10991 => x"01",
         10992 => x"00",
         10993 => x"01",
         10994 => x"01",
         10995 => x"02",
         10996 => x"02",
         10997 => x"2c",
         10998 => x"02",
         10999 => x"2c",
         11000 => x"02",
         11001 => x"02",
         11002 => x"01",
         11003 => x"00",
         11004 => x"01",
         11005 => x"01",
         11006 => x"02",
         11007 => x"02",
         11008 => x"02",
         11009 => x"02",
         11010 => x"01",
         11011 => x"02",
         11012 => x"02",
         11013 => x"02",
         11014 => x"01",
         11015 => x"02",
         11016 => x"02",
         11017 => x"02",
         11018 => x"02",
         11019 => x"01",
         11020 => x"02",
         11021 => x"02",
         11022 => x"02",
         11023 => x"02",
         11024 => x"02",
         11025 => x"02",
         11026 => x"01",
         11027 => x"02",
         11028 => x"02",
         11029 => x"02",
         11030 => x"01",
         11031 => x"01",
         11032 => x"02",
         11033 => x"02",
         11034 => x"02",
         11035 => x"01",
         11036 => x"00",
         11037 => x"03",
         11038 => x"03",
         11039 => x"03",
         11040 => x"03",
         11041 => x"03",
         11042 => x"03",
         11043 => x"03",
         11044 => x"03",
         11045 => x"03",
         11046 => x"03",
         11047 => x"03",
         11048 => x"01",
         11049 => x"00",
         11050 => x"03",
         11051 => x"03",
         11052 => x"03",
         11053 => x"03",
         11054 => x"03",
         11055 => x"03",
         11056 => x"07",
         11057 => x"01",
         11058 => x"01",
         11059 => x"01",
         11060 => x"00",
         11061 => x"04",
         11062 => x"05",
         11063 => x"00",
         11064 => x"1d",
         11065 => x"2c",
         11066 => x"01",
         11067 => x"01",
         11068 => x"06",
         11069 => x"06",
         11070 => x"06",
         11071 => x"06",
         11072 => x"06",
         11073 => x"00",
         11074 => x"1f",
         11075 => x"1f",
         11076 => x"1f",
         11077 => x"1f",
         11078 => x"1f",
         11079 => x"1f",
         11080 => x"1f",
         11081 => x"1f",
         11082 => x"1f",
         11083 => x"1f",
         11084 => x"1f",
         11085 => x"1f",
         11086 => x"1f",
         11087 => x"1f",
         11088 => x"1f",
         11089 => x"1f",
         11090 => x"1f",
         11091 => x"1f",
         11092 => x"1f",
         11093 => x"1f",
         11094 => x"06",
         11095 => x"06",
         11096 => x"00",
         11097 => x"1f",
         11098 => x"1f",
         11099 => x"00",
         11100 => x"21",
         11101 => x"21",
         11102 => x"21",
         11103 => x"05",
         11104 => x"04",
         11105 => x"01",
         11106 => x"01",
         11107 => x"01",
         11108 => x"01",
         11109 => x"08",
         11110 => x"03",
         11111 => x"00",
         11112 => x"00",
         11113 => x"01",
         11114 => x"00",
         11115 => x"00",
         11116 => x"00",
         11117 => x"01",
         11118 => x"00",
         11119 => x"00",
         11120 => x"00",
         11121 => x"01",
         11122 => x"00",
         11123 => x"00",
         11124 => x"00",
         11125 => x"01",
         11126 => x"00",
         11127 => x"00",
         11128 => x"00",
         11129 => x"01",
         11130 => x"00",
         11131 => x"00",
         11132 => x"00",
         11133 => x"01",
         11134 => x"00",
         11135 => x"00",
         11136 => x"00",
         11137 => x"01",
         11138 => x"00",
         11139 => x"00",
         11140 => x"00",
         11141 => x"01",
         11142 => x"00",
         11143 => x"00",
         11144 => x"00",
         11145 => x"01",
         11146 => x"00",
         11147 => x"00",
         11148 => x"00",
         11149 => x"01",
         11150 => x"00",
         11151 => x"00",
         11152 => x"00",
         11153 => x"01",
         11154 => x"00",
         11155 => x"00",
         11156 => x"00",
         11157 => x"01",
         11158 => x"00",
         11159 => x"00",
         11160 => x"00",
         11161 => x"01",
         11162 => x"00",
         11163 => x"00",
         11164 => x"00",
         11165 => x"01",
         11166 => x"00",
         11167 => x"00",
         11168 => x"00",
         11169 => x"01",
         11170 => x"00",
         11171 => x"00",
         11172 => x"00",
         11173 => x"01",
         11174 => x"00",
         11175 => x"00",
         11176 => x"00",
         11177 => x"01",
         11178 => x"00",
         11179 => x"00",
         11180 => x"00",
         11181 => x"01",
         11182 => x"00",
         11183 => x"00",
         11184 => x"00",
         11185 => x"01",
         11186 => x"00",
         11187 => x"00",
         11188 => x"00",
         11189 => x"01",
         11190 => x"00",
         11191 => x"00",
         11192 => x"00",
         11193 => x"01",
         11194 => x"00",
         11195 => x"00",
         11196 => x"00",
         11197 => x"01",
         11198 => x"00",
         11199 => x"00",
         11200 => x"00",
         11201 => x"01",
         11202 => x"00",
         11203 => x"00",
         11204 => x"00",
         11205 => x"01",
         11206 => x"00",
         11207 => x"00",
         11208 => x"00",
         11209 => x"01",
         11210 => x"00",
         11211 => x"00",
         11212 => x"00",
         11213 => x"00",
         11214 => x"00",
         11215 => x"00",
         11216 => x"00",
         11217 => x"00",
         11218 => x"00",
         11219 => x"00",
         11220 => x"00",
         11221 => x"01",
         11222 => x"01",
         11223 => x"00",
         11224 => x"00",
         11225 => x"00",
         11226 => x"00",
         11227 => x"05",
         11228 => x"05",
         11229 => x"05",
         11230 => x"00",
         11231 => x"01",
         11232 => x"01",
         11233 => x"01",
         11234 => x"01",
         11235 => x"00",
         11236 => x"00",
         11237 => x"00",
         11238 => x"00",
         11239 => x"00",
         11240 => x"00",
         11241 => x"00",
         11242 => x"00",
         11243 => x"00",
         11244 => x"00",
         11245 => x"00",
         11246 => x"00",
         11247 => x"00",
         11248 => x"00",
         11249 => x"00",
         11250 => x"00",
         11251 => x"00",
         11252 => x"00",
         11253 => x"00",
         11254 => x"00",
         11255 => x"00",
         11256 => x"00",
         11257 => x"00",
         11258 => x"00",
         11259 => x"00",
         11260 => x"01",
         11261 => x"00",
         11262 => x"01",
         11263 => x"00",
         11264 => x"02",
         11265 => x"00",
         11266 => x"00",
         11267 => x"00",
         11268 => x"00",
         11269 => x"01",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(7 downto 0);
                memBRead(7 downto 0) <= memBWrite(7 downto 0);
            else
                memBRead(7 downto 0) <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(15 downto 8);
                memBRead(15 downto 8) <= memBWrite(15 downto 8);
            else
                memBRead(15 downto 8) <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(23 downto 16);
                memBRead(23 downto 16) <= memBWrite(23 downto 16);
            else
                memBRead(23 downto 16) <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2)))) := memBWrite(31 downto 24);
                memBRead(31 downto 24) <= memBWrite(31 downto 24);
            else
                memBRead(31 downto 24) <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

end arch;
