IOCP_SinglePortBootBRAM.vhd