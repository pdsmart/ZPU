ZPUTA_DualPortBootBRAM.vhd