-- Byte Addressed 32bit/64bit BRAM module for the ZPU Evo implementation.
--
-- This template provides a 32bit wide bus on port A and a 64bit bus
-- on port B. This is typically used for the ZPU Boot BRAM where port B
-- is used exclusively for instruction storage.
--
-- Copyright 2018-2021 - Philip Smart for the ZPU Evo implementation.
-- History:
--   20190618  - Initial 32 bit dual port BRAM described by inference rather than
--               using an IP Megacore. This was to make it more portable but also
--               to allow 8/16/32 bit writes to the memory.
--   20210108  - Updated to 64bit on Port B to allow for the 64bit decoder on the ZPU.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity DualPort3264BootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);

        memBAddr             : in  std_logic_vector(addrbits-1 downto 3);
        memBWrite            : in  std_logic_vector(WORD_64BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBRead             : out std_logic_vector(WORD_64BIT_RANGE)
    );
end DualPort3264BootBRAM;

architecture arch of DualPort3264BootBRAM is

    -- Declare 8 byte wide arrays for byte level addressing.
    type ramArray is array(natural range 0 to (2**(addrbits-3))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"fa",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"05",
            10 => x"52",
            11 => x"00",
            12 => x"08",
            13 => x"81",
            14 => x"06",
            15 => x"0b",
            16 => x"05",
            17 => x"06",
            18 => x"06",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"09",
            25 => x"72",
            26 => x"31",
            27 => x"51",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"93",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"2b",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"06",
            45 => x"b4",
            46 => x"00",
            47 => x"00",
            48 => x"ff",
            49 => x"0a",
            50 => x"51",
            51 => x"00",
            52 => x"51",
            53 => x"05",
            54 => x"72",
            55 => x"00",
            56 => x"05",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"05",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"81",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"08",
            77 => x"05",
            78 => x"52",
            79 => x"00",
            80 => x"08",
            81 => x"06",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"d2",
            86 => x"90",
            87 => x"00",
            88 => x"08",
            89 => x"cd",
            90 => x"90",
            91 => x"00",
            92 => x"81",
            93 => x"05",
            94 => x"74",
            95 => x"51",
            96 => x"81",
            97 => x"ff",
            98 => x"72",
            99 => x"51",
           100 => x"04",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"52",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"72",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"ff",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"8c",
           133 => x"04",
           134 => x"0b",
           135 => x"8c",
           136 => x"04",
           137 => x"0b",
           138 => x"8c",
           139 => x"04",
           140 => x"0b",
           141 => x"8d",
           142 => x"04",
           143 => x"0b",
           144 => x"8d",
           145 => x"04",
           146 => x"0b",
           147 => x"8e",
           148 => x"04",
           149 => x"0b",
           150 => x"8f",
           151 => x"04",
           152 => x"0b",
           153 => x"8f",
           154 => x"04",
           155 => x"0b",
           156 => x"90",
           157 => x"04",
           158 => x"0b",
           159 => x"90",
           160 => x"04",
           161 => x"0b",
           162 => x"91",
           163 => x"04",
           164 => x"0b",
           165 => x"91",
           166 => x"04",
           167 => x"0b",
           168 => x"92",
           169 => x"04",
           170 => x"0b",
           171 => x"92",
           172 => x"04",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"81",
           193 => x"8b",
           194 => x"80",
           195 => x"e6",
           196 => x"80",
           197 => x"97",
           198 => x"80",
           199 => x"e1",
           200 => x"80",
           201 => x"e1",
           202 => x"80",
           203 => x"f6",
           204 => x"80",
           205 => x"da",
           206 => x"c0",
           207 => x"80",
           208 => x"80",
           209 => x"0c",
           210 => x"80",
           211 => x"0c",
           212 => x"80",
           213 => x"0c",
           214 => x"80",
           215 => x"0c",
           216 => x"08",
           217 => x"a4",
           218 => x"a4",
           219 => x"e0",
           220 => x"e0",
           221 => x"82",
           222 => x"82",
           223 => x"04",
           224 => x"2d",
           225 => x"90",
           226 => x"a7",
           227 => x"80",
           228 => x"83",
           229 => x"c0",
           230 => x"81",
           231 => x"80",
           232 => x"0c",
           233 => x"08",
           234 => x"a4",
           235 => x"a4",
           236 => x"e0",
           237 => x"e0",
           238 => x"82",
           239 => x"82",
           240 => x"04",
           241 => x"2d",
           242 => x"90",
           243 => x"a8",
           244 => x"80",
           245 => x"8d",
           246 => x"c0",
           247 => x"82",
           248 => x"80",
           249 => x"0c",
           250 => x"08",
           251 => x"a4",
           252 => x"a4",
           253 => x"e0",
           254 => x"e0",
           255 => x"82",
           256 => x"82",
           257 => x"04",
           258 => x"2d",
           259 => x"90",
           260 => x"87",
           261 => x"80",
           262 => x"83",
           263 => x"c0",
           264 => x"82",
           265 => x"80",
           266 => x"0c",
           267 => x"08",
           268 => x"a4",
           269 => x"a4",
           270 => x"e0",
           271 => x"e0",
           272 => x"82",
           273 => x"82",
           274 => x"04",
           275 => x"2d",
           276 => x"90",
           277 => x"8c",
           278 => x"80",
           279 => x"b4",
           280 => x"c0",
           281 => x"82",
           282 => x"80",
           283 => x"0c",
           284 => x"08",
           285 => x"a4",
           286 => x"a4",
           287 => x"e0",
           288 => x"e0",
           289 => x"82",
           290 => x"82",
           291 => x"04",
           292 => x"2d",
           293 => x"90",
           294 => x"80",
           295 => x"80",
           296 => x"e0",
           297 => x"c0",
           298 => x"81",
           299 => x"80",
           300 => x"0c",
           301 => x"08",
           302 => x"a4",
           303 => x"a4",
           304 => x"e0",
           305 => x"e0",
           306 => x"3c",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"10",
           311 => x"ff",
           312 => x"83",
           313 => x"fc",
           314 => x"80",
           315 => x"06",
           316 => x"0a",
           317 => x"51",
           318 => x"84",
           319 => x"05",
           320 => x"04",
           321 => x"00",
           322 => x"a4",
           323 => x"08",
           324 => x"fc",
           325 => x"05",
           326 => x"05",
           327 => x"54",
           328 => x"70",
           329 => x"82",
           330 => x"82",
           331 => x"0d",
           332 => x"a4",
           333 => x"3d",
           334 => x"08",
           335 => x"81",
           336 => x"38",
           337 => x"05",
           338 => x"0b",
           339 => x"81",
           340 => x"05",
           341 => x"8c",
           342 => x"08",
           343 => x"88",
           344 => x"05",
           345 => x"08",
           346 => x"82",
           347 => x"80",
           348 => x"05",
           349 => x"98",
           350 => x"05",
           351 => x"05",
           352 => x"38",
           353 => x"05",
           354 => x"08",
           355 => x"f8",
           356 => x"82",
           357 => x"05",
           358 => x"82",
           359 => x"05",
           360 => x"ff",
           361 => x"05",
           362 => x"a4",
           363 => x"a4",
           364 => x"a4",
           365 => x"0c",
           366 => x"04",
           367 => x"a4",
           368 => x"e0",
           369 => x"a4",
           370 => x"08",
           371 => x"e0",
           372 => x"a4",
           373 => x"08",
           374 => x"fc",
           375 => x"8c",
           376 => x"e0",
           377 => x"3f",
           378 => x"a4",
           379 => x"08",
           380 => x"88",
           381 => x"34",
           382 => x"70",
           383 => x"0d",
           384 => x"a4",
           385 => x"3d",
           386 => x"70",
           387 => x"82",
           388 => x"82",
           389 => x"82",
           390 => x"54",
           391 => x"82",
           392 => x"e0",
           393 => x"e0",
           394 => x"82",
           395 => x"08",
           396 => x"0d",
           397 => x"05",
           398 => x"08",
           399 => x"e0",
           400 => x"33",
           401 => x"81",
           402 => x"80",
           403 => x"a4",
           404 => x"82",
           405 => x"72",
           406 => x"f8",
           407 => x"72",
           408 => x"a4",
           409 => x"e0",
           410 => x"a4",
           411 => x"51",
           412 => x"82",
           413 => x"af",
           414 => x"a4",
           415 => x"26",
           416 => x"f8",
           417 => x"81",
           418 => x"08",
           419 => x"98",
           420 => x"82",
           421 => x"83",
           422 => x"51",
           423 => x"38",
           424 => x"70",
           425 => x"e0",
           426 => x"39",
           427 => x"70",
           428 => x"83",
           429 => x"51",
           430 => x"a4",
           431 => x"08",
           432 => x"08",
           433 => x"51",
           434 => x"e8",
           435 => x"05",
           436 => x"51",
           437 => x"80",
           438 => x"05",
           439 => x"22",
           440 => x"51",
           441 => x"a4",
           442 => x"70",
           443 => x"2c",
           444 => x"e0",
           445 => x"39",
           446 => x"70",
           447 => x"53",
           448 => x"a4",
           449 => x"70",
           450 => x"38",
           451 => x"05",
           452 => x"33",
           453 => x"05",
           454 => x"05",
           455 => x"82",
           456 => x"82",
           457 => x"51",
           458 => x"a4",
           459 => x"51",
           460 => x"05",
           461 => x"22",
           462 => x"e0",
           463 => x"39",
           464 => x"70",
           465 => x"e0",
           466 => x"39",
           467 => x"70",
           468 => x"e0",
           469 => x"39",
           470 => x"70",
           471 => x"a4",
           472 => x"e0",
           473 => x"39",
           474 => x"70",
           475 => x"a4",
           476 => x"bf",
           477 => x"34",
           478 => x"ff",
           479 => x"08",
           480 => x"e0",
           481 => x"39",
           482 => x"82",
           483 => x"05",
           484 => x"70",
           485 => x"08",
           486 => x"ec",
           487 => x"82",
           488 => x"ef",
           489 => x"08",
           490 => x"84",
           491 => x"0c",
           492 => x"05",
           493 => x"22",
           494 => x"51",
           495 => x"82",
           496 => x"98",
           497 => x"e0",
           498 => x"a4",
           499 => x"72",
           500 => x"99",
           501 => x"08",
           502 => x"08",
           503 => x"05",
           504 => x"22",
           505 => x"22",
           506 => x"e0",
           507 => x"39",
           508 => x"82",
           509 => x"05",
           510 => x"70",
           511 => x"0c",
           512 => x"70",
           513 => x"51",
           514 => x"e0",
           515 => x"2b",
           516 => x"a4",
           517 => x"ec",
           518 => x"82",
           519 => x"39",
           520 => x"51",
           521 => x"53",
           522 => x"23",
           523 => x"53",
           524 => x"73",
           525 => x"a4",
           526 => x"82",
           527 => x"82",
           528 => x"72",
           529 => x"08",
           530 => x"90",
           531 => x"08",
           532 => x"a4",
           533 => x"82",
           534 => x"e0",
           535 => x"82",
           536 => x"08",
           537 => x"53",
           538 => x"82",
           539 => x"e0",
           540 => x"a4",
           541 => x"22",
           542 => x"e0",
           543 => x"a4",
           544 => x"a4",
           545 => x"08",
           546 => x"51",
           547 => x"05",
           548 => x"e0",
           549 => x"82",
           550 => x"80",
           551 => x"a4",
           552 => x"82",
           553 => x"0b",
           554 => x"82",
           555 => x"82",
           556 => x"72",
           557 => x"08",
           558 => x"90",
           559 => x"08",
           560 => x"a4",
           561 => x"82",
           562 => x"e0",
           563 => x"82",
           564 => x"08",
           565 => x"53",
           566 => x"82",
           567 => x"e0",
           568 => x"06",
           569 => x"e4",
           570 => x"e0",
           571 => x"a4",
           572 => x"08",
           573 => x"fc",
           574 => x"54",
           575 => x"08",
           576 => x"08",
           577 => x"d4",
           578 => x"05",
           579 => x"27",
           580 => x"05",
           581 => x"a4",
           582 => x"11",
           583 => x"08",
           584 => x"a4",
           585 => x"b0",
           586 => x"08",
           587 => x"d4",
           588 => x"d0",
           589 => x"08",
           590 => x"a4",
           591 => x"08",
           592 => x"a4",
           593 => x"c7",
           594 => x"e0",
           595 => x"e0",
           596 => x"84",
           597 => x"08",
           598 => x"55",
           599 => x"53",
           600 => x"34",
           601 => x"70",
           602 => x"94",
           603 => x"22",
           604 => x"a4",
           605 => x"08",
           606 => x"81",
           607 => x"80",
           608 => x"05",
           609 => x"08",
           610 => x"cc",
           611 => x"08",
           612 => x"f4",
           613 => x"09",
           614 => x"08",
           615 => x"82",
           616 => x"39",
           617 => x"ff",
           618 => x"c8",
           619 => x"05",
           620 => x"23",
           621 => x"70",
           622 => x"53",
           623 => x"e0",
           624 => x"2b",
           625 => x"fc",
           626 => x"74",
           627 => x"e4",
           628 => x"72",
           629 => x"9d",
           630 => x"33",
           631 => x"33",
           632 => x"e0",
           633 => x"a4",
           634 => x"70",
           635 => x"2e",
           636 => x"05",
           637 => x"70",
           638 => x"51",
           639 => x"08",
           640 => x"53",
           641 => x"23",
           642 => x"05",
           643 => x"70",
           644 => x"51",
           645 => x"08",
           646 => x"53",
           647 => x"23",
           648 => x"70",
           649 => x"38",
           650 => x"ff",
           651 => x"08",
           652 => x"90",
           653 => x"38",
           654 => x"52",
           655 => x"82",
           656 => x"81",
           657 => x"72",
           658 => x"08",
           659 => x"ca",
           660 => x"08",
           661 => x"81",
           662 => x"90",
           663 => x"08",
           664 => x"39",
           665 => x"70",
           666 => x"53",
           667 => x"a4",
           668 => x"8a",
           669 => x"05",
           670 => x"51",
           671 => x"82",
           672 => x"b0",
           673 => x"08",
           674 => x"09",
           675 => x"08",
           676 => x"08",
           677 => x"82",
           678 => x"88",
           679 => x"72",
           680 => x"08",
           681 => x"72",
           682 => x"73",
           683 => x"80",
           684 => x"08",
           685 => x"fa",
           686 => x"e4",
           687 => x"06",
           688 => x"38",
           689 => x"ff",
           690 => x"08",
           691 => x"98",
           692 => x"38",
           693 => x"52",
           694 => x"82",
           695 => x"87",
           696 => x"72",
           697 => x"05",
           698 => x"e0",
           699 => x"2b",
           700 => x"25",
           701 => x"05",
           702 => x"d2",
           703 => x"33",
           704 => x"06",
           705 => x"05",
           706 => x"05",
           707 => x"39",
           708 => x"53",
           709 => x"80",
           710 => x"05",
           711 => x"e0",
           712 => x"ff",
           713 => x"2e",
           714 => x"88",
           715 => x"fc",
           716 => x"a4",
           717 => x"e0",
           718 => x"f2",
           719 => x"08",
           720 => x"2e",
           721 => x"e0",
           722 => x"51",
           723 => x"05",
           724 => x"72",
           725 => x"82",
           726 => x"82",
           727 => x"33",
           728 => x"a4",
           729 => x"e0",
           730 => x"39",
           731 => x"82",
           732 => x"a4",
           733 => x"a4",
           734 => x"e0",
           735 => x"a4",
           736 => x"53",
           737 => x"a4",
           738 => x"70",
           739 => x"2e",
           740 => x"ec",
           741 => x"82",
           742 => x"90",
           743 => x"73",
           744 => x"88",
           745 => x"3f",
           746 => x"05",
           747 => x"05",
           748 => x"82",
           749 => x"b7",
           750 => x"33",
           751 => x"a8",
           752 => x"e4",
           753 => x"08",
           754 => x"a4",
           755 => x"e0",
           756 => x"39",
           757 => x"52",
           758 => x"51",
           759 => x"e0",
           760 => x"08",
           761 => x"0c",
           762 => x"05",
           763 => x"0d",
           764 => x"a4",
           765 => x"3d",
           766 => x"e0",
           767 => x"e0",
           768 => x"dd",
           769 => x"e0",
           770 => x"e0",
           771 => x"02",
           772 => x"80",
           773 => x"0c",
           774 => x"70",
           775 => x"06",
           776 => x"2e",
           777 => x"08",
           778 => x"e0",
           779 => x"33",
           780 => x"81",
           781 => x"0c",
           782 => x"05",
           783 => x"80",
           784 => x"82",
           785 => x"08",
           786 => x"51",
           787 => x"53",
           788 => x"0b",
           789 => x"ff",
           790 => x"fb",
           791 => x"13",
           792 => x"08",
           793 => x"0b",
           794 => x"82",
           795 => x"82",
           796 => x"82",
           797 => x"e0",
           798 => x"a4",
           799 => x"82",
           800 => x"0b",
           801 => x"82",
           802 => x"11",
           803 => x"70",
           804 => x"72",
           805 => x"e0",
           806 => x"39",
           807 => x"53",
           808 => x"05",
           809 => x"88",
           810 => x"08",
           811 => x"53",
           812 => x"a4",
           813 => x"08",
           814 => x"08",
           815 => x"51",
           816 => x"53",
           817 => x"0b",
           818 => x"ff",
           819 => x"05",
           820 => x"05",
           821 => x"05",
           822 => x"0d",
           823 => x"a4",
           824 => x"3d",
           825 => x"e0",
           826 => x"3f",
           827 => x"98",
           828 => x"a4",
           829 => x"82",
           830 => x"e0",
           831 => x"33",
           832 => x"81",
           833 => x"80",
           834 => x"a4",
           835 => x"82",
           836 => x"11",
           837 => x"51",
           838 => x"db",
           839 => x"08",
           840 => x"54",
           841 => x"25",
           842 => x"05",
           843 => x"08",
           844 => x"72",
           845 => x"0c",
           846 => x"8c",
           847 => x"82",
           848 => x"82",
           849 => x"53",
           850 => x"8c",
           851 => x"05",
           852 => x"05",
           853 => x"12",
           854 => x"e0",
           855 => x"e0",
           856 => x"08",
           857 => x"a4",
           858 => x"a4",
           859 => x"39",
           860 => x"05",
           861 => x"08",
           862 => x"82",
           863 => x"08",
           864 => x"0d",
           865 => x"85",
           866 => x"06",
           867 => x"8d",
           868 => x"f8",
           869 => x"a4",
           870 => x"70",
           871 => x"51",
           872 => x"82",
           873 => x"e0",
           874 => x"85",
           875 => x"52",
           876 => x"08",
           877 => x"05",
           878 => x"88",
           879 => x"e0",
           880 => x"52",
           881 => x"88",
           882 => x"2a",
           883 => x"71",
           884 => x"a4",
           885 => x"33",
           886 => x"51",
           887 => x"08",
           888 => x"05",
           889 => x"08",
           890 => x"07",
           891 => x"0b",
           892 => x"81",
           893 => x"05",
           894 => x"52",
           895 => x"88",
           896 => x"05",
           897 => x"71",
           898 => x"e0",
           899 => x"e0",
           900 => x"80",
           901 => x"05",
           902 => x"0c",
           903 => x"85",
           904 => x"05",
           905 => x"05",
           906 => x"38",
           907 => x"90",
           908 => x"ec",
           909 => x"08",
           910 => x"82",
           911 => x"e0",
           912 => x"e0",
           913 => x"34",
           914 => x"05",
           915 => x"88",
           916 => x"8c",
           917 => x"05",
           918 => x"e0",
           919 => x"52",
           920 => x"82",
           921 => x"e0",
           922 => x"02",
           923 => x"82",
           924 => x"e0",
           925 => x"a4",
           926 => x"08",
           927 => x"90",
           928 => x"82",
           929 => x"e0",
           930 => x"ac",
           931 => x"08",
           932 => x"05",
           933 => x"08",
           934 => x"a4",
           935 => x"08",
           936 => x"08",
           937 => x"f8",
           938 => x"05",
           939 => x"05",
           940 => x"08",
           941 => x"05",
           942 => x"08",
           943 => x"05",
           944 => x"08",
           945 => x"a4",
           946 => x"e0",
           947 => x"a4",
           948 => x"e0",
           949 => x"a4",
           950 => x"08",
           951 => x"71",
           952 => x"08",
           953 => x"a4",
           954 => x"08",
           955 => x"a4",
           956 => x"08",
           957 => x"82",
           958 => x"70",
           959 => x"08",
           960 => x"05",
           961 => x"08",
           962 => x"a4",
           963 => x"e0",
           964 => x"39",
           965 => x"70",
           966 => x"0d",
           967 => x"a4",
           968 => x"3d",
           969 => x"08",
           970 => x"82",
           971 => x"71",
           972 => x"08",
           973 => x"05",
           974 => x"70",
           975 => x"e0",
           976 => x"82",
           977 => x"e0",
           978 => x"a4",
           979 => x"e0",
           980 => x"e0",
           981 => x"02",
           982 => x"82",
           983 => x"e0",
           984 => x"a4",
           985 => x"82",
           986 => x"05",
           987 => x"82",
           988 => x"51",
           989 => x"fc",
           990 => x"08",
           991 => x"51",
           992 => x"39",
           993 => x"70",
           994 => x"0d",
           995 => x"a4",
           996 => x"3d",
           997 => x"08",
           998 => x"82",
           999 => x"e0",
          1000 => x"a4",
          1001 => x"e5",
          1002 => x"08",
          1003 => x"05",
          1004 => x"08",
          1005 => x"05",
          1006 => x"08",
          1007 => x"08",
          1008 => x"e0",
          1009 => x"82",
          1010 => x"e0",
          1011 => x"71",
          1012 => x"05",
          1013 => x"fc",
          1014 => x"a4",
          1015 => x"98",
          1016 => x"a4",
          1017 => x"82",
          1018 => x"e0",
          1019 => x"81",
          1020 => x"05",
          1021 => x"08",
          1022 => x"a4",
          1023 => x"08",
          1024 => x"ff",
          1025 => x"2e",
          1026 => x"a4",
          1027 => x"82",
          1028 => x"05",
          1029 => x"70",
          1030 => x"38",
          1031 => x"05",
          1032 => x"08",
          1033 => x"a4",
          1034 => x"08",
          1035 => x"ff",
          1036 => x"05",
          1037 => x"e0",
          1038 => x"52",
          1039 => x"e0",
          1040 => x"39",
          1041 => x"ff",
          1042 => x"0c",
          1043 => x"70",
          1044 => x"0b",
          1045 => x"ae",
          1046 => x"08",
          1047 => x"05",
          1048 => x"82",
          1049 => x"55",
          1050 => x"82",
          1051 => x"e0",
          1052 => x"98",
          1053 => x"0c",
          1054 => x"e0",
          1055 => x"a4",
          1056 => x"a4",
          1057 => x"3f",
          1058 => x"a4",
          1059 => x"08",
          1060 => x"51",
          1061 => x"98",
          1062 => x"05",
          1063 => x"05",
          1064 => x"a4",
          1065 => x"e0",
          1066 => x"a4",
          1067 => x"74",
          1068 => x"08",
          1069 => x"08",
          1070 => x"08",
          1071 => x"08",
          1072 => x"0c",
          1073 => x"08",
          1074 => x"82",
          1075 => x"08",
          1076 => x"0d",
          1077 => x"82",
          1078 => x"e0",
          1079 => x"80",
          1080 => x"0c",
          1081 => x"f8",
          1082 => x"a4",
          1083 => x"e0",
          1084 => x"ff",
          1085 => x"38",
          1086 => x"ff",
          1087 => x"0c",
          1088 => x"ff",
          1089 => x"e0",
          1090 => x"82",
          1091 => x"e0",
          1092 => x"a4",
          1093 => x"e0",
          1094 => x"e0",
          1095 => x"98",
          1096 => x"0c",
          1097 => x"e0",
          1098 => x"a4",
          1099 => x"08",
          1100 => x"90",
          1101 => x"82",
          1102 => x"05",
          1103 => x"82",
          1104 => x"05",
          1105 => x"82",
          1106 => x"2e",
          1107 => x"05",
          1108 => x"fc",
          1109 => x"82",
          1110 => x"05",
          1111 => x"ff",
          1112 => x"05",
          1113 => x"84",
          1114 => x"82",
          1115 => x"0c",
          1116 => x"8c",
          1117 => x"88",
          1118 => x"98",
          1119 => x"84",
          1120 => x"82",
          1121 => x"0c",
          1122 => x"a4",
          1123 => x"08",
          1124 => x"82",
          1125 => x"83",
          1126 => x"82",
          1127 => x"8f",
          1128 => x"08",
          1129 => x"82",
          1130 => x"2e",
          1131 => x"05",
          1132 => x"98",
          1133 => x"08",
          1134 => x"05",
          1135 => x"08",
          1136 => x"fc",
          1137 => x"e0",
          1138 => x"05",
          1139 => x"0c",
          1140 => x"ff",
          1141 => x"f8",
          1142 => x"82",
          1143 => x"da",
          1144 => x"08",
          1145 => x"08",
          1146 => x"94",
          1147 => x"08",
          1148 => x"0c",
          1149 => x"08",
          1150 => x"a4",
          1151 => x"08",
          1152 => x"f8",
          1153 => x"f4",
          1154 => x"05",
          1155 => x"08",
          1156 => x"08",
          1157 => x"05",
          1158 => x"08",
          1159 => x"f8",
          1160 => x"82",
          1161 => x"82",
          1162 => x"05",
          1163 => x"71",
          1164 => x"08",
          1165 => x"88",
          1166 => x"08",
          1167 => x"08",
          1168 => x"8c",
          1169 => x"05",
          1170 => x"08",
          1171 => x"2c",
          1172 => x"82",
          1173 => x"06",
          1174 => x"82",
          1175 => x"e0",
          1176 => x"e0",
          1177 => x"82",
          1178 => x"e0",
          1179 => x"82",
          1180 => x"52",
          1181 => x"cb",
          1182 => x"08",
          1183 => x"05",
          1184 => x"05",
          1185 => x"08",
          1186 => x"0c",
          1187 => x"05",
          1188 => x"0d",
          1189 => x"a4",
          1190 => x"3d",
          1191 => x"08",
          1192 => x"82",
          1193 => x"80",
          1194 => x"0b",
          1195 => x"8a",
          1196 => x"f0",
          1197 => x"05",
          1198 => x"0c",
          1199 => x"05",
          1200 => x"05",
          1201 => x"fc",
          1202 => x"05",
          1203 => x"0c",
          1204 => x"83",
          1205 => x"38",
          1206 => x"05",
          1207 => x"a4",
          1208 => x"08",
          1209 => x"f8",
          1210 => x"08",
          1211 => x"08",
          1212 => x"a4",
          1213 => x"08",
          1214 => x"f8",
          1215 => x"f4",
          1216 => x"05",
          1217 => x"8c",
          1218 => x"e8",
          1219 => x"e0",
          1220 => x"a4",
          1221 => x"08",
          1222 => x"a4",
          1223 => x"a4",
          1224 => x"e0",
          1225 => x"a4",
          1226 => x"08",
          1227 => x"08",
          1228 => x"fc",
          1229 => x"8c",
          1230 => x"e4",
          1231 => x"e0",
          1232 => x"a4",
          1233 => x"08",
          1234 => x"a4",
          1235 => x"a4",
          1236 => x"e0",
          1237 => x"a4",
          1238 => x"08",
          1239 => x"08",
          1240 => x"a4",
          1241 => x"a4",
          1242 => x"81",
          1243 => x"75",
          1244 => x"08",
          1245 => x"53",
          1246 => x"51",
          1247 => x"04",
          1248 => x"a4",
          1249 => x"08",
          1250 => x"08",
          1251 => x"82",
          1252 => x"08",
          1253 => x"08",
          1254 => x"e0",
          1255 => x"0d",
          1256 => x"a4",
          1257 => x"3d",
          1258 => x"08",
          1259 => x"08",
          1260 => x"70",
          1261 => x"0d",
          1262 => x"a4",
          1263 => x"3d",
          1264 => x"fc",
          1265 => x"05",
          1266 => x"a4",
          1267 => x"3f",
          1268 => x"a4",
          1269 => x"82",
          1270 => x"e0",
          1271 => x"a4",
          1272 => x"38",
          1273 => x"51",
          1274 => x"82",
          1275 => x"31",
          1276 => x"52",
          1277 => x"05",
          1278 => x"08",
          1279 => x"0c",
          1280 => x"82",
          1281 => x"e0",
          1282 => x"52",
          1283 => x"08",
          1284 => x"88",
          1285 => x"e8",
          1286 => x"e0",
          1287 => x"52",
          1288 => x"08",
          1289 => x"0b",
          1290 => x"82",
          1291 => x"05",
          1292 => x"f8",
          1293 => x"05",
          1294 => x"08",
          1295 => x"0c",
          1296 => x"82",
          1297 => x"82",
          1298 => x"2b",
          1299 => x"52",
          1300 => x"05",
          1301 => x"08",
          1302 => x"a4",
          1303 => x"a4",
          1304 => x"e0",
          1305 => x"70",
          1306 => x"05",
          1307 => x"08",
          1308 => x"05",
          1309 => x"05",
          1310 => x"08",
          1311 => x"31",
          1312 => x"05",
          1313 => x"e0",
          1314 => x"a4",
          1315 => x"e0",
          1316 => x"a4",
          1317 => x"08",
          1318 => x"08",
          1319 => x"a4",
          1320 => x"08",
          1321 => x"a4",
          1322 => x"51",
          1323 => x"82",
          1324 => x"82",
          1325 => x"82",
          1326 => x"e0",
          1327 => x"a4",
          1328 => x"82",
          1329 => x"0b",
          1330 => x"82",
          1331 => x"e0",
          1332 => x"e0",
          1333 => x"a4",
          1334 => x"08",
          1335 => x"08",
          1336 => x"88",
          1337 => x"05",
          1338 => x"f8",
          1339 => x"88",
          1340 => x"05",
          1341 => x"08",
          1342 => x"05",
          1343 => x"05",
          1344 => x"08",
          1345 => x"32",
          1346 => x"82",
          1347 => x"82",
          1348 => x"51",
          1349 => x"08",
          1350 => x"08",
          1351 => x"05",
          1352 => x"51",
          1353 => x"a4",
          1354 => x"82",
          1355 => x"0b",
          1356 => x"82",
          1357 => x"80",
          1358 => x"05",
          1359 => x"53",
          1360 => x"34",
          1361 => x"2e",
          1362 => x"a4",
          1363 => x"05",
          1364 => x"a4",
          1365 => x"2e",
          1366 => x"82",
          1367 => x"e0",
          1368 => x"81",
          1369 => x"72",
          1370 => x"34",
          1371 => x"53",
          1372 => x"dc",
          1373 => x"08",
          1374 => x"08",
          1375 => x"08",
          1376 => x"f8",
          1377 => x"05",
          1378 => x"08",
          1379 => x"a4",
          1380 => x"84",
          1381 => x"e0",
          1382 => x"a4",
          1383 => x"05",
          1384 => x"33",
          1385 => x"81",
          1386 => x"08",
          1387 => x"88",
          1388 => x"0c",
          1389 => x"e0",
          1390 => x"39",
          1391 => x"53",
          1392 => x"82",
          1393 => x"80",
          1394 => x"33",
          1395 => x"e0",
          1396 => x"b9",
          1397 => x"82",
          1398 => x"d8",
          1399 => x"f4",
          1400 => x"08",
          1401 => x"90",
          1402 => x"33",
          1403 => x"39",
          1404 => x"05",
          1405 => x"e0",
          1406 => x"82",
          1407 => x"e0",
          1408 => x"73",
          1409 => x"08",
          1410 => x"27",
          1411 => x"05",
          1412 => x"e0",
          1413 => x"a4",
          1414 => x"53",
          1415 => x"34",
          1416 => x"53",
          1417 => x"a4",
          1418 => x"53",
          1419 => x"34",
          1420 => x"53",
          1421 => x"82",
          1422 => x"98",
          1423 => x"33",
          1424 => x"54",
          1425 => x"0b",
          1426 => x"80",
          1427 => x"05",
          1428 => x"05",
          1429 => x"05",
          1430 => x"fc",
          1431 => x"05",
          1432 => x"70",
          1433 => x"33",
          1434 => x"fe",
          1435 => x"05",
          1436 => x"82",
          1437 => x"82",
          1438 => x"e0",
          1439 => x"a4",
          1440 => x"81",
          1441 => x"0c",
          1442 => x"82",
          1443 => x"e0",
          1444 => x"02",
          1445 => x"80",
          1446 => x"34",
          1447 => x"53",
          1448 => x"88",
          1449 => x"33",
          1450 => x"05",
          1451 => x"a0",
          1452 => x"e0",
          1453 => x"81",
          1454 => x"e0",
          1455 => x"ad",
          1456 => x"0b",
          1457 => x"82",
          1458 => x"08",
          1459 => x"53",
          1460 => x"05",
          1461 => x"33",
          1462 => x"81",
          1463 => x"05",
          1464 => x"70",
          1465 => x"a4",
          1466 => x"08",
          1467 => x"e8",
          1468 => x"05",
          1469 => x"e0",
          1470 => x"2e",
          1471 => x"82",
          1472 => x"e0",
          1473 => x"81",
          1474 => x"72",
          1475 => x"34",
          1476 => x"a4",
          1477 => x"08",
          1478 => x"71",
          1479 => x"82",
          1480 => x"fe",
          1481 => x"33",
          1482 => x"0b",
          1483 => x"83",
          1484 => x"05",
          1485 => x"82",
          1486 => x"72",
          1487 => x"0b",
          1488 => x"82",
          1489 => x"08",
          1490 => x"a4",
          1491 => x"27",
          1492 => x"05",
          1493 => x"8d",
          1494 => x"ec",
          1495 => x"82",
          1496 => x"0b",
          1497 => x"82",
          1498 => x"a0",
          1499 => x"a4",
          1500 => x"73",
          1501 => x"f8",
          1502 => x"82",
          1503 => x"e0",
          1504 => x"51",
          1505 => x"05",
          1506 => x"33",
          1507 => x"e0",
          1508 => x"51",
          1509 => x"05",
          1510 => x"33",
          1511 => x"0b",
          1512 => x"81",
          1513 => x"05",
          1514 => x"33",
          1515 => x"80",
          1516 => x"0c",
          1517 => x"f4",
          1518 => x"fc",
          1519 => x"f8",
          1520 => x"08",
          1521 => x"88",
          1522 => x"0c",
          1523 => x"72",
          1524 => x"34",
          1525 => x"f0",
          1526 => x"38",
          1527 => x"30",
          1528 => x"82",
          1529 => x"e0",
          1530 => x"53",
          1531 => x"05",
          1532 => x"08",
          1533 => x"82",
          1534 => x"7a",
          1535 => x"80",
          1536 => x"15",
          1537 => x"d2",
          1538 => x"09",
          1539 => x"f1",
          1540 => x"db",
          1541 => x"8d",
          1542 => x"98",
          1543 => x"58",
          1544 => x"8b",
          1545 => x"2e",
          1546 => x"ff",
          1547 => x"38",
          1548 => x"8a",
          1549 => x"e0",
          1550 => x"52",
          1551 => x"84",
          1552 => x"08",
          1553 => x"39",
          1554 => x"82",
          1555 => x"be",
          1556 => x"a0",
          1557 => x"51",
          1558 => x"80",
          1559 => x"cf",
          1560 => x"39",
          1561 => x"82",
          1562 => x"b8",
          1563 => x"af",
          1564 => x"82",
          1565 => x"a4",
          1566 => x"97",
          1567 => x"82",
          1568 => x"fc",
          1569 => x"ce",
          1570 => x"3d",
          1571 => x"e7",
          1572 => x"e8",
          1573 => x"74",
          1574 => x"08",
          1575 => x"e0",
          1576 => x"82",
          1577 => x"87",
          1578 => x"02",
          1579 => x"57",
          1580 => x"73",
          1581 => x"77",
          1582 => x"74",
          1583 => x"55",
          1584 => x"53",
          1585 => x"81",
          1586 => x"57",
          1587 => x"e0",
          1588 => x"82",
          1589 => x"05",
          1590 => x"51",
          1591 => x"08",
          1592 => x"7a",
          1593 => x"19",
          1594 => x"3d",
          1595 => x"76",
          1596 => x"30",
          1597 => x"51",
          1598 => x"c1",
          1599 => x"52",
          1600 => x"75",
          1601 => x"04",
          1602 => x"b7",
          1603 => x"53",
          1604 => x"82",
          1605 => x"2e",
          1606 => x"9c",
          1607 => x"60",
          1608 => x"7e",
          1609 => x"58",
          1610 => x"98",
          1611 => x"0d",
          1612 => x"cf",
          1613 => x"5f",
          1614 => x"38",
          1615 => x"81",
          1616 => x"2e",
          1617 => x"2e",
          1618 => x"d2",
          1619 => x"c4",
          1620 => x"cc",
          1621 => x"74",
          1622 => x"2e",
          1623 => x"80",
          1624 => x"27",
          1625 => x"d0",
          1626 => x"82",
          1627 => x"82",
          1628 => x"53",
          1629 => x"52",
          1630 => x"3f",
          1631 => x"ae",
          1632 => x"74",
          1633 => x"72",
          1634 => x"ad",
          1635 => x"51",
          1636 => x"82",
          1637 => x"ba",
          1638 => x"51",
          1639 => x"78",
          1640 => x"33",
          1641 => x"83",
          1642 => x"27",
          1643 => x"70",
          1644 => x"2e",
          1645 => x"38",
          1646 => x"88",
          1647 => x"51",
          1648 => x"b6",
          1649 => x"3f",
          1650 => x"51",
          1651 => x"98",
          1652 => x"a0",
          1653 => x"51",
          1654 => x"98",
          1655 => x"70",
          1656 => x"72",
          1657 => x"58",
          1658 => x"d6",
          1659 => x"7c",
          1660 => x"38",
          1661 => x"8f",
          1662 => x"9b",
          1663 => x"3f",
          1664 => x"51",
          1665 => x"22",
          1666 => x"54",
          1667 => x"33",
          1668 => x"e8",
          1669 => x"89",
          1670 => x"0d",
          1671 => x"f4",
          1672 => x"c2",
          1673 => x"99",
          1674 => x"06",
          1675 => x"81",
          1676 => x"51",
          1677 => x"3f",
          1678 => x"52",
          1679 => x"99",
          1680 => x"98",
          1681 => x"83",
          1682 => x"80",
          1683 => x"3f",
          1684 => x"80",
          1685 => x"70",
          1686 => x"92",
          1687 => x"c3",
          1688 => x"98",
          1689 => x"06",
          1690 => x"81",
          1691 => x"51",
          1692 => x"3f",
          1693 => x"52",
          1694 => x"98",
          1695 => x"a0",
          1696 => x"87",
          1697 => x"80",
          1698 => x"3f",
          1699 => x"80",
          1700 => x"70",
          1701 => x"92",
          1702 => x"c3",
          1703 => x"97",
          1704 => x"0d",
          1705 => x"05",
          1706 => x"80",
          1707 => x"0b",
          1708 => x"38",
          1709 => x"f7",
          1710 => x"e0",
          1711 => x"08",
          1712 => x"51",
          1713 => x"34",
          1714 => x"73",
          1715 => x"82",
          1716 => x"81",
          1717 => x"80",
          1718 => x"51",
          1719 => x"a8",
          1720 => x"0b",
          1721 => x"82",
          1722 => x"09",
          1723 => x"53",
          1724 => x"80",
          1725 => x"0d",
          1726 => x"5e",
          1727 => x"81",
          1728 => x"82",
          1729 => x"78",
          1730 => x"97",
          1731 => x"52",
          1732 => x"78",
          1733 => x"9a",
          1734 => x"88",
          1735 => x"39",
          1736 => x"51",
          1737 => x"47",
          1738 => x"f1",
          1739 => x"f3",
          1740 => x"2b",
          1741 => x"c2",
          1742 => x"24",
          1743 => x"38",
          1744 => x"2e",
          1745 => x"da",
          1746 => x"2e",
          1747 => x"85",
          1748 => x"38",
          1749 => x"89",
          1750 => x"38",
          1751 => x"78",
          1752 => x"a7",
          1753 => x"38",
          1754 => x"81",
          1755 => x"39",
          1756 => x"8a",
          1757 => x"53",
          1758 => x"82",
          1759 => x"38",
          1760 => x"84",
          1761 => x"98",
          1762 => x"3d",
          1763 => x"51",
          1764 => x"86",
          1765 => x"c4",
          1766 => x"64",
          1767 => x"38",
          1768 => x"5c",
          1769 => x"db",
          1770 => x"ff",
          1771 => x"e0",
          1772 => x"b5",
          1773 => x"05",
          1774 => x"08",
          1775 => x"fe",
          1776 => x"eb",
          1777 => x"2e",
          1778 => x"ff",
          1779 => x"27",
          1780 => x"81",
          1781 => x"05",
          1782 => x"11",
          1783 => x"3f",
          1784 => x"fc",
          1785 => x"ff",
          1786 => x"e0",
          1787 => x"b5",
          1788 => x"05",
          1789 => x"08",
          1790 => x"84",
          1791 => x"79",
          1792 => x"7b",
          1793 => x"92",
          1794 => x"53",
          1795 => x"a3",
          1796 => x"44",
          1797 => x"3f",
          1798 => x"11",
          1799 => x"3f",
          1800 => x"82",
          1801 => x"89",
          1802 => x"cd",
          1803 => x"80",
          1804 => x"45",
          1805 => x"78",
          1806 => x"08",
          1807 => x"59",
          1808 => x"cc",
          1809 => x"33",
          1810 => x"de",
          1811 => x"e4",
          1812 => x"fe",
          1813 => x"e8",
          1814 => x"de",
          1815 => x"80",
          1816 => x"44",
          1817 => x"59",
          1818 => x"c0",
          1819 => x"33",
          1820 => x"de",
          1821 => x"ff",
          1822 => x"82",
          1823 => x"de",
          1824 => x"38",
          1825 => x"82",
          1826 => x"3d",
          1827 => x"51",
          1828 => x"80",
          1829 => x"7a",
          1830 => x"90",
          1831 => x"2a",
          1832 => x"78",
          1833 => x"83",
          1834 => x"ff",
          1835 => x"62",
          1836 => x"3f",
          1837 => x"b5",
          1838 => x"05",
          1839 => x"08",
          1840 => x"fe",
          1841 => x"e7",
          1842 => x"2e",
          1843 => x"05",
          1844 => x"b5",
          1845 => x"05",
          1846 => x"08",
          1847 => x"33",
          1848 => x"a0",
          1849 => x"80",
          1850 => x"3f",
          1851 => x"2e",
          1852 => x"38",
          1853 => x"84",
          1854 => x"98",
          1855 => x"02",
          1856 => x"81",
          1857 => x"d4",
          1858 => x"39",
          1859 => x"84",
          1860 => x"98",
          1861 => x"3d",
          1862 => x"51",
          1863 => x"80",
          1864 => x"c2",
          1865 => x"23",
          1866 => x"53",
          1867 => x"82",
          1868 => x"39",
          1869 => x"d8",
          1870 => x"f8",
          1871 => x"ff",
          1872 => x"59",
          1873 => x"9f",
          1874 => x"d0",
          1875 => x"ff",
          1876 => x"e0",
          1877 => x"59",
          1878 => x"82",
          1879 => x"39",
          1880 => x"3f",
          1881 => x"11",
          1882 => x"3f",
          1883 => x"e4",
          1884 => x"ff",
          1885 => x"e0",
          1886 => x"61",
          1887 => x"b5",
          1888 => x"05",
          1889 => x"08",
          1890 => x"08",
          1891 => x"9d",
          1892 => x"80",
          1893 => x"3f",
          1894 => x"2e",
          1895 => x"38",
          1896 => x"84",
          1897 => x"98",
          1898 => x"71",
          1899 => x"b5",
          1900 => x"b3",
          1901 => x"80",
          1902 => x"ab",
          1903 => x"f5",
          1904 => x"51",
          1905 => x"04",
          1906 => x"84",
          1907 => x"98",
          1908 => x"52",
          1909 => x"3f",
          1910 => x"08",
          1911 => x"98",
          1912 => x"9c",
          1913 => x"c8",
          1914 => x"99",
          1915 => x"51",
          1916 => x"a6",
          1917 => x"97",
          1918 => x"cc",
          1919 => x"f1",
          1920 => x"e0",
          1921 => x"82",
          1922 => x"84",
          1923 => x"98",
          1924 => x"80",
          1925 => x"08",
          1926 => x"08",
          1927 => x"7a",
          1928 => x"89",
          1929 => x"ca",
          1930 => x"c2",
          1931 => x"82",
          1932 => x"80",
          1933 => x"ff",
          1934 => x"b5",
          1935 => x"3f",
          1936 => x"54",
          1937 => x"3d",
          1938 => x"3f",
          1939 => x"c7",
          1940 => x"51",
          1941 => x"58",
          1942 => x"55",
          1943 => x"80",
          1944 => x"51",
          1945 => x"82",
          1946 => x"72",
          1947 => x"80",
          1948 => x"5a",
          1949 => x"8d",
          1950 => x"5c",
          1951 => x"32",
          1952 => x"38",
          1953 => x"38",
          1954 => x"3f",
          1955 => x"39",
          1956 => x"3f",
          1957 => x"0b",
          1958 => x"8c",
          1959 => x"52",
          1960 => x"98",
          1961 => x"87",
          1962 => x"3f",
          1963 => x"0c",
          1964 => x"55",
          1965 => x"e7",
          1966 => x"75",
          1967 => x"73",
          1968 => x"98",
          1969 => x"0b",
          1970 => x"83",
          1971 => x"82",
          1972 => x"02",
          1973 => x"82",
          1974 => x"13",
          1975 => x"0c",
          1976 => x"82",
          1977 => x"82",
          1978 => x"80",
          1979 => x"51",
          1980 => x"04",
          1981 => x"55",
          1982 => x"81",
          1983 => x"2e",
          1984 => x"53",
          1985 => x"2e",
          1986 => x"53",
          1987 => x"09",
          1988 => x"12",
          1989 => x"a2",
          1990 => x"2e",
          1991 => x"81",
          1992 => x"70",
          1993 => x"80",
          1994 => x"72",
          1995 => x"81",
          1996 => x"32",
          1997 => x"51",
          1998 => x"80",
          1999 => x"75",
          2000 => x"0c",
          2001 => x"76",
          2002 => x"86",
          2003 => x"b2",
          2004 => x"80",
          2005 => x"e0",
          2006 => x"3d",
          2007 => x"52",
          2008 => x"98",
          2009 => x"82",
          2010 => x"84",
          2011 => x"26",
          2012 => x"84",
          2013 => x"86",
          2014 => x"26",
          2015 => x"86",
          2016 => x"38",
          2017 => x"87",
          2018 => x"87",
          2019 => x"c0",
          2020 => x"c0",
          2021 => x"c0",
          2022 => x"c0",
          2023 => x"c0",
          2024 => x"c0",
          2025 => x"a4",
          2026 => x"80",
          2027 => x"52",
          2028 => x"0d",
          2029 => x"c0",
          2030 => x"c0",
          2031 => x"87",
          2032 => x"1c",
          2033 => x"79",
          2034 => x"08",
          2035 => x"98",
          2036 => x"87",
          2037 => x"1c",
          2038 => x"7b",
          2039 => x"08",
          2040 => x"0c",
          2041 => x"83",
          2042 => x"57",
          2043 => x"55",
          2044 => x"53",
          2045 => x"c8",
          2046 => x"3d",
          2047 => x"05",
          2048 => x"09",
          2049 => x"83",
          2050 => x"07",
          2051 => x"38",
          2052 => x"3f",
          2053 => x"98",
          2054 => x"81",
          2055 => x"2e",
          2056 => x"72",
          2057 => x"76",
          2058 => x"38",
          2059 => x"0d",
          2060 => x"54",
          2061 => x"8a",
          2062 => x"70",
          2063 => x"54",
          2064 => x"82",
          2065 => x"fb",
          2066 => x"de",
          2067 => x"55",
          2068 => x"80",
          2069 => x"51",
          2070 => x"06",
          2071 => x"38",
          2072 => x"51",
          2073 => x"81",
          2074 => x"38",
          2075 => x"51",
          2076 => x"06",
          2077 => x"80",
          2078 => x"52",
          2079 => x"0c",
          2080 => x"02",
          2081 => x"2a",
          2082 => x"34",
          2083 => x"02",
          2084 => x"09",
          2085 => x"51",
          2086 => x"81",
          2087 => x"84",
          2088 => x"c0",
          2089 => x"2a",
          2090 => x"80",
          2091 => x"81",
          2092 => x"81",
          2093 => x"80",
          2094 => x"81",
          2095 => x"75",
          2096 => x"80",
          2097 => x"c0",
          2098 => x"0b",
          2099 => x"04",
          2100 => x"33",
          2101 => x"70",
          2102 => x"ff",
          2103 => x"70",
          2104 => x"87",
          2105 => x"86",
          2106 => x"08",
          2107 => x"54",
          2108 => x"91",
          2109 => x"d7",
          2110 => x"51",
          2111 => x"93",
          2112 => x"ff",
          2113 => x"87",
          2114 => x"86",
          2115 => x"72",
          2116 => x"ff",
          2117 => x"38",
          2118 => x"0d",
          2119 => x"33",
          2120 => x"c0",
          2121 => x"38",
          2122 => x"70",
          2123 => x"51",
          2124 => x"ff",
          2125 => x"70",
          2126 => x"90",
          2127 => x"82",
          2128 => x"04",
          2129 => x"81",
          2130 => x"fe",
          2131 => x"81",
          2132 => x"84",
          2133 => x"c0",
          2134 => x"2a",
          2135 => x"52",
          2136 => x"ff",
          2137 => x"70",
          2138 => x"90",
          2139 => x"98",
          2140 => x"98",
          2141 => x"0d",
          2142 => x"2a",
          2143 => x"84",
          2144 => x"82",
          2145 => x"08",
          2146 => x"94",
          2147 => x"9e",
          2148 => x"c0",
          2149 => x"87",
          2150 => x"0c",
          2151 => x"cc",
          2152 => x"de",
          2153 => x"82",
          2154 => x"08",
          2155 => x"bc",
          2156 => x"9e",
          2157 => x"c0",
          2158 => x"87",
          2159 => x"de",
          2160 => x"82",
          2161 => x"08",
          2162 => x"8c",
          2163 => x"82",
          2164 => x"9e",
          2165 => x"51",
          2166 => x"81",
          2167 => x"0b",
          2168 => x"80",
          2169 => x"2e",
          2170 => x"fa",
          2171 => x"08",
          2172 => x"52",
          2173 => x"71",
          2174 => x"c0",
          2175 => x"06",
          2176 => x"38",
          2177 => x"80",
          2178 => x"a0",
          2179 => x"80",
          2180 => x"de",
          2181 => x"90",
          2182 => x"52",
          2183 => x"52",
          2184 => x"87",
          2185 => x"80",
          2186 => x"83",
          2187 => x"34",
          2188 => x"70",
          2189 => x"70",
          2190 => x"82",
          2191 => x"9e",
          2192 => x"51",
          2193 => x"81",
          2194 => x"0b",
          2195 => x"c0",
          2196 => x"2e",
          2197 => x"82",
          2198 => x"08",
          2199 => x"70",
          2200 => x"82",
          2201 => x"08",
          2202 => x"51",
          2203 => x"80",
          2204 => x"84",
          2205 => x"2e",
          2206 => x"85",
          2207 => x"83",
          2208 => x"51",
          2209 => x"87",
          2210 => x"51",
          2211 => x"81",
          2212 => x"c0",
          2213 => x"51",
          2214 => x"0d",
          2215 => x"51",
          2216 => x"33",
          2217 => x"c8",
          2218 => x"c8",
          2219 => x"de",
          2220 => x"38",
          2221 => x"08",
          2222 => x"ff",
          2223 => x"54",
          2224 => x"cc",
          2225 => x"52",
          2226 => x"3f",
          2227 => x"2e",
          2228 => x"de",
          2229 => x"94",
          2230 => x"fd",
          2231 => x"82",
          2232 => x"11",
          2233 => x"88",
          2234 => x"73",
          2235 => x"08",
          2236 => x"82",
          2237 => x"82",
          2238 => x"8e",
          2239 => x"c9",
          2240 => x"df",
          2241 => x"38",
          2242 => x"88",
          2243 => x"85",
          2244 => x"82",
          2245 => x"51",
          2246 => x"33",
          2247 => x"ca",
          2248 => x"de",
          2249 => x"38",
          2250 => x"3f",
          2251 => x"2e",
          2252 => x"a3",
          2253 => x"73",
          2254 => x"51",
          2255 => x"33",
          2256 => x"ca",
          2257 => x"cb",
          2258 => x"de",
          2259 => x"ff",
          2260 => x"52",
          2261 => x"3f",
          2262 => x"e0",
          2263 => x"88",
          2264 => x"e8",
          2265 => x"86",
          2266 => x"bd",
          2267 => x"f7",
          2268 => x"c0",
          2269 => x"e0",
          2270 => x"ff",
          2271 => x"54",
          2272 => x"f0",
          2273 => x"51",
          2274 => x"08",
          2275 => x"54",
          2276 => x"cc",
          2277 => x"de",
          2278 => x"38",
          2279 => x"c0",
          2280 => x"82",
          2281 => x"76",
          2282 => x"08",
          2283 => x"b0",
          2284 => x"87",
          2285 => x"92",
          2286 => x"26",
          2287 => x"cc",
          2288 => x"bc",
          2289 => x"97",
          2290 => x"82",
          2291 => x"d8",
          2292 => x"ff",
          2293 => x"71",
          2294 => x"c0",
          2295 => x"08",
          2296 => x"3d",
          2297 => x"79",
          2298 => x"13",
          2299 => x"51",
          2300 => x"33",
          2301 => x"82",
          2302 => x"05",
          2303 => x"52",
          2304 => x"38",
          2305 => x"85",
          2306 => x"02",
          2307 => x"55",
          2308 => x"82",
          2309 => x"a3",
          2310 => x"a0",
          2311 => x"fc",
          2312 => x"3f",
          2313 => x"34",
          2314 => x"77",
          2315 => x"34",
          2316 => x"7c",
          2317 => x"88",
          2318 => x"33",
          2319 => x"70",
          2320 => x"74",
          2321 => x"fd",
          2322 => x"29",
          2323 => x"54",
          2324 => x"e0",
          2325 => x"33",
          2326 => x"70",
          2327 => x"a7",
          2328 => x"ff",
          2329 => x"81",
          2330 => x"74",
          2331 => x"87",
          2332 => x"77",
          2333 => x"08",
          2334 => x"df",
          2335 => x"3d",
          2336 => x"75",
          2337 => x"e4",
          2338 => x"3f",
          2339 => x"e8",
          2340 => x"0d",
          2341 => x"08",
          2342 => x"51",
          2343 => x"14",
          2344 => x"e6",
          2345 => x"82",
          2346 => x"95",
          2347 => x"82",
          2348 => x"80",
          2349 => x"0d",
          2350 => x"52",
          2351 => x"e9",
          2352 => x"38",
          2353 => x"52",
          2354 => x"c1",
          2355 => x"ba",
          2356 => x"82",
          2357 => x"e0",
          2358 => x"98",
          2359 => x"80",
          2360 => x"17",
          2361 => x"c0",
          2362 => x"ff",
          2363 => x"3d",
          2364 => x"5a",
          2365 => x"82",
          2366 => x"3f",
          2367 => x"ff",
          2368 => x"80",
          2369 => x"81",
          2370 => x"80",
          2371 => x"9d",
          2372 => x"58",
          2373 => x"25",
          2374 => x"05",
          2375 => x"74",
          2376 => x"2a",
          2377 => x"38",
          2378 => x"08",
          2379 => x"89",
          2380 => x"89",
          2381 => x"a0",
          2382 => x"9b",
          2383 => x"ab",
          2384 => x"ab",
          2385 => x"74",
          2386 => x"0c",
          2387 => x"7c",
          2388 => x"59",
          2389 => x"06",
          2390 => x"77",
          2391 => x"5b",
          2392 => x"a0",
          2393 => x"75",
          2394 => x"29",
          2395 => x"55",
          2396 => x"08",
          2397 => x"a9",
          2398 => x"c5",
          2399 => x"2e",
          2400 => x"b5",
          2401 => x"1a",
          2402 => x"05",
          2403 => x"08",
          2404 => x"78",
          2405 => x"e0",
          2406 => x"85",
          2407 => x"70",
          2408 => x"27",
          2409 => x"e0",
          2410 => x"3d",
          2411 => x"b4",
          2412 => x"af",
          2413 => x"df",
          2414 => x"38",
          2415 => x"73",
          2416 => x"81",
          2417 => x"56",
          2418 => x"51",
          2419 => x"82",
          2420 => x"80",
          2421 => x"52",
          2422 => x"f3",
          2423 => x"8c",
          2424 => x"d3",
          2425 => x"08",
          2426 => x"f8",
          2427 => x"9a",
          2428 => x"82",
          2429 => x"06",
          2430 => x"51",
          2431 => x"08",
          2432 => x"25",
          2433 => x"05",
          2434 => x"80",
          2435 => x"51",
          2436 => x"ff",
          2437 => x"38",
          2438 => x"06",
          2439 => x"df",
          2440 => x"e4",
          2441 => x"3f",
          2442 => x"3f",
          2443 => x"98",
          2444 => x"38",
          2445 => x"33",
          2446 => x"f7",
          2447 => x"2c",
          2448 => x"82",
          2449 => x"33",
          2450 => x"59",
          2451 => x"80",
          2452 => x"74",
          2453 => x"05",
          2454 => x"24",
          2455 => x"77",
          2456 => x"08",
          2457 => x"d7",
          2458 => x"56",
          2459 => x"81",
          2460 => x"81",
          2461 => x"26",
          2462 => x"51",
          2463 => x"81",
          2464 => x"39",
          2465 => x"38",
          2466 => x"34",
          2467 => x"f7",
          2468 => x"2c",
          2469 => x"cd",
          2470 => x"57",
          2471 => x"81",
          2472 => x"14",
          2473 => x"d4",
          2474 => x"92",
          2475 => x"82",
          2476 => x"75",
          2477 => x"fd",
          2478 => x"e0",
          2479 => x"dc",
          2480 => x"38",
          2481 => x"27",
          2482 => x"2c",
          2483 => x"74",
          2484 => x"74",
          2485 => x"05",
          2486 => x"56",
          2487 => x"33",
          2488 => x"dc",
          2489 => x"74",
          2490 => x"7e",
          2491 => x"82",
          2492 => x"70",
          2493 => x"05",
          2494 => x"5a",
          2495 => x"38",
          2496 => x"70",
          2497 => x"74",
          2498 => x"05",
          2499 => x"56",
          2500 => x"82",
          2501 => x"98",
          2502 => x"56",
          2503 => x"82",
          2504 => x"97",
          2505 => x"81",
          2506 => x"f7",
          2507 => x"24",
          2508 => x"34",
          2509 => x"dc",
          2510 => x"f3",
          2511 => x"dc",
          2512 => x"73",
          2513 => x"d8",
          2514 => x"d8",
          2515 => x"dc",
          2516 => x"51",
          2517 => x"33",
          2518 => x"f7",
          2519 => x"74",
          2520 => x"14",
          2521 => x"52",
          2522 => x"74",
          2523 => x"05",
          2524 => x"58",
          2525 => x"82",
          2526 => x"95",
          2527 => x"98",
          2528 => x"33",
          2529 => x"fa",
          2530 => x"88",
          2531 => x"80",
          2532 => x"98",
          2533 => x"55",
          2534 => x"39",
          2535 => x"80",
          2536 => x"8a",
          2537 => x"d8",
          2538 => x"e0",
          2539 => x"96",
          2540 => x"80",
          2541 => x"79",
          2542 => x"7a",
          2543 => x"80",
          2544 => x"e0",
          2545 => x"f7",
          2546 => x"b8",
          2547 => x"51",
          2548 => x"33",
          2549 => x"34",
          2550 => x"82",
          2551 => x"55",
          2552 => x"ff",
          2553 => x"74",
          2554 => x"ff",
          2555 => x"ad",
          2556 => x"74",
          2557 => x"33",
          2558 => x"80",
          2559 => x"98",
          2560 => x"55",
          2561 => x"fc",
          2562 => x"3f",
          2563 => x"70",
          2564 => x"51",
          2565 => x"38",
          2566 => x"ff",
          2567 => x"29",
          2568 => x"82",
          2569 => x"75",
          2570 => x"f7",
          2571 => x"f7",
          2572 => x"27",
          2573 => x"52",
          2574 => x"34",
          2575 => x"92",
          2576 => x"81",
          2577 => x"56",
          2578 => x"b8",
          2579 => x"82",
          2580 => x"0b",
          2581 => x"f7",
          2582 => x"38",
          2583 => x"2e",
          2584 => x"3f",
          2585 => x"34",
          2586 => x"81",
          2587 => x"9c",
          2588 => x"7a",
          2589 => x"11",
          2590 => x"38",
          2591 => x"e0",
          2592 => x"e0",
          2593 => x"53",
          2594 => x"3f",
          2595 => x"08",
          2596 => x"74",
          2597 => x"7a",
          2598 => x"82",
          2599 => x"a4",
          2600 => x"82",
          2601 => x"82",
          2602 => x"05",
          2603 => x"bd",
          2604 => x"82",
          2605 => x"74",
          2606 => x"99",
          2607 => x"f7",
          2608 => x"ff",
          2609 => x"51",
          2610 => x"73",
          2611 => x"82",
          2612 => x"f7",
          2613 => x"79",
          2614 => x"82",
          2615 => x"82",
          2616 => x"77",
          2617 => x"08",
          2618 => x"dc",
          2619 => x"ff",
          2620 => x"f7",
          2621 => x"e0",
          2622 => x"51",
          2623 => x"33",
          2624 => x"34",
          2625 => x"fa",
          2626 => x"80",
          2627 => x"80",
          2628 => x"ff",
          2629 => x"54",
          2630 => x"76",
          2631 => x"54",
          2632 => x"34",
          2633 => x"15",
          2634 => x"88",
          2635 => x"fe",
          2636 => x"06",
          2637 => x"74",
          2638 => x"82",
          2639 => x"e0",
          2640 => x"55",
          2641 => x"34",
          2642 => x"73",
          2643 => x"38",
          2644 => x"83",
          2645 => x"82",
          2646 => x"f9",
          2647 => x"84",
          2648 => x"e0",
          2649 => x"74",
          2650 => x"12",
          2651 => x"05",
          2652 => x"06",
          2653 => x"59",
          2654 => x"71",
          2655 => x"e0",
          2656 => x"54",
          2657 => x"34",
          2658 => x"33",
          2659 => x"70",
          2660 => x"52",
          2661 => x"ff",
          2662 => x"71",
          2663 => x"53",
          2664 => x"08",
          2665 => x"17",
          2666 => x"0d",
          2667 => x"9e",
          2668 => x"86",
          2669 => x"2b",
          2670 => x"52",
          2671 => x"85",
          2672 => x"88",
          2673 => x"13",
          2674 => x"88",
          2675 => x"12",
          2676 => x"07",
          2677 => x"12",
          2678 => x"07",
          2679 => x"70",
          2680 => x"82",
          2681 => x"12",
          2682 => x"ff",
          2683 => x"53",
          2684 => x"14",
          2685 => x"0d",
          2686 => x"08",
          2687 => x"81",
          2688 => x"88",
          2689 => x"71",
          2690 => x"5f",
          2691 => x"54",
          2692 => x"51",
          2693 => x"70",
          2694 => x"8b",
          2695 => x"70",
          2696 => x"07",
          2697 => x"51",
          2698 => x"72",
          2699 => x"82",
          2700 => x"e0",
          2701 => x"12",
          2702 => x"07",
          2703 => x"33",
          2704 => x"70",
          2705 => x"57",
          2706 => x"71",
          2707 => x"fb",
          2708 => x"84",
          2709 => x"72",
          2710 => x"71",
          2711 => x"5b",
          2712 => x"33",
          2713 => x"02",
          2714 => x"70",
          2715 => x"71",
          2716 => x"e0",
          2717 => x"12",
          2718 => x"07",
          2719 => x"12",
          2720 => x"07",
          2721 => x"70",
          2722 => x"82",
          2723 => x"83",
          2724 => x"e0",
          2725 => x"04",
          2726 => x"08",
          2727 => x"06",
          2728 => x"82",
          2729 => x"11",
          2730 => x"8b",
          2731 => x"70",
          2732 => x"71",
          2733 => x"53",
          2734 => x"25",
          2735 => x"51",
          2736 => x"14",
          2737 => x"71",
          2738 => x"2a",
          2739 => x"14",
          2740 => x"87",
          2741 => x"19",
          2742 => x"88",
          2743 => x"5b",
          2744 => x"85",
          2745 => x"53",
          2746 => x"87",
          2747 => x"76",
          2748 => x"82",
          2749 => x"12",
          2750 => x"80",
          2751 => x"55",
          2752 => x"15",
          2753 => x"0d",
          2754 => x"38",
          2755 => x"38",
          2756 => x"0d",
          2757 => x"58",
          2758 => x"83",
          2759 => x"84",
          2760 => x"2b",
          2761 => x"81",
          2762 => x"cb",
          2763 => x"81",
          2764 => x"81",
          2765 => x"ff",
          2766 => x"51",
          2767 => x"38",
          2768 => x"5a",
          2769 => x"71",
          2770 => x"38",
          2771 => x"7a",
          2772 => x"82",
          2773 => x"12",
          2774 => x"ff",
          2775 => x"55",
          2776 => x"80",
          2777 => x"74",
          2778 => x"77",
          2779 => x"75",
          2780 => x"82",
          2781 => x"f7",
          2782 => x"1c",
          2783 => x"8b",
          2784 => x"5e",
          2785 => x"ff",
          2786 => x"56",
          2787 => x"ff",
          2788 => x"e0",
          2789 => x"72",
          2790 => x"71",
          2791 => x"5b",
          2792 => x"19",
          2793 => x"88",
          2794 => x"12",
          2795 => x"07",
          2796 => x"78",
          2797 => x"82",
          2798 => x"84",
          2799 => x"2b",
          2800 => x"52",
          2801 => x"85",
          2802 => x"84",
          2803 => x"8d",
          2804 => x"52",
          2805 => x"db",
          2806 => x"38",
          2807 => x"98",
          2808 => x"84",
          2809 => x"66",
          2810 => x"e0",
          2811 => x"84",
          2812 => x"7e",
          2813 => x"08",
          2814 => x"7b",
          2815 => x"ba",
          2816 => x"e0",
          2817 => x"e0",
          2818 => x"70",
          2819 => x"73",
          2820 => x"88",
          2821 => x"ff",
          2822 => x"73",
          2823 => x"33",
          2824 => x"53",
          2825 => x"54",
          2826 => x"80",
          2827 => x"06",
          2828 => x"42",
          2829 => x"71",
          2830 => x"70",
          2831 => x"71",
          2832 => x"56",
          2833 => x"75",
          2834 => x"54",
          2835 => x"18",
          2836 => x"8f",
          2837 => x"83",
          2838 => x"7f",
          2839 => x"78",
          2840 => x"7f",
          2841 => x"38",
          2842 => x"33",
          2843 => x"f4",
          2844 => x"b7",
          2845 => x"ff",
          2846 => x"2b",
          2847 => x"53",
          2848 => x"e0",
          2849 => x"ff",
          2850 => x"60",
          2851 => x"38",
          2852 => x"88",
          2853 => x"33",
          2854 => x"f4",
          2855 => x"df",
          2856 => x"ff",
          2857 => x"2b",
          2858 => x"53",
          2859 => x"e0",
          2860 => x"05",
          2861 => x"06",
          2862 => x"f9",
          2863 => x"82",
          2864 => x"7d",
          2865 => x"51",
          2866 => x"98",
          2867 => x"38",
          2868 => x"8f",
          2869 => x"88",
          2870 => x"3f",
          2871 => x"94",
          2872 => x"77",
          2873 => x"82",
          2874 => x"08",
          2875 => x"52",
          2876 => x"e1",
          2877 => x"3d",
          2878 => x"05",
          2879 => x"87",
          2880 => x"71",
          2881 => x"04",
          2882 => x"02",
          2883 => x"83",
          2884 => x"72",
          2885 => x"53",
          2886 => x"38",
          2887 => x"c0",
          2888 => x"85",
          2889 => x"52",
          2890 => x"70",
          2891 => x"8c",
          2892 => x"fc",
          2893 => x"87",
          2894 => x"2e",
          2895 => x"34",
          2896 => x"82",
          2897 => x"f3",
          2898 => x"05",
          2899 => x"83",
          2900 => x"e0",
          2901 => x"71",
          2902 => x"2b",
          2903 => x"92",
          2904 => x"41",
          2905 => x"87",
          2906 => x"84",
          2907 => x"70",
          2908 => x"2e",
          2909 => x"70",
          2910 => x"80",
          2911 => x"2e",
          2912 => x"26",
          2913 => x"87",
          2914 => x"38",
          2915 => x"80",
          2916 => x"99",
          2917 => x"8c",
          2918 => x"51",
          2919 => x"8d",
          2920 => x"81",
          2921 => x"2e",
          2922 => x"52",
          2923 => x"ed",
          2924 => x"71",
          2925 => x"53",
          2926 => x"0d",
          2927 => x"02",
          2928 => x"58",
          2929 => x"fc",
          2930 => x"06",
          2931 => x"81",
          2932 => x"2b",
          2933 => x"92",
          2934 => x"40",
          2935 => x"c0",
          2936 => x"76",
          2937 => x"2a",
          2938 => x"80",
          2939 => x"5c",
          2940 => x"81",
          2941 => x"80",
          2942 => x"08",
          2943 => x"8c",
          2944 => x"77",
          2945 => x"0c",
          2946 => x"08",
          2947 => x"38",
          2948 => x"70",
          2949 => x"5b",
          2950 => x"fc",
          2951 => x"7d",
          2952 => x"80",
          2953 => x"38",
          2954 => x"98",
          2955 => x"0d",
          2956 => x"02",
          2957 => x"54",
          2958 => x"98",
          2959 => x"80",
          2960 => x"8c",
          2961 => x"dc",
          2962 => x"84",
          2963 => x"54",
          2964 => x"39",
          2965 => x"cb",
          2966 => x"81",
          2967 => x"8a",
          2968 => x"71",
          2969 => x"52",
          2970 => x"c0",
          2971 => x"82",
          2972 => x"39",
          2973 => x"77",
          2974 => x"72",
          2975 => x"73",
          2976 => x"04",
          2977 => x"71",
          2978 => x"98",
          2979 => x"fd",
          2980 => x"12",
          2981 => x"07",
          2982 => x"2b",
          2983 => x"0c",
          2984 => x"3d",
          2985 => x"84",
          2986 => x"72",
          2987 => x"2a",
          2988 => x"04",
          2989 => x"70",
          2990 => x"88",
          2991 => x"54",
          2992 => x"70",
          2993 => x"51",
          2994 => x"fe",
          2995 => x"51",
          2996 => x"81",
          2997 => x"55",
          2998 => x"3d",
          2999 => x"76",
          3000 => x"05",
          3001 => x"38",
          3002 => x"78",
          3003 => x"81",
          3004 => x"56",
          3005 => x"52",
          3006 => x"71",
          3007 => x"98",
          3008 => x"0d",
          3009 => x"73",
          3010 => x"33",
          3011 => x"e0",
          3012 => x"0b",
          3013 => x"0d",
          3014 => x"52",
          3015 => x"3f",
          3016 => x"38",
          3017 => x"52",
          3018 => x"e0",
          3019 => x"72",
          3020 => x"72",
          3021 => x"3d",
          3022 => x"80",
          3023 => x"7a",
          3024 => x"16",
          3025 => x"17",
          3026 => x"e0",
          3027 => x"b7",
          3028 => x"34",
          3029 => x"31",
          3030 => x"77",
          3031 => x"74",
          3032 => x"81",
          3033 => x"16",
          3034 => x"81",
          3035 => x"3d",
          3036 => x"56",
          3037 => x"2e",
          3038 => x"82",
          3039 => x"08",
          3040 => x"16",
          3041 => x"3f",
          3042 => x"38",
          3043 => x"0c",
          3044 => x"0d",
          3045 => x"57",
          3046 => x"58",
          3047 => x"76",
          3048 => x"06",
          3049 => x"78",
          3050 => x"38",
          3051 => x"52",
          3052 => x"3f",
          3053 => x"51",
          3054 => x"d2",
          3055 => x"8a",
          3056 => x"51",
          3057 => x"84",
          3058 => x"17",
          3059 => x"c8",
          3060 => x"b4",
          3061 => x"81",
          3062 => x"84",
          3063 => x"17",
          3064 => x"98",
          3065 => x"77",
          3066 => x"04",
          3067 => x"12",
          3068 => x"56",
          3069 => x"22",
          3070 => x"57",
          3071 => x"3d",
          3072 => x"70",
          3073 => x"81",
          3074 => x"81",
          3075 => x"72",
          3076 => x"24",
          3077 => x"81",
          3078 => x"38",
          3079 => x"70",
          3080 => x"74",
          3081 => x"98",
          3082 => x"06",
          3083 => x"89",
          3084 => x"54",
          3085 => x"e0",
          3086 => x"ff",
          3087 => x"2b",
          3088 => x"2a",
          3089 => x"e2",
          3090 => x"da",
          3091 => x"05",
          3092 => x"e0",
          3093 => x"83",
          3094 => x"f8",
          3095 => x"ff",
          3096 => x"2a",
          3097 => x"fc",
          3098 => x"38",
          3099 => x"05",
          3100 => x"e0",
          3101 => x"39",
          3102 => x"89",
          3103 => x"7c",
          3104 => x"77",
          3105 => x"08",
          3106 => x"72",
          3107 => x"24",
          3108 => x"82",
          3109 => x"38",
          3110 => x"70",
          3111 => x"76",
          3112 => x"98",
          3113 => x"d9",
          3114 => x"05",
          3115 => x"54",
          3116 => x"77",
          3117 => x"8f",
          3118 => x"34",
          3119 => x"2a",
          3120 => x"fa",
          3121 => x"82",
          3122 => x"83",
          3123 => x"2a",
          3124 => x"2a",
          3125 => x"06",
          3126 => x"ec",
          3127 => x"05",
          3128 => x"e0",
          3129 => x"80",
          3130 => x"52",
          3131 => x"b8",
          3132 => x"76",
          3133 => x"75",
          3134 => x"08",
          3135 => x"77",
          3136 => x"fc",
          3137 => x"51",
          3138 => x"98",
          3139 => x"72",
          3140 => x"17",
          3141 => x"3d",
          3142 => x"7e",
          3143 => x"75",
          3144 => x"27",
          3145 => x"ff",
          3146 => x"3f",
          3147 => x"98",
          3148 => x"54",
          3149 => x"39",
          3150 => x"39",
          3151 => x"82",
          3152 => x"08",
          3153 => x"98",
          3154 => x"98",
          3155 => x"74",
          3156 => x"e0",
          3157 => x"fe",
          3158 => x"74",
          3159 => x"17",
          3160 => x"73",
          3161 => x"26",
          3162 => x"e0",
          3163 => x"3d",
          3164 => x"5b",
          3165 => x"77",
          3166 => x"78",
          3167 => x"79",
          3168 => x"55",
          3169 => x"e0",
          3170 => x"e0",
          3171 => x"9c",
          3172 => x"82",
          3173 => x"70",
          3174 => x"38",
          3175 => x"e2",
          3176 => x"76",
          3177 => x"7a",
          3178 => x"e0",
          3179 => x"86",
          3180 => x"e0",
          3181 => x"07",
          3182 => x"98",
          3183 => x"81",
          3184 => x"2e",
          3185 => x"74",
          3186 => x"27",
          3187 => x"80",
          3188 => x"9c",
          3189 => x"56",
          3190 => x"52",
          3191 => x"98",
          3192 => x"82",
          3193 => x"06",
          3194 => x"82",
          3195 => x"72",
          3196 => x"51",
          3197 => x"78",
          3198 => x"73",
          3199 => x"52",
          3200 => x"98",
          3201 => x"82",
          3202 => x"55",
          3203 => x"80",
          3204 => x"76",
          3205 => x"08",
          3206 => x"0c",
          3207 => x"08",
          3208 => x"ff",
          3209 => x"81",
          3210 => x"39",
          3211 => x"8c",
          3212 => x"98",
          3213 => x"55",
          3214 => x"0d",
          3215 => x"55",
          3216 => x"58",
          3217 => x"d8",
          3218 => x"3f",
          3219 => x"08",
          3220 => x"77",
          3221 => x"8a",
          3222 => x"56",
          3223 => x"97",
          3224 => x"52",
          3225 => x"82",
          3226 => x"8a",
          3227 => x"72",
          3228 => x"56",
          3229 => x"0d",
          3230 => x"08",
          3231 => x"26",
          3232 => x"72",
          3233 => x"88",
          3234 => x"33",
          3235 => x"16",
          3236 => x"2a",
          3237 => x"58",
          3238 => x"16",
          3239 => x"8a",
          3240 => x"72",
          3241 => x"51",
          3242 => x"54",
          3243 => x"38",
          3244 => x"8b",
          3245 => x"08",
          3246 => x"74",
          3247 => x"75",
          3248 => x"08",
          3249 => x"98",
          3250 => x"2e",
          3251 => x"39",
          3252 => x"74",
          3253 => x"18",
          3254 => x"0c",
          3255 => x"7a",
          3256 => x"59",
          3257 => x"86",
          3258 => x"14",
          3259 => x"81",
          3260 => x"77",
          3261 => x"0c",
          3262 => x"76",
          3263 => x"74",
          3264 => x"39",
          3265 => x"2a",
          3266 => x"52",
          3267 => x"98",
          3268 => x"e0",
          3269 => x"55",
          3270 => x"f4",
          3271 => x"08",
          3272 => x"77",
          3273 => x"39",
          3274 => x"86",
          3275 => x"55",
          3276 => x"c4",
          3277 => x"81",
          3278 => x"98",
          3279 => x"98",
          3280 => x"82",
          3281 => x"15",
          3282 => x"3f",
          3283 => x"76",
          3284 => x"9c",
          3285 => x"98",
          3286 => x"0d",
          3287 => x"80",
          3288 => x"e0",
          3289 => x"80",
          3290 => x"98",
          3291 => x"3f",
          3292 => x"98",
          3293 => x"08",
          3294 => x"58",
          3295 => x"83",
          3296 => x"55",
          3297 => x"07",
          3298 => x"16",
          3299 => x"88",
          3300 => x"56",
          3301 => x"82",
          3302 => x"08",
          3303 => x"2e",
          3304 => x"73",
          3305 => x"04",
          3306 => x"54",
          3307 => x"83",
          3308 => x"53",
          3309 => x"90",
          3310 => x"82",
          3311 => x"53",
          3312 => x"0d",
          3313 => x"83",
          3314 => x"55",
          3315 => x"51",
          3316 => x"8b",
          3317 => x"51",
          3318 => x"fd",
          3319 => x"53",
          3320 => x"05",
          3321 => x"05",
          3322 => x"51",
          3323 => x"e0",
          3324 => x"3d",
          3325 => x"08",
          3326 => x"98",
          3327 => x"98",
          3328 => x"3f",
          3329 => x"98",
          3330 => x"70",
          3331 => x"5b",
          3332 => x"06",
          3333 => x"86",
          3334 => x"73",
          3335 => x"38",
          3336 => x"73",
          3337 => x"81",
          3338 => x"38",
          3339 => x"54",
          3340 => x"83",
          3341 => x"38",
          3342 => x"8f",
          3343 => x"73",
          3344 => x"72",
          3345 => x"74",
          3346 => x"ac",
          3347 => x"2e",
          3348 => x"15",
          3349 => x"06",
          3350 => x"16",
          3351 => x"98",
          3352 => x"80",
          3353 => x"06",
          3354 => x"7b",
          3355 => x"75",
          3356 => x"98",
          3357 => x"80",
          3358 => x"80",
          3359 => x"53",
          3360 => x"39",
          3361 => x"06",
          3362 => x"27",
          3363 => x"70",
          3364 => x"2e",
          3365 => x"38",
          3366 => x"ff",
          3367 => x"84",
          3368 => x"39",
          3369 => x"3f",
          3370 => x"53",
          3371 => x"ac",
          3372 => x"51",
          3373 => x"5b",
          3374 => x"19",
          3375 => x"0b",
          3376 => x"0c",
          3377 => x"60",
          3378 => x"51",
          3379 => x"58",
          3380 => x"81",
          3381 => x"1a",
          3382 => x"ea",
          3383 => x"82",
          3384 => x"19",
          3385 => x"38",
          3386 => x"33",
          3387 => x"54",
          3388 => x"2e",
          3389 => x"81",
          3390 => x"38",
          3391 => x"09",
          3392 => x"33",
          3393 => x"55",
          3394 => x"2a",
          3395 => x"2e",
          3396 => x"bf",
          3397 => x"0c",
          3398 => x"81",
          3399 => x"56",
          3400 => x"ac",
          3401 => x"5d",
          3402 => x"83",
          3403 => x"38",
          3404 => x"f3",
          3405 => x"82",
          3406 => x"e5",
          3407 => x"ff",
          3408 => x"38",
          3409 => x"75",
          3410 => x"98",
          3411 => x"55",
          3412 => x"3f",
          3413 => x"81",
          3414 => x"39",
          3415 => x"06",
          3416 => x"27",
          3417 => x"2a",
          3418 => x"80",
          3419 => x"38",
          3420 => x"73",
          3421 => x"06",
          3422 => x"73",
          3423 => x"51",
          3424 => x"81",
          3425 => x"38",
          3426 => x"95",
          3427 => x"19",
          3428 => x"98",
          3429 => x"5c",
          3430 => x"78",
          3431 => x"08",
          3432 => x"fc",
          3433 => x"90",
          3434 => x"70",
          3435 => x"56",
          3436 => x"38",
          3437 => x"56",
          3438 => x"1d",
          3439 => x"5d",
          3440 => x"53",
          3441 => x"87",
          3442 => x"06",
          3443 => x"80",
          3444 => x"8c",
          3445 => x"7d",
          3446 => x"7b",
          3447 => x"22",
          3448 => x"73",
          3449 => x"ff",
          3450 => x"74",
          3451 => x"2a",
          3452 => x"56",
          3453 => x"75",
          3454 => x"57",
          3455 => x"75",
          3456 => x"57",
          3457 => x"b9",
          3458 => x"73",
          3459 => x"84",
          3460 => x"94",
          3461 => x"74",
          3462 => x"33",
          3463 => x"19",
          3464 => x"82",
          3465 => x"ff",
          3466 => x"81",
          3467 => x"27",
          3468 => x"54",
          3469 => x"05",
          3470 => x"a0",
          3471 => x"17",
          3472 => x"75",
          3473 => x"79",
          3474 => x"08",
          3475 => x"7b",
          3476 => x"80",
          3477 => x"98",
          3478 => x"2e",
          3479 => x"80",
          3480 => x"80",
          3481 => x"81",
          3482 => x"80",
          3483 => x"51",
          3484 => x"08",
          3485 => x"c5",
          3486 => x"e0",
          3487 => x"59",
          3488 => x"85",
          3489 => x"54",
          3490 => x"98",
          3491 => x"fa",
          3492 => x"82",
          3493 => x"98",
          3494 => x"3f",
          3495 => x"98",
          3496 => x"9c",
          3497 => x"57",
          3498 => x"8b",
          3499 => x"17",
          3500 => x"16",
          3501 => x"f3",
          3502 => x"ff",
          3503 => x"22",
          3504 => x"82",
          3505 => x"df",
          3506 => x"ff",
          3507 => x"d4",
          3508 => x"38",
          3509 => x"73",
          3510 => x"77",
          3511 => x"80",
          3512 => x"e0",
          3513 => x"80",
          3514 => x"d7",
          3515 => x"e2",
          3516 => x"82",
          3517 => x"82",
          3518 => x"51",
          3519 => x"52",
          3520 => x"9c",
          3521 => x"55",
          3522 => x"83",
          3523 => x"98",
          3524 => x"0d",
          3525 => x"13",
          3526 => x"2e",
          3527 => x"b1",
          3528 => x"e0",
          3529 => x"08",
          3530 => x"e0",
          3531 => x"ab",
          3532 => x"34",
          3533 => x"08",
          3534 => x"08",
          3535 => x"e0",
          3536 => x"80",
          3537 => x"81",
          3538 => x"e0",
          3539 => x"3d",
          3540 => x"5c",
          3541 => x"08",
          3542 => x"08",
          3543 => x"71",
          3544 => x"57",
          3545 => x"9d",
          3546 => x"1b",
          3547 => x"d0",
          3548 => x"51",
          3549 => x"74",
          3550 => x"11",
          3551 => x"83",
          3552 => x"51",
          3553 => x"08",
          3554 => x"75",
          3555 => x"38",
          3556 => x"74",
          3557 => x"74",
          3558 => x"25",
          3559 => x"73",
          3560 => x"39",
          3561 => x"57",
          3562 => x"11",
          3563 => x"f1",
          3564 => x"30",
          3565 => x"94",
          3566 => x"80",
          3567 => x"1c",
          3568 => x"56",
          3569 => x"85",
          3570 => x"e5",
          3571 => x"72",
          3572 => x"8b",
          3573 => x"38",
          3574 => x"81",
          3575 => x"58",
          3576 => x"ff",
          3577 => x"80",
          3578 => x"53",
          3579 => x"bf",
          3580 => x"e1",
          3581 => x"5a",
          3582 => x"96",
          3583 => x"ff",
          3584 => x"aa",
          3585 => x"51",
          3586 => x"84",
          3587 => x"53",
          3588 => x"8a",
          3589 => x"06",
          3590 => x"58",
          3591 => x"71",
          3592 => x"b5",
          3593 => x"0b",
          3594 => x"11",
          3595 => x"89",
          3596 => x"13",
          3597 => x"9c",
          3598 => x"e0",
          3599 => x"d9",
          3600 => x"19",
          3601 => x"82",
          3602 => x"3d",
          3603 => x"08",
          3604 => x"55",
          3605 => x"55",
          3606 => x"80",
          3607 => x"88",
          3608 => x"80",
          3609 => x"af",
          3610 => x"56",
          3611 => x"80",
          3612 => x"dc",
          3613 => x"33",
          3614 => x"ff",
          3615 => x"7d",
          3616 => x"08",
          3617 => x"08",
          3618 => x"92",
          3619 => x"82",
          3620 => x"38",
          3621 => x"08",
          3622 => x"e0",
          3623 => x"75",
          3624 => x"08",
          3625 => x"70",
          3626 => x"07",
          3627 => x"75",
          3628 => x"ff",
          3629 => x"c4",
          3630 => x"08",
          3631 => x"81",
          3632 => x"74",
          3633 => x"81",
          3634 => x"56",
          3635 => x"83",
          3636 => x"70",
          3637 => x"51",
          3638 => x"76",
          3639 => x"09",
          3640 => x"73",
          3641 => x"78",
          3642 => x"38",
          3643 => x"09",
          3644 => x"54",
          3645 => x"38",
          3646 => x"80",
          3647 => x"78",
          3648 => x"75",
          3649 => x"58",
          3650 => x"07",
          3651 => x"39",
          3652 => x"1a",
          3653 => x"71",
          3654 => x"2a",
          3655 => x"ae",
          3656 => x"19",
          3657 => x"11",
          3658 => x"38",
          3659 => x"07",
          3660 => x"70",
          3661 => x"73",
          3662 => x"81",
          3663 => x"55",
          3664 => x"8f",
          3665 => x"73",
          3666 => x"76",
          3667 => x"38",
          3668 => x"54",
          3669 => x"1a",
          3670 => x"80",
          3671 => x"55",
          3672 => x"eb",
          3673 => x"51",
          3674 => x"88",
          3675 => x"1f",
          3676 => x"94",
          3677 => x"ae",
          3678 => x"51",
          3679 => x"80",
          3680 => x"d1",
          3681 => x"26",
          3682 => x"70",
          3683 => x"7e",
          3684 => x"2e",
          3685 => x"38",
          3686 => x"07",
          3687 => x"78",
          3688 => x"81",
          3689 => x"80",
          3690 => x"07",
          3691 => x"ce",
          3692 => x"ff",
          3693 => x"06",
          3694 => x"38",
          3695 => x"11",
          3696 => x"a4",
          3697 => x"8a",
          3698 => x"fe",
          3699 => x"88",
          3700 => x"18",
          3701 => x"92",
          3702 => x"d4",
          3703 => x"2e",
          3704 => x"58",
          3705 => x"73",
          3706 => x"5c",
          3707 => x"8e",
          3708 => x"83",
          3709 => x"18",
          3710 => x"18",
          3711 => x"54",
          3712 => x"86",
          3713 => x"88",
          3714 => x"82",
          3715 => x"06",
          3716 => x"83",
          3717 => x"06",
          3718 => x"81",
          3719 => x"9f",
          3720 => x"2e",
          3721 => x"82",
          3722 => x"80",
          3723 => x"76",
          3724 => x"3f",
          3725 => x"56",
          3726 => x"be",
          3727 => x"09",
          3728 => x"2a",
          3729 => x"51",
          3730 => x"81",
          3731 => x"38",
          3732 => x"56",
          3733 => x"73",
          3734 => x"82",
          3735 => x"ac",
          3736 => x"70",
          3737 => x"2e",
          3738 => x"06",
          3739 => x"e4",
          3740 => x"1f",
          3741 => x"98",
          3742 => x"0d",
          3743 => x"73",
          3744 => x"2e",
          3745 => x"57",
          3746 => x"ba",
          3747 => x"ba",
          3748 => x"73",
          3749 => x"51",
          3750 => x"82",
          3751 => x"56",
          3752 => x"80",
          3753 => x"08",
          3754 => x"58",
          3755 => x"ff",
          3756 => x"26",
          3757 => x"06",
          3758 => x"99",
          3759 => x"ff",
          3760 => x"2a",
          3761 => x"06",
          3762 => x"30",
          3763 => x"07",
          3764 => x"54",
          3765 => x"81",
          3766 => x"25",
          3767 => x"24",
          3768 => x"78",
          3769 => x"51",
          3770 => x"0d",
          3771 => x"0b",
          3772 => x"0c",
          3773 => x"84",
          3774 => x"38",
          3775 => x"82",
          3776 => x"54",
          3777 => x"09",
          3778 => x"b8",
          3779 => x"2e",
          3780 => x"74",
          3781 => x"25",
          3782 => x"38",
          3783 => x"b5",
          3784 => x"80",
          3785 => x"e0",
          3786 => x"80",
          3787 => x"dc",
          3788 => x"3f",
          3789 => x"98",
          3790 => x"74",
          3791 => x"04",
          3792 => x"80",
          3793 => x"0c",
          3794 => x"98",
          3795 => x"e0",
          3796 => x"e0",
          3797 => x"05",
          3798 => x"80",
          3799 => x"76",
          3800 => x"72",
          3801 => x"51",
          3802 => x"81",
          3803 => x"72",
          3804 => x"38",
          3805 => x"53",
          3806 => x"f2",
          3807 => x"82",
          3808 => x"81",
          3809 => x"3f",
          3810 => x"70",
          3811 => x"86",
          3812 => x"74",
          3813 => x"8a",
          3814 => x"53",
          3815 => x"e0",
          3816 => x"82",
          3817 => x"9c",
          3818 => x"72",
          3819 => x"74",
          3820 => x"33",
          3821 => x"38",
          3822 => x"82",
          3823 => x"84",
          3824 => x"56",
          3825 => x"18",
          3826 => x"70",
          3827 => x"71",
          3828 => x"51",
          3829 => x"57",
          3830 => x"73",
          3831 => x"08",
          3832 => x"e0",
          3833 => x"2e",
          3834 => x"81",
          3835 => x"8c",
          3836 => x"83",
          3837 => x"84",
          3838 => x"81",
          3839 => x"51",
          3840 => x"83",
          3841 => x"2e",
          3842 => x"ce",
          3843 => x"98",
          3844 => x"8d",
          3845 => x"3f",
          3846 => x"15",
          3847 => x"34",
          3848 => x"81",
          3849 => x"72",
          3850 => x"ff",
          3851 => x"33",
          3852 => x"72",
          3853 => x"06",
          3854 => x"56",
          3855 => x"c9",
          3856 => x"82",
          3857 => x"8f",
          3858 => x"38",
          3859 => x"82",
          3860 => x"55",
          3861 => x"c8",
          3862 => x"80",
          3863 => x"e0",
          3864 => x"8d",
          3865 => x"88",
          3866 => x"05",
          3867 => x"38",
          3868 => x"51",
          3869 => x"08",
          3870 => x"82",
          3871 => x"ff",
          3872 => x"57",
          3873 => x"82",
          3874 => x"81",
          3875 => x"2e",
          3876 => x"16",
          3877 => x"70",
          3878 => x"0c",
          3879 => x"06",
          3880 => x"c0",
          3881 => x"ff",
          3882 => x"38",
          3883 => x"51",
          3884 => x"ac",
          3885 => x"39",
          3886 => x"38",
          3887 => x"53",
          3888 => x"15",
          3889 => x"51",
          3890 => x"8d",
          3891 => x"cc",
          3892 => x"0b",
          3893 => x"15",
          3894 => x"81",
          3895 => x"c8",
          3896 => x"ff",
          3897 => x"06",
          3898 => x"51",
          3899 => x"80",
          3900 => x"15",
          3901 => x"3f",
          3902 => x"06",
          3903 => x"81",
          3904 => x"c6",
          3905 => x"8b",
          3906 => x"b3",
          3907 => x"3f",
          3908 => x"e4",
          3909 => x"84",
          3910 => x"e0",
          3911 => x"14",
          3912 => x"08",
          3913 => x"f7",
          3914 => x"f7",
          3915 => x"f7",
          3916 => x"98",
          3917 => x"98",
          3918 => x"0d",
          3919 => x"ba",
          3920 => x"b2",
          3921 => x"aa",
          3922 => x"57",
          3923 => x"9a",
          3924 => x"ca",
          3925 => x"52",
          3926 => x"55",
          3927 => x"0c",
          3928 => x"3d",
          3929 => x"05",
          3930 => x"52",
          3931 => x"0b",
          3932 => x"82",
          3933 => x"e0",
          3934 => x"2e",
          3935 => x"73",
          3936 => x"78",
          3937 => x"92",
          3938 => x"84",
          3939 => x"98",
          3940 => x"88",
          3941 => x"02",
          3942 => x"59",
          3943 => x"38",
          3944 => x"cc",
          3945 => x"58",
          3946 => x"55",
          3947 => x"7a",
          3948 => x"56",
          3949 => x"55",
          3950 => x"80",
          3951 => x"57",
          3952 => x"77",
          3953 => x"ab",
          3954 => x"84",
          3955 => x"51",
          3956 => x"55",
          3957 => x"06",
          3958 => x"2a",
          3959 => x"2e",
          3960 => x"77",
          3961 => x"77",
          3962 => x"73",
          3963 => x"7a",
          3964 => x"08",
          3965 => x"8e",
          3966 => x"a0",
          3967 => x"52",
          3968 => x"62",
          3969 => x"54",
          3970 => x"2e",
          3971 => x"51",
          3972 => x"d0",
          3973 => x"98",
          3974 => x"ca",
          3975 => x"02",
          3976 => x"81",
          3977 => x"86",
          3978 => x"81",
          3979 => x"80",
          3980 => x"73",
          3981 => x"92",
          3982 => x"3f",
          3983 => x"90",
          3984 => x"08",
          3985 => x"81",
          3986 => x"38",
          3987 => x"11",
          3988 => x"0c",
          3989 => x"3f",
          3990 => x"08",
          3991 => x"5a",
          3992 => x"82",
          3993 => x"7a",
          3994 => x"23",
          3995 => x"1a",
          3996 => x"0b",
          3997 => x"81",
          3998 => x"8d",
          3999 => x"81",
          4000 => x"1a",
          4001 => x"7b",
          4002 => x"78",
          4003 => x"08",
          4004 => x"83",
          4005 => x"ff",
          4006 => x"55",
          4007 => x"76",
          4008 => x"27",
          4009 => x"5a",
          4010 => x"74",
          4011 => x"73",
          4012 => x"51",
          4013 => x"85",
          4014 => x"2a",
          4015 => x"0c",
          4016 => x"73",
          4017 => x"04",
          4018 => x"40",
          4019 => x"3d",
          4020 => x"3f",
          4021 => x"98",
          4022 => x"74",
          4023 => x"c7",
          4024 => x"87",
          4025 => x"95",
          4026 => x"56",
          4027 => x"34",
          4028 => x"08",
          4029 => x"27",
          4030 => x"82",
          4031 => x"ff",
          4032 => x"7e",
          4033 => x"2a",
          4034 => x"87",
          4035 => x"98",
          4036 => x"3f",
          4037 => x"27",
          4038 => x"a3",
          4039 => x"08",
          4040 => x"e0",
          4041 => x"82",
          4042 => x"59",
          4043 => x"77",
          4044 => x"55",
          4045 => x"31",
          4046 => x"81",
          4047 => x"82",
          4048 => x"83",
          4049 => x"a0",
          4050 => x"74",
          4051 => x"b8",
          4052 => x"89",
          4053 => x"3f",
          4054 => x"9c",
          4055 => x"06",
          4056 => x"76",
          4057 => x"08",
          4058 => x"e0",
          4059 => x"94",
          4060 => x"05",
          4061 => x"7b",
          4062 => x"76",
          4063 => x"0c",
          4064 => x"75",
          4065 => x"04",
          4066 => x"40",
          4067 => x"3d",
          4068 => x"3f",
          4069 => x"98",
          4070 => x"74",
          4071 => x"bf",
          4072 => x"70",
          4073 => x"74",
          4074 => x"82",
          4075 => x"9f",
          4076 => x"56",
          4077 => x"11",
          4078 => x"75",
          4079 => x"38",
          4080 => x"56",
          4081 => x"11",
          4082 => x"5c",
          4083 => x"88",
          4084 => x"52",
          4085 => x"51",
          4086 => x"55",
          4087 => x"b2",
          4088 => x"74",
          4089 => x"19",
          4090 => x"88",
          4091 => x"9c",
          4092 => x"38",
          4093 => x"e0",
          4094 => x"08",
          4095 => x"82",
          4096 => x"38",
          4097 => x"2a",
          4098 => x"38",
          4099 => x"5b",
          4100 => x"7b",
          4101 => x"52",
          4102 => x"3f",
          4103 => x"7e",
          4104 => x"74",
          4105 => x"b4",
          4106 => x"05",
          4107 => x"3f",
          4108 => x"78",
          4109 => x"18",
          4110 => x"7e",
          4111 => x"98",
          4112 => x"12",
          4113 => x"18",
          4114 => x"31",
          4115 => x"7b",
          4116 => x"ff",
          4117 => x"fd",
          4118 => x"18",
          4119 => x"51",
          4120 => x"0b",
          4121 => x"08",
          4122 => x"08",
          4123 => x"08",
          4124 => x"83",
          4125 => x"fd",
          4126 => x"07",
          4127 => x"75",
          4128 => x"04",
          4129 => x"05",
          4130 => x"82",
          4131 => x"08",
          4132 => x"86",
          4133 => x"73",
          4134 => x"08",
          4135 => x"82",
          4136 => x"08",
          4137 => x"11",
          4138 => x"16",
          4139 => x"75",
          4140 => x"08",
          4141 => x"3f",
          4142 => x"51",
          4143 => x"15",
          4144 => x"81",
          4145 => x"bb",
          4146 => x"17",
          4147 => x"90",
          4148 => x"8a",
          4149 => x"70",
          4150 => x"98",
          4151 => x"38",
          4152 => x"f1",
          4153 => x"82",
          4154 => x"98",
          4155 => x"0c",
          4156 => x"84",
          4157 => x"80",
          4158 => x"38",
          4159 => x"34",
          4160 => x"83",
          4161 => x"53",
          4162 => x"51",
          4163 => x"55",
          4164 => x"76",
          4165 => x"51",
          4166 => x"55",
          4167 => x"80",
          4168 => x"56",
          4169 => x"98",
          4170 => x"05",
          4171 => x"51",
          4172 => x"76",
          4173 => x"3f",
          4174 => x"8e",
          4175 => x"09",
          4176 => x"82",
          4177 => x"ff",
          4178 => x"80",
          4179 => x"34",
          4180 => x"05",
          4181 => x"3f",
          4182 => x"98",
          4183 => x"3d",
          4184 => x"d8",
          4185 => x"08",
          4186 => x"a0",
          4187 => x"c4",
          4188 => x"82",
          4189 => x"d9",
          4190 => x"ea",
          4191 => x"e0",
          4192 => x"3d",
          4193 => x"82",
          4194 => x"76",
          4195 => x"e0",
          4196 => x"82",
          4197 => x"b6",
          4198 => x"e0",
          4199 => x"08",
          4200 => x"82",
          4201 => x"52",
          4202 => x"98",
          4203 => x"2e",
          4204 => x"06",
          4205 => x"76",
          4206 => x"b8",
          4207 => x"76",
          4208 => x"51",
          4209 => x"38",
          4210 => x"81",
          4211 => x"f5",
          4212 => x"81",
          4213 => x"78",
          4214 => x"e1",
          4215 => x"58",
          4216 => x"75",
          4217 => x"08",
          4218 => x"f4",
          4219 => x"8d",
          4220 => x"11",
          4221 => x"82",
          4222 => x"d2",
          4223 => x"5c",
          4224 => x"38",
          4225 => x"55",
          4226 => x"73",
          4227 => x"76",
          4228 => x"33",
          4229 => x"15",
          4230 => x"05",
          4231 => x"06",
          4232 => x"e0",
          4233 => x"73",
          4234 => x"7a",
          4235 => x"76",
          4236 => x"0d",
          4237 => x"3d",
          4238 => x"eb",
          4239 => x"82",
          4240 => x"15",
          4241 => x"15",
          4242 => x"90",
          4243 => x"06",
          4244 => x"56",
          4245 => x"17",
          4246 => x"38",
          4247 => x"59",
          4248 => x"76",
          4249 => x"3f",
          4250 => x"54",
          4251 => x"3f",
          4252 => x"38",
          4253 => x"18",
          4254 => x"57",
          4255 => x"08",
          4256 => x"51",
          4257 => x"08",
          4258 => x"81",
          4259 => x"2e",
          4260 => x"88",
          4261 => x"80",
          4262 => x"80",
          4263 => x"08",
          4264 => x"70",
          4265 => x"5a",
          4266 => x"52",
          4267 => x"e0",
          4268 => x"95",
          4269 => x"39",
          4270 => x"3f",
          4271 => x"2e",
          4272 => x"79",
          4273 => x"38",
          4274 => x"94",
          4275 => x"83",
          4276 => x"38",
          4277 => x"3f",
          4278 => x"0b",
          4279 => x"39",
          4280 => x"bb",
          4281 => x"08",
          4282 => x"15",
          4283 => x"16",
          4284 => x"53",
          4285 => x"06",
          4286 => x"9c",
          4287 => x"16",
          4288 => x"0c",
          4289 => x"79",
          4290 => x"8b",
          4291 => x"52",
          4292 => x"3f",
          4293 => x"98",
          4294 => x"7a",
          4295 => x"e0",
          4296 => x"80",
          4297 => x"2b",
          4298 => x"86",
          4299 => x"06",
          4300 => x"38",
          4301 => x"e0",
          4302 => x"0c",
          4303 => x"23",
          4304 => x"3f",
          4305 => x"2e",
          4306 => x"86",
          4307 => x"76",
          4308 => x"0c",
          4309 => x"76",
          4310 => x"53",
          4311 => x"87",
          4312 => x"86",
          4313 => x"79",
          4314 => x"56",
          4315 => x"08",
          4316 => x"38",
          4317 => x"52",
          4318 => x"e0",
          4319 => x"e0",
          4320 => x"3f",
          4321 => x"98",
          4322 => x"38",
          4323 => x"08",
          4324 => x"f6",
          4325 => x"8c",
          4326 => x"70",
          4327 => x"82",
          4328 => x"54",
          4329 => x"0d",
          4330 => x"53",
          4331 => x"56",
          4332 => x"55",
          4333 => x"52",
          4334 => x"98",
          4335 => x"38",
          4336 => x"2b",
          4337 => x"86",
          4338 => x"38",
          4339 => x"74",
          4340 => x"04",
          4341 => x"80",
          4342 => x"3d",
          4343 => x"08",
          4344 => x"38",
          4345 => x"08",
          4346 => x"58",
          4347 => x"7c",
          4348 => x"ce",
          4349 => x"e0",
          4350 => x"81",
          4351 => x"82",
          4352 => x"f0",
          4353 => x"e0",
          4354 => x"e0",
          4355 => x"e0",
          4356 => x"08",
          4357 => x"7f",
          4358 => x"77",
          4359 => x"15",
          4360 => x"75",
          4361 => x"52",
          4362 => x"98",
          4363 => x"d6",
          4364 => x"1a",
          4365 => x"09",
          4366 => x"ff",
          4367 => x"83",
          4368 => x"25",
          4369 => x"9b",
          4370 => x"3f",
          4371 => x"70",
          4372 => x"59",
          4373 => x"7a",
          4374 => x"7c",
          4375 => x"11",
          4376 => x"15",
          4377 => x"3d",
          4378 => x"3d",
          4379 => x"95",
          4380 => x"e0",
          4381 => x"33",
          4382 => x"33",
          4383 => x"55",
          4384 => x"90",
          4385 => x"18",
          4386 => x"38",
          4387 => x"08",
          4388 => x"82",
          4389 => x"56",
          4390 => x"76",
          4391 => x"98",
          4392 => x"38",
          4393 => x"2e",
          4394 => x"a4",
          4395 => x"e0",
          4396 => x"38",
          4397 => x"08",
          4398 => x"82",
          4399 => x"8c",
          4400 => x"07",
          4401 => x"2e",
          4402 => x"55",
          4403 => x"0d",
          4404 => x"3d",
          4405 => x"d9",
          4406 => x"82",
          4407 => x"46",
          4408 => x"52",
          4409 => x"08",
          4410 => x"38",
          4411 => x"2a",
          4412 => x"55",
          4413 => x"54",
          4414 => x"80",
          4415 => x"54",
          4416 => x"52",
          4417 => x"e0",
          4418 => x"06",
          4419 => x"d6",
          4420 => x"98",
          4421 => x"5a",
          4422 => x"8a",
          4423 => x"3f",
          4424 => x"98",
          4425 => x"08",
          4426 => x"82",
          4427 => x"08",
          4428 => x"82",
          4429 => x"82",
          4430 => x"51",
          4431 => x"82",
          4432 => x"98",
          4433 => x"75",
          4434 => x"90",
          4435 => x"ff",
          4436 => x"55",
          4437 => x"f9",
          4438 => x"82",
          4439 => x"e8",
          4440 => x"bc",
          4441 => x"3f",
          4442 => x"98",
          4443 => x"52",
          4444 => x"3f",
          4445 => x"98",
          4446 => x"39",
          4447 => x"81",
          4448 => x"05",
          4449 => x"55",
          4450 => x"5a",
          4451 => x"ff",
          4452 => x"75",
          4453 => x"38",
          4454 => x"2e",
          4455 => x"82",
          4456 => x"06",
          4457 => x"73",
          4458 => x"52",
          4459 => x"e0",
          4460 => x"81",
          4461 => x"19",
          4462 => x"ae",
          4463 => x"0b",
          4464 => x"0a",
          4465 => x"d8",
          4466 => x"51",
          4467 => x"b8",
          4468 => x"a3",
          4469 => x"d9",
          4470 => x"11",
          4471 => x"54",
          4472 => x"ff",
          4473 => x"54",
          4474 => x"88",
          4475 => x"ff",
          4476 => x"78",
          4477 => x"90",
          4478 => x"0b",
          4479 => x"a9",
          4480 => x"39",
          4481 => x"ac",
          4482 => x"9a",
          4483 => x"3d",
          4484 => x"53",
          4485 => x"3d",
          4486 => x"08",
          4487 => x"38",
          4488 => x"3d",
          4489 => x"e0",
          4490 => x"82",
          4491 => x"81",
          4492 => x"af",
          4493 => x"aa",
          4494 => x"9f",
          4495 => x"70",
          4496 => x"3d",
          4497 => x"82",
          4498 => x"08",
          4499 => x"09",
          4500 => x"08",
          4501 => x"39",
          4502 => x"81",
          4503 => x"bd",
          4504 => x"82",
          4505 => x"56",
          4506 => x"52",
          4507 => x"02",
          4508 => x"16",
          4509 => x"51",
          4510 => x"07",
          4511 => x"81",
          4512 => x"70",
          4513 => x"55",
          4514 => x"64",
          4515 => x"51",
          4516 => x"08",
          4517 => x"82",
          4518 => x"80",
          4519 => x"78",
          4520 => x"98",
          4521 => x"55",
          4522 => x"81",
          4523 => x"81",
          4524 => x"76",
          4525 => x"81",
          4526 => x"e0",
          4527 => x"a5",
          4528 => x"e0",
          4529 => x"a3",
          4530 => x"74",
          4531 => x"04",
          4532 => x"33",
          4533 => x"57",
          4534 => x"52",
          4535 => x"e0",
          4536 => x"80",
          4537 => x"3d",
          4538 => x"e0",
          4539 => x"b8",
          4540 => x"a0",
          4541 => x"75",
          4542 => x"33",
          4543 => x"57",
          4544 => x"54",
          4545 => x"ff",
          4546 => x"55",
          4547 => x"0d",
          4548 => x"53",
          4549 => x"51",
          4550 => x"55",
          4551 => x"76",
          4552 => x"51",
          4553 => x"55",
          4554 => x"80",
          4555 => x"86",
          4556 => x"86",
          4557 => x"54",
          4558 => x"76",
          4559 => x"51",
          4560 => x"08",
          4561 => x"3d",
          4562 => x"5c",
          4563 => x"52",
          4564 => x"e0",
          4565 => x"70",
          4566 => x"51",
          4567 => x"38",
          4568 => x"80",
          4569 => x"5f",
          4570 => x"ff",
          4571 => x"57",
          4572 => x"74",
          4573 => x"82",
          4574 => x"08",
          4575 => x"e0",
          4576 => x"18",
          4577 => x"74",
          4578 => x"78",
          4579 => x"54",
          4580 => x"38",
          4581 => x"55",
          4582 => x"39",
          4583 => x"38",
          4584 => x"70",
          4585 => x"80",
          4586 => x"bc",
          4587 => x"ff",
          4588 => x"57",
          4589 => x"70",
          4590 => x"83",
          4591 => x"84",
          4592 => x"b8",
          4593 => x"e0",
          4594 => x"98",
          4595 => x"0d",
          4596 => x"52",
          4597 => x"e0",
          4598 => x"54",
          4599 => x"8b",
          4600 => x"58",
          4601 => x"33",
          4602 => x"86",
          4603 => x"9c",
          4604 => x"ff",
          4605 => x"98",
          4606 => x"52",
          4607 => x"3f",
          4608 => x"06",
          4609 => x"52",
          4610 => x"3f",
          4611 => x"ff",
          4612 => x"88",
          4613 => x"38",
          4614 => x"75",
          4615 => x"73",
          4616 => x"16",
          4617 => x"34",
          4618 => x"56",
          4619 => x"3d",
          4620 => x"2e",
          4621 => x"38",
          4622 => x"33",
          4623 => x"06",
          4624 => x"38",
          4625 => x"3d",
          4626 => x"82",
          4627 => x"08",
          4628 => x"ff",
          4629 => x"54",
          4630 => x"80",
          4631 => x"80",
          4632 => x"2e",
          4633 => x"54",
          4634 => x"52",
          4635 => x"e0",
          4636 => x"b1",
          4637 => x"52",
          4638 => x"54",
          4639 => x"77",
          4640 => x"78",
          4641 => x"51",
          4642 => x"08",
          4643 => x"0c",
          4644 => x"60",
          4645 => x"33",
          4646 => x"40",
          4647 => x"98",
          4648 => x"bd",
          4649 => x"b5",
          4650 => x"1a",
          4651 => x"33",
          4652 => x"55",
          4653 => x"97",
          4654 => x"58",
          4655 => x"70",
          4656 => x"56",
          4657 => x"7d",
          4658 => x"2a",
          4659 => x"08",
          4660 => x"77",
          4661 => x"26",
          4662 => x"59",
          4663 => x"9c",
          4664 => x"9c",
          4665 => x"55",
          4666 => x"99",
          4667 => x"ff",
          4668 => x"38",
          4669 => x"81",
          4670 => x"80",
          4671 => x"ff",
          4672 => x"7d",
          4673 => x"55",
          4674 => x"56",
          4675 => x"38",
          4676 => x"51",
          4677 => x"08",
          4678 => x"38",
          4679 => x"5c",
          4680 => x"5c",
          4681 => x"80",
          4682 => x"7c",
          4683 => x"c0",
          4684 => x"15",
          4685 => x"54",
          4686 => x"31",
          4687 => x"07",
          4688 => x"73",
          4689 => x"04",
          4690 => x"05",
          4691 => x"45",
          4692 => x"80",
          4693 => x"a0",
          4694 => x"82",
          4695 => x"74",
          4696 => x"82",
          4697 => x"05",
          4698 => x"8d",
          4699 => x"7f",
          4700 => x"98",
          4701 => x"56",
          4702 => x"76",
          4703 => x"8a",
          4704 => x"fc",
          4705 => x"92",
          4706 => x"38",
          4707 => x"74",
          4708 => x"15",
          4709 => x"38",
          4710 => x"84",
          4711 => x"80",
          4712 => x"06",
          4713 => x"56",
          4714 => x"89",
          4715 => x"43",
          4716 => x"30",
          4717 => x"91",
          4718 => x"2e",
          4719 => x"7a",
          4720 => x"81",
          4721 => x"38",
          4722 => x"3f",
          4723 => x"06",
          4724 => x"2e",
          4725 => x"90",
          4726 => x"57",
          4727 => x"b6",
          4728 => x"e0",
          4729 => x"ff",
          4730 => x"48",
          4731 => x"81",
          4732 => x"81",
          4733 => x"38",
          4734 => x"e0",
          4735 => x"38",
          4736 => x"75",
          4737 => x"48",
          4738 => x"b8",
          4739 => x"8a",
          4740 => x"06",
          4741 => x"62",
          4742 => x"8d",
          4743 => x"2e",
          4744 => x"93",
          4745 => x"80",
          4746 => x"81",
          4747 => x"67",
          4748 => x"dc",
          4749 => x"38",
          4750 => x"dc",
          4751 => x"57",
          4752 => x"76",
          4753 => x"51",
          4754 => x"08",
          4755 => x"2a",
          4756 => x"e0",
          4757 => x"46",
          4758 => x"ec",
          4759 => x"67",
          4760 => x"cc",
          4761 => x"38",
          4762 => x"cc",
          4763 => x"57",
          4764 => x"76",
          4765 => x"51",
          4766 => x"08",
          4767 => x"08",
          4768 => x"82",
          4769 => x"08",
          4770 => x"59",
          4771 => x"5d",
          4772 => x"11",
          4773 => x"71",
          4774 => x"52",
          4775 => x"09",
          4776 => x"18",
          4777 => x"79",
          4778 => x"58",
          4779 => x"38",
          4780 => x"70",
          4781 => x"3f",
          4782 => x"2e",
          4783 => x"98",
          4784 => x"38",
          4785 => x"59",
          4786 => x"7d",
          4787 => x"38",
          4788 => x"08",
          4789 => x"1a",
          4790 => x"74",
          4791 => x"55",
          4792 => x"fd",
          4793 => x"f5",
          4794 => x"79",
          4795 => x"f1",
          4796 => x"81",
          4797 => x"55",
          4798 => x"81",
          4799 => x"38",
          4800 => x"ff",
          4801 => x"e4",
          4802 => x"84",
          4803 => x"aa",
          4804 => x"ff",
          4805 => x"8e",
          4806 => x"7d",
          4807 => x"84",
          4808 => x"51",
          4809 => x"83",
          4810 => x"ff",
          4811 => x"8d",
          4812 => x"1b",
          4813 => x"95",
          4814 => x"ff",
          4815 => x"1b",
          4816 => x"9c",
          4817 => x"83",
          4818 => x"82",
          4819 => x"51",
          4820 => x"1b",
          4821 => x"ac",
          4822 => x"52",
          4823 => x"86",
          4824 => x"3f",
          4825 => x"a9",
          4826 => x"82",
          4827 => x"ae",
          4828 => x"1b",
          4829 => x"ff",
          4830 => x"8c",
          4831 => x"34",
          4832 => x"82",
          4833 => x"8d",
          4834 => x"fe",
          4835 => x"3f",
          4836 => x"51",
          4837 => x"e0",
          4838 => x"2e",
          4839 => x"54",
          4840 => x"ff",
          4841 => x"52",
          4842 => x"8b",
          4843 => x"8c",
          4844 => x"52",
          4845 => x"3f",
          4846 => x"ff",
          4847 => x"1b",
          4848 => x"d5",
          4849 => x"75",
          4850 => x"51",
          4851 => x"1f",
          4852 => x"d1",
          4853 => x"ff",
          4854 => x"7d",
          4855 => x"f8",
          4856 => x"ff",
          4857 => x"3f",
          4858 => x"39",
          4859 => x"2e",
          4860 => x"51",
          4861 => x"57",
          4862 => x"76",
          4863 => x"ff",
          4864 => x"82",
          4865 => x"98",
          4866 => x"3f",
          4867 => x"74",
          4868 => x"2e",
          4869 => x"2e",
          4870 => x"62",
          4871 => x"75",
          4872 => x"b1",
          4873 => x"38",
          4874 => x"74",
          4875 => x"93",
          4876 => x"26",
          4877 => x"83",
          4878 => x"38",
          4879 => x"51",
          4880 => x"e0",
          4881 => x"29",
          4882 => x"75",
          4883 => x"52",
          4884 => x"81",
          4885 => x"77",
          4886 => x"52",
          4887 => x"d4",
          4888 => x"3f",
          4889 => x"81",
          4890 => x"16",
          4891 => x"16",
          4892 => x"52",
          4893 => x"0b",
          4894 => x"82",
          4895 => x"34",
          4896 => x"7e",
          4897 => x"d8",
          4898 => x"ff",
          4899 => x"7a",
          4900 => x"81",
          4901 => x"80",
          4902 => x"a5",
          4903 => x"90",
          4904 => x"81",
          4905 => x"56",
          4906 => x"0d",
          4907 => x"59",
          4908 => x"57",
          4909 => x"f8",
          4910 => x"52",
          4911 => x"2e",
          4912 => x"33",
          4913 => x"76",
          4914 => x"57",
          4915 => x"38",
          4916 => x"38",
          4917 => x"8d",
          4918 => x"02",
          4919 => x"77",
          4920 => x"8d",
          4921 => x"08",
          4922 => x"17",
          4923 => x"77",
          4924 => x"25",
          4925 => x"75",
          4926 => x"ca",
          4927 => x"70",
          4928 => x"51",
          4929 => x"19",
          4930 => x"f9",
          4931 => x"56",
          4932 => x"fc",
          4933 => x"75",
          4934 => x"98",
          4935 => x"2e",
          4936 => x"08",
          4937 => x"e0",
          4938 => x"3d",
          4939 => x"52",
          4940 => x"74",
          4941 => x"0d",
          4942 => x"86",
          4943 => x"73",
          4944 => x"51",
          4945 => x"fd",
          4946 => x"05",
          4947 => x"ff",
          4948 => x"06",
          4949 => x"73",
          4950 => x"81",
          4951 => x"38",
          4952 => x"2e",
          4953 => x"ff",
          4954 => x"8d",
          4955 => x"70",
          4956 => x"12",
          4957 => x"82",
          4958 => x"fe",
          4959 => x"84",
          4960 => x"53",
          4961 => x"53",
          4962 => x"81",
          4963 => x"8b",
          4964 => x"70",
          4965 => x"0c",
          4966 => x"77",
          4967 => x"a7",
          4968 => x"d5",
          4969 => x"85",
          4970 => x"82",
          4971 => x"25",
          4972 => x"70",
          4973 => x"57",
          4974 => x"06",
          4975 => x"71",
          4976 => x"80",
          4977 => x"b8",
          4978 => x"31",
          4979 => x"51",
          4980 => x"06",
          4981 => x"f0",
          4982 => x"9a",
          4983 => x"12",
          4984 => x"39",
          4985 => x"a0",
          4986 => x"52",
          4987 => x"10",
          4988 => x"70",
          4989 => x"04",
          4990 => x"ff",
          4991 => x"00",
          4992 => x"85",
          4993 => x"93",
          4994 => x"a1",
          4995 => x"af",
          4996 => x"bd",
          4997 => x"cb",
          4998 => x"d7",
          4999 => x"e3",
          5000 => x"ef",
          5001 => x"fb",
          5002 => x"87",
          5003 => x"93",
          5004 => x"79",
          5005 => x"8a",
          5006 => x"61",
          5007 => x"52",
          5008 => x"95",
          5009 => x"b1",
          5010 => x"4c",
          5011 => x"b3",
          5012 => x"4c",
          5013 => x"b1",
          5014 => x"b3",
          5015 => x"91",
          5016 => x"ab",
          5017 => x"b5",
          5018 => x"bf",
          5019 => x"ca",
          5020 => x"4e",
          5021 => x"94",
          5022 => x"4e",
          5023 => x"4e",
          5024 => x"4e",
          5025 => x"51",
          5026 => x"7c",
          5027 => x"4e",
          5028 => x"4e",
          5029 => x"4e",
          5030 => x"4e",
          5031 => x"4e",
          5032 => x"4e",
          5033 => x"4e",
          5034 => x"4e",
          5035 => x"4e",
          5036 => x"4e",
          5037 => x"4e",
          5038 => x"4e",
          5039 => x"4e",
          5040 => x"4e",
          5041 => x"4e",
          5042 => x"4e",
          5043 => x"4e",
          5044 => x"4e",
          5045 => x"dc",
          5046 => x"4e",
          5047 => x"4e",
          5048 => x"4e",
          5049 => x"4e",
          5050 => x"4e",
          5051 => x"4e",
          5052 => x"4e",
          5053 => x"0c",
          5054 => x"e3",
          5055 => x"e3",
          5056 => x"73",
          5057 => x"4e",
          5058 => x"4e",
          5059 => x"20",
          5060 => x"4e",
          5061 => x"45",
          5062 => x"53",
          5063 => x"4e",
          5064 => x"69",
          5065 => x"63",
          5066 => x"69",
          5067 => x"61",
          5068 => x"65",
          5069 => x"65",
          5070 => x"70",
          5071 => x"66",
          5072 => x"6d",
          5073 => x"00",
          5074 => x"00",
          5075 => x"00",
          5076 => x"00",
          5077 => x"00",
          5078 => x"74",
          5079 => x"65",
          5080 => x"6f",
          5081 => x"73",
          5082 => x"73",
          5083 => x"6f",
          5084 => x"00",
          5085 => x"72",
          5086 => x"65",
          5087 => x"72",
          5088 => x"6b",
          5089 => x"61",
          5090 => x"66",
          5091 => x"6e",
          5092 => x"70",
          5093 => x"6e",
          5094 => x"61",
          5095 => x"65",
          5096 => x"00",
          5097 => x"64",
          5098 => x"00",
          5099 => x"72",
          5100 => x"69",
          5101 => x"00",
          5102 => x"6e",
          5103 => x"61",
          5104 => x"00",
          5105 => x"72",
          5106 => x"74",
          5107 => x"00",
          5108 => x"75",
          5109 => x"20",
          5110 => x"2e",
          5111 => x"6b",
          5112 => x"61",
          5113 => x"00",
          5114 => x"61",
          5115 => x"69",
          5116 => x"6d",
          5117 => x"6f",
          5118 => x"00",
          5119 => x"61",
          5120 => x"00",
          5121 => x"2c",
          5122 => x"69",
          5123 => x"65",
          5124 => x"00",
          5125 => x"20",
          5126 => x"00",
          5127 => x"63",
          5128 => x"6d",
          5129 => x"00",
          5130 => x"79",
          5131 => x"69",
          5132 => x"00",
          5133 => x"65",
          5134 => x"72",
          5135 => x"00",
          5136 => x"2e",
          5137 => x"6e",
          5138 => x"6f",
          5139 => x"75",
          5140 => x"25",
          5141 => x"75",
          5142 => x"73",
          5143 => x"00",
          5144 => x"00",
          5145 => x"00",
          5146 => x"58",
          5147 => x"20",
          5148 => x"00",
          5149 => x"00",
          5150 => x"00",
          5151 => x"00",
          5152 => x"00",
          5153 => x"30",
          5154 => x"31",
          5155 => x"55",
          5156 => x"30",
          5157 => x"25",
          5158 => x"00",
          5159 => x"65",
          5160 => x"61",
          5161 => x"00",
          5162 => x"6e",
          5163 => x"00",
          5164 => x"65",
          5165 => x"00",
          5166 => x"44",
          5167 => x"75",
          5168 => x"54",
          5169 => x"74",
          5170 => x"00",
          5171 => x"58",
          5172 => x"75",
          5173 => x"54",
          5174 => x"74",
          5175 => x"00",
          5176 => x"58",
          5177 => x"75",
          5178 => x"54",
          5179 => x"74",
          5180 => x"00",
          5181 => x"20",
          5182 => x"72",
          5183 => x"62",
          5184 => x"6d",
          5185 => x"00",
          5186 => x"63",
          5187 => x"00",
          5188 => x"2e",
          5189 => x"00",
          5190 => x"74",
          5191 => x"61",
          5192 => x"20",
          5193 => x"20",
          5194 => x"69",
          5195 => x"75",
          5196 => x"00",
          5197 => x"61",
          5198 => x"2e",
          5199 => x"79",
          5200 => x"00",
          5201 => x"6e",
          5202 => x"00",
          5203 => x"30",
          5204 => x"38",
          5205 => x"29",
          5206 => x"70",
          5207 => x"00",
          5208 => x"74",
          5209 => x"6c",
          5210 => x"00",
          5211 => x"6c",
          5212 => x"00",
          5213 => x"30",
          5214 => x"00",
          5215 => x"6e",
          5216 => x"40",
          5217 => x"2e",
          5218 => x"6c",
          5219 => x"65",
          5220 => x"78",
          5221 => x"00",
          5222 => x"74",
          5223 => x"6f",
          5224 => x"2e",
          5225 => x"74",
          5226 => x"61",
          5227 => x"69",
          5228 => x"00",
          5229 => x"62",
          5230 => x"2e",
          5231 => x"00",
          5232 => x"5c",
          5233 => x"73",
          5234 => x"5c",
          5235 => x"00",
          5236 => x"00",
          5237 => x"6d",
          5238 => x"00",
          5239 => x"65",
          5240 => x"64",
          5241 => x"74",
          5242 => x"73",
          5243 => x"64",
          5244 => x"6e",
          5245 => x"00",
          5246 => x"67",
          5247 => x"75",
          5248 => x"00",
          5249 => x"64",
          5250 => x"25",
          5251 => x"00",
          5252 => x"66",
          5253 => x"6f",
          5254 => x"72",
          5255 => x"63",
          5256 => x"00",
          5257 => x"65",
          5258 => x"6d",
          5259 => x"00",
          5260 => x"53",
          5261 => x"25",
          5262 => x"58",
          5263 => x"20",
          5264 => x"20",
          5265 => x"3a",
          5266 => x"00",
          5267 => x"4e",
          5268 => x"25",
          5269 => x"58",
          5270 => x"20",
          5271 => x"20",
          5272 => x"3a",
          5273 => x"00",
          5274 => x"20",
          5275 => x"25",
          5276 => x"58",
          5277 => x"20",
          5278 => x"20",
          5279 => x"63",
          5280 => x"64",
          5281 => x"20",
          5282 => x"20",
          5283 => x"72",
          5284 => x"64",
          5285 => x"20",
          5286 => x"52",
          5287 => x"6e",
          5288 => x"64",
          5289 => x"20",
          5290 => x"45",
          5291 => x"00",
          5292 => x"49",
          5293 => x"20",
          5294 => x"00",
          5295 => x"00",
          5296 => x"00",
          5297 => x"65",
          5298 => x"20",
          5299 => x"65",
          5300 => x"72",
          5301 => x"73",
          5302 => x"0a",
          5303 => x"20",
          5304 => x"6f",
          5305 => x"74",
          5306 => x"73",
          5307 => x"0a",
          5308 => x"20",
          5309 => x"74",
          5310 => x"72",
          5311 => x"20",
          5312 => x"0a",
          5313 => x"63",
          5314 => x"20",
          5315 => x"20",
          5316 => x"20",
          5317 => x"20",
          5318 => x"0a",
          5319 => x"20",
          5320 => x"43",
          5321 => x"65",
          5322 => x"20",
          5323 => x"30",
          5324 => x"00",
          5325 => x"41",
          5326 => x"20",
          5327 => x"20",
          5328 => x"25",
          5329 => x"48",
          5330 => x"20",
          5331 => x"65",
          5332 => x"43",
          5333 => x"65",
          5334 => x"30",
          5335 => x"00",
          5336 => x"00",
          5337 => x"00",
          5338 => x"00",
          5339 => x"6d",
          5340 => x"6e",
          5341 => x"44",
          5342 => x"02",
          5343 => x"00",
          5344 => x"3c",
          5345 => x"04",
          5346 => x"00",
          5347 => x"34",
          5348 => x"06",
          5349 => x"00",
          5350 => x"2c",
          5351 => x"01",
          5352 => x"00",
          5353 => x"24",
          5354 => x"0b",
          5355 => x"00",
          5356 => x"1c",
          5357 => x"0a",
          5358 => x"00",
          5359 => x"14",
          5360 => x"0c",
          5361 => x"00",
          5362 => x"0c",
          5363 => x"0f",
          5364 => x"00",
          5365 => x"04",
          5366 => x"10",
          5367 => x"00",
          5368 => x"fc",
          5369 => x"12",
          5370 => x"00",
          5371 => x"f4",
          5372 => x"14",
          5373 => x"00",
          5374 => x"00",
          5375 => x"00",
          5376 => x"7e",
          5377 => x"7e",
          5378 => x"7e",
          5379 => x"7e",
          5380 => x"00",
          5381 => x"00",
          5382 => x"00",
          5383 => x"00",
          5384 => x"00",
          5385 => x"74",
          5386 => x"74",
          5387 => x"00",
          5388 => x"25",
          5389 => x"6c",
          5390 => x"65",
          5391 => x"20",
          5392 => x"20",
          5393 => x"20",
          5394 => x"00",
          5395 => x"6f",
          5396 => x"61",
          5397 => x"6f",
          5398 => x"2c",
          5399 => x"69",
          5400 => x"00",
          5401 => x"7f",
          5402 => x"3d",
          5403 => x"00",
          5404 => x"00",
          5405 => x"53",
          5406 => x"4e",
          5407 => x"46",
          5408 => x"00",
          5409 => x"20",
          5410 => x"20",
          5411 => x"c0",
          5412 => x"00",
          5413 => x"07",
          5414 => x"1c",
          5415 => x"41",
          5416 => x"49",
          5417 => x"4f",
          5418 => x"9b",
          5419 => x"55",
          5420 => x"ab",
          5421 => x"b3",
          5422 => x"bb",
          5423 => x"c3",
          5424 => x"cb",
          5425 => x"d3",
          5426 => x"db",
          5427 => x"e3",
          5428 => x"eb",
          5429 => x"f3",
          5430 => x"fb",
          5431 => x"3b",
          5432 => x"3a",
          5433 => x"00",
          5434 => x"40",
          5435 => x"00",
          5436 => x"08",
          5437 => x"00",
          5438 => x"e2",
          5439 => x"e7",
          5440 => x"ef",
          5441 => x"c5",
          5442 => x"f4",
          5443 => x"f9",
          5444 => x"a2",
          5445 => x"92",
          5446 => x"fa",
          5447 => x"ba",
          5448 => x"bd",
          5449 => x"bb",
          5450 => x"02",
          5451 => x"56",
          5452 => x"57",
          5453 => x"10",
          5454 => x"1c",
          5455 => x"5f",
          5456 => x"66",
          5457 => x"67",
          5458 => x"59",
          5459 => x"6b",
          5460 => x"88",
          5461 => x"80",
          5462 => x"c0",
          5463 => x"c4",
          5464 => x"b4",
          5465 => x"29",
          5466 => x"64",
          5467 => x"48",
          5468 => x"1a",
          5469 => x"a0",
          5470 => x"17",
          5471 => x"01",
          5472 => x"32",
          5473 => x"4a",
          5474 => x"80",
          5475 => x"82",
          5476 => x"86",
          5477 => x"8a",
          5478 => x"8e",
          5479 => x"91",
          5480 => x"96",
          5481 => x"3d",
          5482 => x"20",
          5483 => x"a2",
          5484 => x"a6",
          5485 => x"aa",
          5486 => x"ae",
          5487 => x"b2",
          5488 => x"b5",
          5489 => x"ba",
          5490 => x"be",
          5491 => x"c2",
          5492 => x"c4",
          5493 => x"ca",
          5494 => x"10",
          5495 => x"de",
          5496 => x"f1",
          5497 => x"28",
          5498 => x"09",
          5499 => x"3d",
          5500 => x"41",
          5501 => x"53",
          5502 => x"55",
          5503 => x"8f",
          5504 => x"5d",
          5505 => x"61",
          5506 => x"65",
          5507 => x"96",
          5508 => x"6d",
          5509 => x"71",
          5510 => x"9f",
          5511 => x"79",
          5512 => x"64",
          5513 => x"81",
          5514 => x"85",
          5515 => x"44",
          5516 => x"8d",
          5517 => x"91",
          5518 => x"fd",
          5519 => x"04",
          5520 => x"8a",
          5521 => x"02",
          5522 => x"08",
          5523 => x"8e",
          5524 => x"f2",
          5525 => x"f4",
          5526 => x"f7",
          5527 => x"30",
          5528 => x"60",
          5529 => x"c1",
          5530 => x"c0",
          5531 => x"26",
          5532 => x"01",
          5533 => x"a0",
          5534 => x"10",
          5535 => x"30",
          5536 => x"51",
          5537 => x"5b",
          5538 => x"5f",
          5539 => x"0e",
          5540 => x"c9",
          5541 => x"db",
          5542 => x"eb",
          5543 => x"08",
          5544 => x"08",
          5545 => x"b9",
          5546 => x"01",
          5547 => x"e0",
          5548 => x"ec",
          5549 => x"4e",
          5550 => x"10",
          5551 => x"d0",
          5552 => x"60",
          5553 => x"75",
          5554 => x"00",
          5555 => x"00",
          5556 => x"40",
          5557 => x"00",
          5558 => x"48",
          5559 => x"00",
          5560 => x"50",
          5561 => x"00",
          5562 => x"58",
          5563 => x"00",
          5564 => x"60",
          5565 => x"00",
          5566 => x"68",
          5567 => x"00",
          5568 => x"70",
          5569 => x"00",
          5570 => x"78",
          5571 => x"00",
          5572 => x"80",
          5573 => x"00",
          5574 => x"88",
          5575 => x"00",
          5576 => x"8c",
          5577 => x"00",
          5578 => x"90",
          5579 => x"00",
          5580 => x"94",
          5581 => x"00",
          5582 => x"98",
          5583 => x"00",
          5584 => x"9c",
          5585 => x"00",
          5586 => x"a0",
          5587 => x"00",
          5588 => x"a4",
          5589 => x"00",
          5590 => x"ac",
          5591 => x"00",
          5592 => x"b0",
          5593 => x"00",
          5594 => x"b8",
          5595 => x"00",
          5596 => x"c0",
          5597 => x"00",
          5598 => x"c8",
          5599 => x"00",
          5600 => x"d0",
          5601 => x"00",
          5602 => x"d8",
          5603 => x"00",
          5604 => x"e0",
          5605 => x"00",
          5606 => x"00",
          5607 => x"ff",
          5608 => x"ff",
          5609 => x"ff",
          5610 => x"00",
          5611 => x"ff",
          5612 => x"00",
          5613 => x"00",
          5614 => x"00",
          5615 => x"00",
          5616 => x"01",
          5617 => x"00",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"00",
          5630 => x"00",
          5631 => x"00",
          5632 => x"00",
          5633 => x"00",
          5634 => x"04",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"87",
             1 => x"ed",
             2 => x"00",
             3 => x"00",
             4 => x"8c",
             5 => x"90",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"82",
            10 => x"06",
            11 => x"00",
            12 => x"06",
            13 => x"09",
            14 => x"09",
            15 => x"0b",
            16 => x"81",
            17 => x"09",
            18 => x"81",
            19 => x"00",
            20 => x"24",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"05",
            26 => x"0a",
            27 => x"53",
            28 => x"26",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"9f",
            45 => x"93",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"09",
            50 => x"53",
            51 => x"00",
            52 => x"53",
            53 => x"81",
            54 => x"07",
            55 => x"00",
            56 => x"81",
            57 => x"09",
            58 => x"00",
            59 => x"00",
            60 => x"81",
            61 => x"09",
            62 => x"04",
            63 => x"00",
            64 => x"81",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"09",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"51",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"83",
            78 => x"06",
            79 => x"00",
            80 => x"06",
            81 => x"83",
            82 => x"0b",
            83 => x"00",
            84 => x"8c",
            85 => x"80",
            86 => x"56",
            87 => x"04",
            88 => x"8c",
            89 => x"80",
            90 => x"56",
            91 => x"04",
            92 => x"70",
            93 => x"ff",
            94 => x"72",
            95 => x"51",
            96 => x"70",
            97 => x"06",
            98 => x"09",
            99 => x"51",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"05",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"04",
           126 => x"ff",
           127 => x"ff",
           128 => x"06",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"85",
           134 => x"0b",
           135 => x"0b",
           136 => x"c6",
           137 => x"0b",
           138 => x"0b",
           139 => x"88",
           140 => x"0b",
           141 => x"0b",
           142 => x"c9",
           143 => x"0b",
           144 => x"0b",
           145 => x"8d",
           146 => x"0b",
           147 => x"0b",
           148 => x"d1",
           149 => x"0b",
           150 => x"0b",
           151 => x"95",
           152 => x"0b",
           153 => x"0b",
           154 => x"d9",
           155 => x"0b",
           156 => x"0b",
           157 => x"9d",
           158 => x"0b",
           159 => x"0b",
           160 => x"e1",
           161 => x"0b",
           162 => x"0b",
           163 => x"a5",
           164 => x"0b",
           165 => x"0b",
           166 => x"e9",
           167 => x"0b",
           168 => x"0b",
           169 => x"ad",
           170 => x"0b",
           171 => x"0b",
           172 => x"f1",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"8c",
           193 => x"81",
           194 => x"c0",
           195 => x"b3",
           196 => x"c0",
           197 => x"b0",
           198 => x"c0",
           199 => x"af",
           200 => x"c0",
           201 => x"94",
           202 => x"c0",
           203 => x"b1",
           204 => x"c0",
           205 => x"80",
           206 => x"80",
           207 => x"0c",
           208 => x"08",
           209 => x"a4",
           210 => x"08",
           211 => x"a4",
           212 => x"08",
           213 => x"a4",
           214 => x"08",
           215 => x"a4",
           216 => x"a4",
           217 => x"e0",
           218 => x"e0",
           219 => x"82",
           220 => x"82",
           221 => x"04",
           222 => x"2d",
           223 => x"90",
           224 => x"e5",
           225 => x"80",
           226 => x"f6",
           227 => x"c0",
           228 => x"82",
           229 => x"80",
           230 => x"0c",
           231 => x"08",
           232 => x"a4",
           233 => x"a4",
           234 => x"e0",
           235 => x"e0",
           236 => x"82",
           237 => x"82",
           238 => x"04",
           239 => x"2d",
           240 => x"90",
           241 => x"88",
           242 => x"80",
           243 => x"8d",
           244 => x"c0",
           245 => x"82",
           246 => x"80",
           247 => x"0c",
           248 => x"08",
           249 => x"a4",
           250 => x"a4",
           251 => x"e0",
           252 => x"e0",
           253 => x"82",
           254 => x"82",
           255 => x"04",
           256 => x"2d",
           257 => x"90",
           258 => x"9d",
           259 => x"80",
           260 => x"84",
           261 => x"c0",
           262 => x"82",
           263 => x"80",
           264 => x"0c",
           265 => x"08",
           266 => x"a4",
           267 => x"a4",
           268 => x"e0",
           269 => x"e0",
           270 => x"82",
           271 => x"82",
           272 => x"04",
           273 => x"2d",
           274 => x"90",
           275 => x"c6",
           276 => x"80",
           277 => x"a5",
           278 => x"c0",
           279 => x"82",
           280 => x"80",
           281 => x"0c",
           282 => x"08",
           283 => x"a4",
           284 => x"a4",
           285 => x"e0",
           286 => x"e0",
           287 => x"82",
           288 => x"82",
           289 => x"04",
           290 => x"2d",
           291 => x"90",
           292 => x"88",
           293 => x"80",
           294 => x"82",
           295 => x"c0",
           296 => x"80",
           297 => x"80",
           298 => x"0c",
           299 => x"08",
           300 => x"a4",
           301 => x"a4",
           302 => x"e0",
           303 => x"e0",
           304 => x"82",
           305 => x"82",
           306 => x"04",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"10",
           311 => x"81",
           312 => x"05",
           313 => x"72",
           314 => x"72",
           315 => x"72",
           316 => x"10",
           317 => x"53",
           318 => x"fc",
           319 => x"84",
           320 => x"f0",
           321 => x"04",
           322 => x"e0",
           323 => x"a4",
           324 => x"08",
           325 => x"fc",
           326 => x"88",
           327 => x"52",
           328 => x"08",
           329 => x"0c",
           330 => x"70",
           331 => x"3d",
           332 => x"e0",
           333 => x"fb",
           334 => x"05",
           335 => x"70",
           336 => x"8f",
           337 => x"8c",
           338 => x"80",
           339 => x"0c",
           340 => x"8c",
           341 => x"08",
           342 => x"a4",
           343 => x"08",
           344 => x"fc",
           345 => x"05",
           346 => x"0b",
           347 => x"25",
           348 => x"90",
           349 => x"e0",
           350 => x"f8",
           351 => x"f8",
           352 => x"8d",
           353 => x"f4",
           354 => x"a4",
           355 => x"08",
           356 => x"34",
           357 => x"ff",
           358 => x"0c",
           359 => x"81",
           360 => x"0c",
           361 => x"fc",
           362 => x"e0",
           363 => x"e0",
           364 => x"e0",
           365 => x"98",
           366 => x"0c",
           367 => x"e0",
           368 => x"82",
           369 => x"e0",
           370 => x"a4",
           371 => x"82",
           372 => x"e0",
           373 => x"a4",
           374 => x"08",
           375 => x"08",
           376 => x"08",
           377 => x"8d",
           378 => x"e0",
           379 => x"a4",
           380 => x"08",
           381 => x"74",
           382 => x"08",
           383 => x"3d",
           384 => x"e0",
           385 => x"fb",
           386 => x"05",
           387 => x"0c",
           388 => x"54",
           389 => x"53",
           390 => x"52",
           391 => x"70",
           392 => x"82",
           393 => x"82",
           394 => x"0d",
           395 => x"a4",
           396 => x"3d",
           397 => x"e4",
           398 => x"05",
           399 => x"82",
           400 => x"11",
           401 => x"70",
           402 => x"72",
           403 => x"e0",
           404 => x"39",
           405 => x"53",
           406 => x"08",
           407 => x"53",
           408 => x"e0",
           409 => x"82",
           410 => x"e0",
           411 => x"06",
           412 => x"38",
           413 => x"53",
           414 => x"e0",
           415 => x"b9",
           416 => x"08",
           417 => x"09",
           418 => x"a4",
           419 => x"70",
           420 => x"38",
           421 => x"70",
           422 => x"06",
           423 => x"99",
           424 => x"22",
           425 => x"82",
           426 => x"d0",
           427 => x"33",
           428 => x"70",
           429 => x"51",
           430 => x"e0",
           431 => x"a4",
           432 => x"a4",
           433 => x"11",
           434 => x"08",
           435 => x"e8",
           436 => x"2c",
           437 => x"38",
           438 => x"e8",
           439 => x"05",
           440 => x"51",
           441 => x"e0",
           442 => x"2b",
           443 => x"88",
           444 => x"82",
           445 => x"b8",
           446 => x"22",
           447 => x"51",
           448 => x"e0",
           449 => x"2b",
           450 => x"8a",
           451 => x"e8",
           452 => x"05",
           453 => x"c4",
           454 => x"c4",
           455 => x"38",
           456 => x"70",
           457 => x"08",
           458 => x"e0",
           459 => x"07",
           460 => x"e4",
           461 => x"05",
           462 => x"82",
           463 => x"a8",
           464 => x"22",
           465 => x"82",
           466 => x"90",
           467 => x"22",
           468 => x"82",
           469 => x"f8",
           470 => x"22",
           471 => x"e0",
           472 => x"82",
           473 => x"d8",
           474 => x"22",
           475 => x"e0",
           476 => x"39",
           477 => x"05",
           478 => x"22",
           479 => x"a4",
           480 => x"82",
           481 => x"a8",
           482 => x"08",
           483 => x"84",
           484 => x"0c",
           485 => x"a4",
           486 => x"08",
           487 => x"72",
           488 => x"8c",
           489 => x"05",
           490 => x"08",
           491 => x"05",
           492 => x"fc",
           493 => x"05",
           494 => x"51",
           495 => x"38",
           496 => x"70",
           497 => x"82",
           498 => x"53",
           499 => x"53",
           500 => x"23",
           501 => x"05",
           502 => x"98",
           503 => x"f4",
           504 => x"05",
           505 => x"05",
           506 => x"82",
           507 => x"d8",
           508 => x"08",
           509 => x"84",
           510 => x"0c",
           511 => x"05",
           512 => x"22",
           513 => x"51",
           514 => x"82",
           515 => x"98",
           516 => x"e0",
           517 => x"a2",
           518 => x"72",
           519 => x"99",
           520 => x"08",
           521 => x"08",
           522 => x"05",
           523 => x"22",
           524 => x"22",
           525 => x"e0",
           526 => x"39",
           527 => x"70",
           528 => x"53",
           529 => x"a4",
           530 => x"08",
           531 => x"a4",
           532 => x"e0",
           533 => x"39",
           534 => x"82",
           535 => x"05",
           536 => x"70",
           537 => x"0c",
           538 => x"08",
           539 => x"82",
           540 => x"25",
           541 => x"05",
           542 => x"82",
           543 => x"e0",
           544 => x"e0",
           545 => x"a4",
           546 => x"06",
           547 => x"e4",
           548 => x"82",
           549 => x"39",
           550 => x"70",
           551 => x"e0",
           552 => x"0b",
           553 => x"90",
           554 => x"23",
           555 => x"70",
           556 => x"53",
           557 => x"a4",
           558 => x"08",
           559 => x"a4",
           560 => x"e0",
           561 => x"39",
           562 => x"82",
           563 => x"05",
           564 => x"70",
           565 => x"0c",
           566 => x"08",
           567 => x"82",
           568 => x"cf",
           569 => x"08",
           570 => x"82",
           571 => x"e0",
           572 => x"a4",
           573 => x"08",
           574 => x"56",
           575 => x"98",
           576 => x"a4",
           577 => x"08",
           578 => x"f0",
           579 => x"73",
           580 => x"f0",
           581 => x"e0",
           582 => x"df",
           583 => x"a4",
           584 => x"e0",
           585 => x"33",
           586 => x"a4",
           587 => x"08",
           588 => x"08",
           589 => x"a4",
           590 => x"e0",
           591 => x"a4",
           592 => x"e0",
           593 => x"a0",
           594 => x"82",
           595 => x"82",
           596 => x"2e",
           597 => x"a4",
           598 => x"54",
           599 => x"51",
           600 => x"05",
           601 => x"22",
           602 => x"2e",
           603 => x"05",
           604 => x"e0",
           605 => x"a4",
           606 => x"70",
           607 => x"2e",
           608 => x"ec",
           609 => x"a4",
           610 => x"08",
           611 => x"a4",
           612 => x"08",
           613 => x"2e",
           614 => x"a4",
           615 => x"72",
           616 => x"93",
           617 => x"08",
           618 => x"08",
           619 => x"c8",
           620 => x"05",
           621 => x"22",
           622 => x"51",
           623 => x"82",
           624 => x"98",
           625 => x"08",
           626 => x"72",
           627 => x"08",
           628 => x"53",
           629 => x"23",
           630 => x"05",
           631 => x"05",
           632 => x"82",
           633 => x"e0",
           634 => x"2a",
           635 => x"80",
           636 => x"e8",
           637 => x"2b",
           638 => x"51",
           639 => x"a4",
           640 => x"51",
           641 => x"05",
           642 => x"fc",
           643 => x"2b",
           644 => x"51",
           645 => x"a4",
           646 => x"51",
           647 => x"05",
           648 => x"22",
           649 => x"b0",
           650 => x"22",
           651 => x"a4",
           652 => x"70",
           653 => x"90",
           654 => x"08",
           655 => x"39",
           656 => x"70",
           657 => x"53",
           658 => x"a4",
           659 => x"8a",
           660 => x"a4",
           661 => x"70",
           662 => x"2e",
           663 => x"05",
           664 => x"a3",
           665 => x"22",
           666 => x"51",
           667 => x"e0",
           668 => x"51",
           669 => x"e4",
           670 => x"06",
           671 => x"38",
           672 => x"52",
           673 => x"a4",
           674 => x"2e",
           675 => x"a4",
           676 => x"a4",
           677 => x"3f",
           678 => x"70",
           679 => x"53",
           680 => x"a4",
           681 => x"54",
           682 => x"23",
           683 => x"53",
           684 => x"a4",
           685 => x"88",
           686 => x"08",
           687 => x"81",
           688 => x"b0",
           689 => x"33",
           690 => x"a4",
           691 => x"70",
           692 => x"90",
           693 => x"08",
           694 => x"39",
           695 => x"70",
           696 => x"53",
           697 => x"ec",
           698 => x"82",
           699 => x"90",
           700 => x"73",
           701 => x"88",
           702 => x"3f",
           703 => x"05",
           704 => x"81",
           705 => x"88",
           706 => x"fc",
           707 => x"ee",
           708 => x"33",
           709 => x"06",
           710 => x"f4",
           711 => x"82",
           712 => x"83",
           713 => x"ff",
           714 => x"08",
           715 => x"08",
           716 => x"e0",
           717 => x"82",
           718 => x"86",
           719 => x"a4",
           720 => x"d3",
           721 => x"82",
           722 => x"11",
           723 => x"f4",
           724 => x"53",
           725 => x"38",
           726 => x"52",
           727 => x"70",
           728 => x"e0",
           729 => x"82",
           730 => x"b7",
           731 => x"08",
           732 => x"e0",
           733 => x"e0",
           734 => x"82",
           735 => x"e0",
           736 => x"52",
           737 => x"e0",
           738 => x"2a",
           739 => x"80",
           740 => x"08",
           741 => x"72",
           742 => x"73",
           743 => x"80",
           744 => x"08",
           745 => x"9b",
           746 => x"88",
           747 => x"f8",
           748 => x"0b",
           749 => x"ea",
           750 => x"05",
           751 => x"06",
           752 => x"08",
           753 => x"a4",
           754 => x"e0",
           755 => x"82",
           756 => x"80",
           757 => x"08",
           758 => x"33",
           759 => x"82",
           760 => x"11",
           761 => x"05",
           762 => x"e0",
           763 => x"3d",
           764 => x"e0",
           765 => x"fd",
           766 => x"82",
           767 => x"82",
           768 => x"e4",
           769 => x"82",
           770 => x"82",
           771 => x"08",
           772 => x"0d",
           773 => x"05",
           774 => x"33",
           775 => x"81",
           776 => x"80",
           777 => x"a4",
           778 => x"82",
           779 => x"72",
           780 => x"08",
           781 => x"05",
           782 => x"fc",
           783 => x"72",
           784 => x"08",
           785 => x"a4",
           786 => x"08",
           787 => x"08",
           788 => x"ff",
           789 => x"0c",
           790 => x"82",
           791 => x"90",
           792 => x"98",
           793 => x"ff",
           794 => x"0c",
           795 => x"70",
           796 => x"53",
           797 => x"82",
           798 => x"e0",
           799 => x"02",
           800 => x"80",
           801 => x"0c",
           802 => x"85",
           803 => x"32",
           804 => x"53",
           805 => x"82",
           806 => x"f3",
           807 => x"08",
           808 => x"88",
           809 => x"08",
           810 => x"a4",
           811 => x"06",
           812 => x"e0",
           813 => x"a4",
           814 => x"a4",
           815 => x"08",
           816 => x"08",
           817 => x"ff",
           818 => x"0c",
           819 => x"f8",
           820 => x"f4",
           821 => x"f4",
           822 => x"3d",
           823 => x"e0",
           824 => x"fe",
           825 => x"82",
           826 => x"93",
           827 => x"e0",
           828 => x"e0",
           829 => x"02",
           830 => x"82",
           831 => x"11",
           832 => x"70",
           833 => x"72",
           834 => x"e0",
           835 => x"39",
           836 => x"85",
           837 => x"06",
           838 => x"80",
           839 => x"05",
           840 => x"08",
           841 => x"08",
           842 => x"8c",
           843 => x"a4",
           844 => x"54",
           845 => x"74",
           846 => x"08",
           847 => x"0c",
           848 => x"70",
           849 => x"51",
           850 => x"08",
           851 => x"8c",
           852 => x"88",
           853 => x"90",
           854 => x"82",
           855 => x"82",
           856 => x"11",
           857 => x"e0",
           858 => x"e0",
           859 => x"8a",
           860 => x"fc",
           861 => x"05",
           862 => x"0d",
           863 => x"a4",
           864 => x"3d",
           865 => x"08",
           866 => x"81",
           867 => x"2e",
           868 => x"08",
           869 => x"e0",
           870 => x"33",
           871 => x"51",
           872 => x"38",
           873 => x"82",
           874 => x"53",
           875 => x"51",
           876 => x"a4",
           877 => x"81",
           878 => x"08",
           879 => x"82",
           880 => x"51",
           881 => x"08",
           882 => x"82",
           883 => x"52",
           884 => x"e0",
           885 => x"70",
           886 => x"0c",
           887 => x"05",
           888 => x"88",
           889 => x"05",
           890 => x"a0",
           891 => x"ff",
           892 => x"0c",
           893 => x"88",
           894 => x"0c",
           895 => x"08",
           896 => x"88",
           897 => x"52",
           898 => x"82",
           899 => x"82",
           900 => x"25",
           901 => x"88",
           902 => x"05",
           903 => x"08",
           904 => x"f0",
           905 => x"fc",
           906 => x"95",
           907 => x"08",
           908 => x"08",
           909 => x"a4",
           910 => x"71",
           911 => x"82",
           912 => x"82",
           913 => x"13",
           914 => x"f8",
           915 => x"08",
           916 => x"05",
           917 => x"fc",
           918 => x"82",
           919 => x"51",
           920 => x"08",
           921 => x"82",
           922 => x"08",
           923 => x"0d",
           924 => x"82",
           925 => x"e0",
           926 => x"a4",
           927 => x"08",
           928 => x"38",
           929 => x"82",
           930 => x"81",
           931 => x"05",
           932 => x"08",
           933 => x"05",
           934 => x"e0",
           935 => x"a4",
           936 => x"a4",
           937 => x"08",
           938 => x"90",
           939 => x"f8",
           940 => x"05",
           941 => x"90",
           942 => x"05",
           943 => x"90",
           944 => x"05",
           945 => x"e0",
           946 => x"82",
           947 => x"e0",
           948 => x"82",
           949 => x"e0",
           950 => x"a4",
           951 => x"33",
           952 => x"a4",
           953 => x"e0",
           954 => x"a4",
           955 => x"e0",
           956 => x"a4",
           957 => x"38",
           958 => x"51",
           959 => x"05",
           960 => x"f8",
           961 => x"05",
           962 => x"e0",
           963 => x"82",
           964 => x"ad",
           965 => x"08",
           966 => x"3d",
           967 => x"e0",
           968 => x"fe",
           969 => x"05",
           970 => x"0c",
           971 => x"52",
           972 => x"05",
           973 => x"fc",
           974 => x"51",
           975 => x"82",
           976 => x"05",
           977 => x"82",
           978 => x"e0",
           979 => x"82",
           980 => x"82",
           981 => x"08",
           982 => x"0d",
           983 => x"82",
           984 => x"e0",
           985 => x"33",
           986 => x"81",
           987 => x"0c",
           988 => x"53",
           989 => x"08",
           990 => x"a4",
           991 => x"06",
           992 => x"be",
           993 => x"08",
           994 => x"3d",
           995 => x"e0",
           996 => x"fd",
           997 => x"05",
           998 => x"0c",
           999 => x"82",
          1000 => x"e0",
          1001 => x"80",
          1002 => x"05",
          1003 => x"90",
          1004 => x"05",
          1005 => x"90",
          1006 => x"05",
          1007 => x"a4",
          1008 => x"82",
          1009 => x"05",
          1010 => x"82",
          1011 => x"52",
          1012 => x"fc",
          1013 => x"08",
          1014 => x"e0",
          1015 => x"e0",
          1016 => x"e0",
          1017 => x"02",
          1018 => x"82",
          1019 => x"2e",
          1020 => x"8c",
          1021 => x"a4",
          1022 => x"e0",
          1023 => x"a4",
          1024 => x"81",
          1025 => x"71",
          1026 => x"e0",
          1027 => x"33",
          1028 => x"81",
          1029 => x"0c",
          1030 => x"8d",
          1031 => x"fc",
          1032 => x"a4",
          1033 => x"e0",
          1034 => x"a4",
          1035 => x"38",
          1036 => x"90",
          1037 => x"82",
          1038 => x"33",
          1039 => x"82",
          1040 => x"d7",
          1041 => x"08",
          1042 => x"05",
          1043 => x"08",
          1044 => x"81",
          1045 => x"0c",
          1046 => x"05",
          1047 => x"8c",
          1048 => x"70",
          1049 => x"53",
          1050 => x"0b",
          1051 => x"82",
          1052 => x"e0",
          1053 => x"a4",
          1054 => x"82",
          1055 => x"e0",
          1056 => x"e0",
          1057 => x"8d",
          1058 => x"e0",
          1059 => x"a4",
          1060 => x"53",
          1061 => x"e0",
          1062 => x"fc",
          1063 => x"fc",
          1064 => x"e0",
          1065 => x"82",
          1066 => x"e0",
          1067 => x"80",
          1068 => x"05",
          1069 => x"05",
          1070 => x"05",
          1071 => x"98",
          1072 => x"05",
          1073 => x"05",
          1074 => x"0d",
          1075 => x"a4",
          1076 => x"3d",
          1077 => x"08",
          1078 => x"82",
          1079 => x"38",
          1080 => x"05",
          1081 => x"08",
          1082 => x"e0",
          1083 => x"82",
          1084 => x"81",
          1085 => x"9f",
          1086 => x"08",
          1087 => x"05",
          1088 => x"08",
          1089 => x"82",
          1090 => x"05",
          1091 => x"82",
          1092 => x"e0",
          1093 => x"82",
          1094 => x"82",
          1095 => x"e0",
          1096 => x"a4",
          1097 => x"82",
          1098 => x"e0",
          1099 => x"a4",
          1100 => x"08",
          1101 => x"38",
          1102 => x"81",
          1103 => x"0c",
          1104 => x"ff",
          1105 => x"0c",
          1106 => x"80",
          1107 => x"8c",
          1108 => x"08",
          1109 => x"34",
          1110 => x"81",
          1111 => x"0c",
          1112 => x"88",
          1113 => x"51",
          1114 => x"04",
          1115 => x"a4",
          1116 => x"08",
          1117 => x"08",
          1118 => x"e0",
          1119 => x"53",
          1120 => x"04",
          1121 => x"a4",
          1122 => x"e0",
          1123 => x"a4",
          1124 => x"38",
          1125 => x"51",
          1126 => x"70",
          1127 => x"52",
          1128 => x"05",
          1129 => x"0c",
          1130 => x"80",
          1131 => x"88",
          1132 => x"e0",
          1133 => x"05",
          1134 => x"e0",
          1135 => x"a4",
          1136 => x"08",
          1137 => x"08",
          1138 => x"e0",
          1139 => x"05",
          1140 => x"08",
          1141 => x"08",
          1142 => x"0b",
          1143 => x"82",
          1144 => x"05",
          1145 => x"a4",
          1146 => x"06",
          1147 => x"05",
          1148 => x"05",
          1149 => x"a4",
          1150 => x"e0",
          1151 => x"a4",
          1152 => x"08",
          1153 => x"08",
          1154 => x"fc",
          1155 => x"05",
          1156 => x"05",
          1157 => x"88",
          1158 => x"a4",
          1159 => x"08",
          1160 => x"38",
          1161 => x"10",
          1162 => x"ff",
          1163 => x"08",
          1164 => x"a4",
          1165 => x"08",
          1166 => x"a4",
          1167 => x"a4",
          1168 => x"08",
          1169 => x"f4",
          1170 => x"a4",
          1171 => x"71",
          1172 => x"0c",
          1173 => x"81",
          1174 => x"0c",
          1175 => x"82",
          1176 => x"82",
          1177 => x"31",
          1178 => x"82",
          1179 => x"05",
          1180 => x"51",
          1181 => x"fe",
          1182 => x"05",
          1183 => x"f0",
          1184 => x"88",
          1185 => x"05",
          1186 => x"05",
          1187 => x"e8",
          1188 => x"3d",
          1189 => x"e0",
          1190 => x"f8",
          1191 => x"05",
          1192 => x"0c",
          1193 => x"fc",
          1194 => x"90",
          1195 => x"0c",
          1196 => x"08",
          1197 => x"f0",
          1198 => x"05",
          1199 => x"f8",
          1200 => x"fc",
          1201 => x"08",
          1202 => x"f8",
          1203 => x"05",
          1204 => x"08",
          1205 => x"8c",
          1206 => x"ec",
          1207 => x"e0",
          1208 => x"a4",
          1209 => x"08",
          1210 => x"a4",
          1211 => x"a4",
          1212 => x"e0",
          1213 => x"a4",
          1214 => x"08",
          1215 => x"08",
          1216 => x"fc",
          1217 => x"70",
          1218 => x"08",
          1219 => x"82",
          1220 => x"e0",
          1221 => x"a4",
          1222 => x"e0",
          1223 => x"e0",
          1224 => x"82",
          1225 => x"e0",
          1226 => x"a4",
          1227 => x"a4",
          1228 => x"08",
          1229 => x"70",
          1230 => x"08",
          1231 => x"82",
          1232 => x"e0",
          1233 => x"a4",
          1234 => x"e0",
          1235 => x"e0",
          1236 => x"82",
          1237 => x"e0",
          1238 => x"a4",
          1239 => x"a4",
          1240 => x"e0",
          1241 => x"e0",
          1242 => x"70",
          1243 => x"70",
          1244 => x"05",
          1245 => x"0c",
          1246 => x"53",
          1247 => x"0c",
          1248 => x"e0",
          1249 => x"a4",
          1250 => x"a4",
          1251 => x"3f",
          1252 => x"a4",
          1253 => x"a4",
          1254 => x"82",
          1255 => x"3d",
          1256 => x"e0",
          1257 => x"fe",
          1258 => x"05",
          1259 => x"05",
          1260 => x"08",
          1261 => x"3d",
          1262 => x"e0",
          1263 => x"f6",
          1264 => x"08",
          1265 => x"8c",
          1266 => x"e0",
          1267 => x"8e",
          1268 => x"e0",
          1269 => x"39",
          1270 => x"82",
          1271 => x"e0",
          1272 => x"a3",
          1273 => x"08",
          1274 => x"08",
          1275 => x"71",
          1276 => x"0c",
          1277 => x"e4",
          1278 => x"05",
          1279 => x"05",
          1280 => x"08",
          1281 => x"82",
          1282 => x"05",
          1283 => x"05",
          1284 => x"08",
          1285 => x"08",
          1286 => x"82",
          1287 => x"05",
          1288 => x"05",
          1289 => x"80",
          1290 => x"0c",
          1291 => x"f8",
          1292 => x"08",
          1293 => x"88",
          1294 => x"05",
          1295 => x"05",
          1296 => x"08",
          1297 => x"31",
          1298 => x"71",
          1299 => x"0c",
          1300 => x"f0",
          1301 => x"05",
          1302 => x"e0",
          1303 => x"e0",
          1304 => x"82",
          1305 => x"2a",
          1306 => x"f4",
          1307 => x"05",
          1308 => x"f0",
          1309 => x"88",
          1310 => x"05",
          1311 => x"08",
          1312 => x"fc",
          1313 => x"82",
          1314 => x"e0",
          1315 => x"82",
          1316 => x"e0",
          1317 => x"a4",
          1318 => x"a4",
          1319 => x"e0",
          1320 => x"a4",
          1321 => x"e0",
          1322 => x"55",
          1323 => x"39",
          1324 => x"70",
          1325 => x"52",
          1326 => x"82",
          1327 => x"e0",
          1328 => x"02",
          1329 => x"9f",
          1330 => x"0c",
          1331 => x"82",
          1332 => x"82",
          1333 => x"e0",
          1334 => x"a4",
          1335 => x"a4",
          1336 => x"08",
          1337 => x"f8",
          1338 => x"08",
          1339 => x"08",
          1340 => x"8c",
          1341 => x"05",
          1342 => x"f4",
          1343 => x"8c",
          1344 => x"05",
          1345 => x"08",
          1346 => x"0c",
          1347 => x"54",
          1348 => x"53",
          1349 => x"98",
          1350 => x"05",
          1351 => x"f8",
          1352 => x"0c",
          1353 => x"e0",
          1354 => x"02",
          1355 => x"80",
          1356 => x"34",
          1357 => x"53",
          1358 => x"88",
          1359 => x"33",
          1360 => x"05",
          1361 => x"a0",
          1362 => x"e0",
          1363 => x"81",
          1364 => x"e0",
          1365 => x"ad",
          1366 => x"0b",
          1367 => x"82",
          1368 => x"08",
          1369 => x"53",
          1370 => x"05",
          1371 => x"33",
          1372 => x"81",
          1373 => x"05",
          1374 => x"70",
          1375 => x"a4",
          1376 => x"08",
          1377 => x"e8",
          1378 => x"05",
          1379 => x"e0",
          1380 => x"2e",
          1381 => x"82",
          1382 => x"e0",
          1383 => x"81",
          1384 => x"72",
          1385 => x"34",
          1386 => x"a4",
          1387 => x"08",
          1388 => x"71",
          1389 => x"82",
          1390 => x"fe",
          1391 => x"33",
          1392 => x"0b",
          1393 => x"83",
          1394 => x"05",
          1395 => x"82",
          1396 => x"72",
          1397 => x"0b",
          1398 => x"82",
          1399 => x"08",
          1400 => x"a4",
          1401 => x"27",
          1402 => x"05",
          1403 => x"8d",
          1404 => x"ec",
          1405 => x"82",
          1406 => x"0b",
          1407 => x"82",
          1408 => x"a0",
          1409 => x"a4",
          1410 => x"73",
          1411 => x"f8",
          1412 => x"82",
          1413 => x"e0",
          1414 => x"51",
          1415 => x"05",
          1416 => x"33",
          1417 => x"e0",
          1418 => x"51",
          1419 => x"05",
          1420 => x"33",
          1421 => x"0b",
          1422 => x"81",
          1423 => x"05",
          1424 => x"33",
          1425 => x"80",
          1426 => x"0c",
          1427 => x"f4",
          1428 => x"fc",
          1429 => x"f8",
          1430 => x"08",
          1431 => x"88",
          1432 => x"0c",
          1433 => x"72",
          1434 => x"34",
          1435 => x"f0",
          1436 => x"38",
          1437 => x"30",
          1438 => x"82",
          1439 => x"e0",
          1440 => x"53",
          1441 => x"05",
          1442 => x"08",
          1443 => x"82",
          1444 => x"08",
          1445 => x"0d",
          1446 => x"05",
          1447 => x"08",
          1448 => x"08",
          1449 => x"72",
          1450 => x"f8",
          1451 => x"72",
          1452 => x"82",
          1453 => x"08",
          1454 => x"82",
          1455 => x"72",
          1456 => x"81",
          1457 => x"34",
          1458 => x"70",
          1459 => x"51",
          1460 => x"f8",
          1461 => x"05",
          1462 => x"06",
          1463 => x"88",
          1464 => x"0c",
          1465 => x"e0",
          1466 => x"a4",
          1467 => x"08",
          1468 => x"e8",
          1469 => x"82",
          1470 => x"f8",
          1471 => x"0b",
          1472 => x"82",
          1473 => x"08",
          1474 => x"53",
          1475 => x"05",
          1476 => x"e0",
          1477 => x"a4",
          1478 => x"05",
          1479 => x"33",
          1480 => x"80",
          1481 => x"05",
          1482 => x"81",
          1483 => x"0c",
          1484 => x"f8",
          1485 => x"38",
          1486 => x"53",
          1487 => x"80",
          1488 => x"0c",
          1489 => x"a4",
          1490 => x"e0",
          1491 => x"73",
          1492 => x"f8",
          1493 => x"38",
          1494 => x"08",
          1495 => x"0b",
          1496 => x"80",
          1497 => x"0c",
          1498 => x"53",
          1499 => x"e0",
          1500 => x"e0",
          1501 => x"08",
          1502 => x"72",
          1503 => x"82",
          1504 => x"11",
          1505 => x"f8",
          1506 => x"05",
          1507 => x"82",
          1508 => x"11",
          1509 => x"f8",
          1510 => x"05",
          1511 => x"80",
          1512 => x"0c",
          1513 => x"f8",
          1514 => x"05",
          1515 => x"38",
          1516 => x"05",
          1517 => x"08",
          1518 => x"08",
          1519 => x"08",
          1520 => x"a4",
          1521 => x"08",
          1522 => x"71",
          1523 => x"53",
          1524 => x"05",
          1525 => x"08",
          1526 => x"90",
          1527 => x"08",
          1528 => x"0c",
          1529 => x"82",
          1530 => x"0c",
          1531 => x"ec",
          1532 => x"05",
          1533 => x"0d",
          1534 => x"0d",
          1535 => x"74",
          1536 => x"77",
          1537 => x"80",
          1538 => x"2e",
          1539 => x"55",
          1540 => x"82",
          1541 => x"dc",
          1542 => x"e0",
          1543 => x"52",
          1544 => x"08",
          1545 => x"81",
          1546 => x"81",
          1547 => x"c4",
          1548 => x"0c",
          1549 => x"82",
          1550 => x"73",
          1551 => x"71",
          1552 => x"71",
          1553 => x"80",
          1554 => x"39",
          1555 => x"82",
          1556 => x"be",
          1557 => x"b0",
          1558 => x"51",
          1559 => x"80",
          1560 => x"c8",
          1561 => x"39",
          1562 => x"bf",
          1563 => x"51",
          1564 => x"39",
          1565 => x"c0",
          1566 => x"51",
          1567 => x"39",
          1568 => x"c0",
          1569 => x"51",
          1570 => x"fb",
          1571 => x"87",
          1572 => x"87",
          1573 => x"52",
          1574 => x"98",
          1575 => x"82",
          1576 => x"52",
          1577 => x"3f",
          1578 => x"66",
          1579 => x"5b",
          1580 => x"07",
          1581 => x"56",
          1582 => x"56",
          1583 => x"51",
          1584 => x"81",
          1585 => x"56",
          1586 => x"08",
          1587 => x"82",
          1588 => x"0c",
          1589 => x"d4",
          1590 => x"75",
          1591 => x"98",
          1592 => x"38",
          1593 => x"74",
          1594 => x"96",
          1595 => x"3f",
          1596 => x"7b",
          1597 => x"57",
          1598 => x"82",
          1599 => x"08",
          1600 => x"56",
          1601 => x"0d",
          1602 => x"05",
          1603 => x"80",
          1604 => x"3f",
          1605 => x"80",
          1606 => x"38",
          1607 => x"55",
          1608 => x"52",
          1609 => x"08",
          1610 => x"e0",
          1611 => x"3d",
          1612 => x"80",
          1613 => x"41",
          1614 => x"a4",
          1615 => x"08",
          1616 => x"a8",
          1617 => x"d0",
          1618 => x"82",
          1619 => x"c1",
          1620 => x"c1",
          1621 => x"55",
          1622 => x"90",
          1623 => x"38",
          1624 => x"7a",
          1625 => x"c1",
          1626 => x"39",
          1627 => x"3f",
          1628 => x"19",
          1629 => x"08",
          1630 => x"99",
          1631 => x"ff",
          1632 => x"39",
          1633 => x"38",
          1634 => x"ff",
          1635 => x"ec",
          1636 => x"55",
          1637 => x"cd",
          1638 => x"f0",
          1639 => x"74",
          1640 => x"70",
          1641 => x"27",
          1642 => x"74",
          1643 => x"06",
          1644 => x"80",
          1645 => x"8a",
          1646 => x"51",
          1647 => x"a0",
          1648 => x"ff",
          1649 => x"8c",
          1650 => x"80",
          1651 => x"08",
          1652 => x"76",
          1653 => x"80",
          1654 => x"08",
          1655 => x"32",
          1656 => x"70",
          1657 => x"58",
          1658 => x"24",
          1659 => x"38",
          1660 => x"b4",
          1661 => x"0c",
          1662 => x"02",
          1663 => x"be",
          1664 => x"fc",
          1665 => x"e8",
          1666 => x"84",
          1667 => x"e9",
          1668 => x"ab",
          1669 => x"a2",
          1670 => x"3d",
          1671 => x"a6",
          1672 => x"82",
          1673 => x"51",
          1674 => x"81",
          1675 => x"38",
          1676 => x"cc",
          1677 => x"95",
          1678 => x"51",
          1679 => x"51",
          1680 => x"9a",
          1681 => x"72",
          1682 => x"71",
          1683 => x"e5",
          1684 => x"3f",
          1685 => x"2a",
          1686 => x"2e",
          1687 => x"82",
          1688 => x"51",
          1689 => x"81",
          1690 => x"38",
          1691 => x"94",
          1692 => x"9d",
          1693 => x"51",
          1694 => x"51",
          1695 => x"99",
          1696 => x"72",
          1697 => x"71",
          1698 => x"ed",
          1699 => x"3f",
          1700 => x"2a",
          1701 => x"2e",
          1702 => x"82",
          1703 => x"51",
          1704 => x"3d",
          1705 => x"84",
          1706 => x"56",
          1707 => x"0b",
          1708 => x"a9",
          1709 => x"82",
          1710 => x"82",
          1711 => x"98",
          1712 => x"51",
          1713 => x"9c",
          1714 => x"54",
          1715 => x"38",
          1716 => x"51",
          1717 => x"08",
          1718 => x"08",
          1719 => x"f7",
          1720 => x"0b",
          1721 => x"0b",
          1722 => x"2e",
          1723 => x"9c",
          1724 => x"3f",
          1725 => x"3d",
          1726 => x"41",
          1727 => x"5f",
          1728 => x"3f",
          1729 => x"59",
          1730 => x"38",
          1731 => x"a8",
          1732 => x"53",
          1733 => x"89",
          1734 => x"2e",
          1735 => x"e5",
          1736 => x"e4",
          1737 => x"70",
          1738 => x"fd",
          1739 => x"51",
          1740 => x"90",
          1741 => x"80",
          1742 => x"c2",
          1743 => x"d2",
          1744 => x"80",
          1745 => x"80",
          1746 => x"c0",
          1747 => x"24",
          1748 => x"8c",
          1749 => x"2e",
          1750 => x"92",
          1751 => x"38",
          1752 => x"8a",
          1753 => x"8d",
          1754 => x"78",
          1755 => x"90",
          1756 => x"38",
          1757 => x"11",
          1758 => x"3f",
          1759 => x"c5",
          1760 => x"ff",
          1761 => x"e0",
          1762 => x"b5",
          1763 => x"05",
          1764 => x"08",
          1765 => x"82",
          1766 => x"64",
          1767 => x"ec",
          1768 => x"05",
          1769 => x"81",
          1770 => x"53",
          1771 => x"82",
          1772 => x"38",
          1773 => x"84",
          1774 => x"98",
          1775 => x"3d",
          1776 => x"51",
          1777 => x"80",
          1778 => x"51",
          1779 => x"64",
          1780 => x"70",
          1781 => x"81",
          1782 => x"80",
          1783 => x"e4",
          1784 => x"fc",
          1785 => x"53",
          1786 => x"82",
          1787 => x"38",
          1788 => x"84",
          1789 => x"98",
          1790 => x"c5",
          1791 => x"5a",
          1792 => x"33",
          1793 => x"2e",
          1794 => x"33",
          1795 => x"ff",
          1796 => x"05",
          1797 => x"8e",
          1798 => x"80",
          1799 => x"e4",
          1800 => x"38",
          1801 => x"2e",
          1802 => x"80",
          1803 => x"78",
          1804 => x"08",
          1805 => x"59",
          1806 => x"c4",
          1807 => x"33",
          1808 => x"de",
          1809 => x"fa",
          1810 => x"82",
          1811 => x"de",
          1812 => x"3d",
          1813 => x"51",
          1814 => x"80",
          1815 => x"78",
          1816 => x"08",
          1817 => x"33",
          1818 => x"de",
          1819 => x"fe",
          1820 => x"82",
          1821 => x"de",
          1822 => x"38",
          1823 => x"82",
          1824 => x"88",
          1825 => x"39",
          1826 => x"b5",
          1827 => x"05",
          1828 => x"08",
          1829 => x"5c",
          1830 => x"7a",
          1831 => x"9f",
          1832 => x"5a",
          1833 => x"2e",
          1834 => x"51",
          1835 => x"54",
          1836 => x"f6",
          1837 => x"39",
          1838 => x"84",
          1839 => x"98",
          1840 => x"3d",
          1841 => x"51",
          1842 => x"80",
          1843 => x"cf",
          1844 => x"45",
          1845 => x"84",
          1846 => x"98",
          1847 => x"70",
          1848 => x"ff",
          1849 => x"53",
          1850 => x"8e",
          1851 => x"ae",
          1852 => x"9f",
          1853 => x"ff",
          1854 => x"e0",
          1855 => x"59",
          1856 => x"64",
          1857 => x"c5",
          1858 => x"a6",
          1859 => x"ff",
          1860 => x"e0",
          1861 => x"b5",
          1862 => x"05",
          1863 => x"08",
          1864 => x"80",
          1865 => x"5b",
          1866 => x"11",
          1867 => x"3f",
          1868 => x"dd",
          1869 => x"c5",
          1870 => x"fb",
          1871 => x"51",
          1872 => x"33",
          1873 => x"78",
          1874 => x"42",
          1875 => x"53",
          1876 => x"82",
          1877 => x"61",
          1878 => x"70",
          1879 => x"a9",
          1880 => x"d4",
          1881 => x"f4",
          1882 => x"fb",
          1883 => x"f6",
          1884 => x"53",
          1885 => x"82",
          1886 => x"61",
          1887 => x"42",
          1888 => x"84",
          1889 => x"98",
          1890 => x"70",
          1891 => x"ff",
          1892 => x"53",
          1893 => x"b6",
          1894 => x"ae",
          1895 => x"9b",
          1896 => x"ff",
          1897 => x"e0",
          1898 => x"61",
          1899 => x"ff",
          1900 => x"b9",
          1901 => x"ff",
          1902 => x"e3",
          1903 => x"2e",
          1904 => x"f4",
          1905 => x"78",
          1906 => x"ff",
          1907 => x"e0",
          1908 => x"64",
          1909 => x"e1",
          1910 => x"98",
          1911 => x"e0",
          1912 => x"ff",
          1913 => x"c6",
          1914 => x"9c",
          1915 => x"e4",
          1916 => x"ff",
          1917 => x"39",
          1918 => x"f4",
          1919 => x"c9",
          1920 => x"82",
          1921 => x"38",
          1922 => x"ff",
          1923 => x"e0",
          1924 => x"78",
          1925 => x"98",
          1926 => x"98",
          1927 => x"5b",
          1928 => x"24",
          1929 => x"80",
          1930 => x"80",
          1931 => x"55",
          1932 => x"c7",
          1933 => x"51",
          1934 => x"52",
          1935 => x"ac",
          1936 => x"fc",
          1937 => x"b5",
          1938 => x"e1",
          1939 => x"82",
          1940 => x"05",
          1941 => x"b4",
          1942 => x"65",
          1943 => x"90",
          1944 => x"05",
          1945 => x"08",
          1946 => x"70",
          1947 => x"5f",
          1948 => x"81",
          1949 => x"2e",
          1950 => x"06",
          1951 => x"81",
          1952 => x"89",
          1953 => x"89",
          1954 => x"84",
          1955 => x"a5",
          1956 => x"f4",
          1957 => x"80",
          1958 => x"94",
          1959 => x"80",
          1960 => x"e0",
          1961 => x"53",
          1962 => x"80",
          1963 => x"75",
          1964 => x"54",
          1965 => x"ca",
          1966 => x"2b",
          1967 => x"52",
          1968 => x"e0",
          1969 => x"83",
          1970 => x"80",
          1971 => x"81",
          1972 => x"83",
          1973 => x"5c",
          1974 => x"88",
          1975 => x"fc",
          1976 => x"3f",
          1977 => x"3f",
          1978 => x"3f",
          1979 => x"81",
          1980 => x"80",
          1981 => x"54",
          1982 => x"2e",
          1983 => x"a0",
          1984 => x"13",
          1985 => x"a2",
          1986 => x"13",
          1987 => x"2e",
          1988 => x"81",
          1989 => x"70",
          1990 => x"80",
          1991 => x"39",
          1992 => x"54",
          1993 => x"70",
          1994 => x"80",
          1995 => x"09",
          1996 => x"a2",
          1997 => x"07",
          1998 => x"38",
          1999 => x"71",
          2000 => x"98",
          2001 => x"0d",
          2002 => x"38",
          2003 => x"d7",
          2004 => x"38",
          2005 => x"82",
          2006 => x"fc",
          2007 => x"05",
          2008 => x"81",
          2009 => x"51",
          2010 => x"38",
          2011 => x"97",
          2012 => x"51",
          2013 => x"38",
          2014 => x"bb",
          2015 => x"55",
          2016 => x"d9",
          2017 => x"73",
          2018 => x"0b",
          2019 => x"87",
          2020 => x"87",
          2021 => x"87",
          2022 => x"87",
          2023 => x"87",
          2024 => x"87",
          2025 => x"98",
          2026 => x"0c",
          2027 => x"80",
          2028 => x"3d",
          2029 => x"87",
          2030 => x"87",
          2031 => x"23",
          2032 => x"82",
          2033 => x"5a",
          2034 => x"b0",
          2035 => x"c0",
          2036 => x"34",
          2037 => x"86",
          2038 => x"5c",
          2039 => x"a0",
          2040 => x"7d",
          2041 => x"7b",
          2042 => x"33",
          2043 => x"33",
          2044 => x"33",
          2045 => x"82",
          2046 => x"8f",
          2047 => x"97",
          2048 => x"2e",
          2049 => x"72",
          2050 => x"74",
          2051 => x"86",
          2052 => x"f0",
          2053 => x"70",
          2054 => x"09",
          2055 => x"81",
          2056 => x"54",
          2057 => x"25",
          2058 => x"ab",
          2059 => x"3d",
          2060 => x"83",
          2061 => x"ff",
          2062 => x"2b",
          2063 => x"56",
          2064 => x"72",
          2065 => x"04",
          2066 => x"82",
          2067 => x"58",
          2068 => x"75",
          2069 => x"94",
          2070 => x"81",
          2071 => x"8c",
          2072 => x"51",
          2073 => x"70",
          2074 => x"8d",
          2075 => x"51",
          2076 => x"ff",
          2077 => x"70",
          2078 => x"90",
          2079 => x"98",
          2080 => x"0d",
          2081 => x"9f",
          2082 => x"b0",
          2083 => x"0d",
          2084 => x"2e",
          2085 => x"8d",
          2086 => x"70",
          2087 => x"94",
          2088 => x"87",
          2089 => x"96",
          2090 => x"72",
          2091 => x"70",
          2092 => x"74",
          2093 => x"72",
          2094 => x"70",
          2095 => x"38",
          2096 => x"94",
          2097 => x"87",
          2098 => x"80",
          2099 => x"0d",
          2100 => x"74",
          2101 => x"57",
          2102 => x"81",
          2103 => x"33",
          2104 => x"58",
          2105 => x"2e",
          2106 => x"70",
          2107 => x"53",
          2108 => x"71",
          2109 => x"70",
          2110 => x"06",
          2111 => x"71",
          2112 => x"70",
          2113 => x"51",
          2114 => x"2e",
          2115 => x"77",
          2116 => x"81",
          2117 => x"86",
          2118 => x"3d",
          2119 => x"b0",
          2120 => x"87",
          2121 => x"86",
          2122 => x"08",
          2123 => x"51",
          2124 => x"81",
          2125 => x"52",
          2126 => x"94",
          2127 => x"06",
          2128 => x"0d",
          2129 => x"08",
          2130 => x"04",
          2131 => x"70",
          2132 => x"94",
          2133 => x"87",
          2134 => x"82",
          2135 => x"ff",
          2136 => x"81",
          2137 => x"52",
          2138 => x"94",
          2139 => x"70",
          2140 => x"e0",
          2141 => x"3d",
          2142 => x"9c",
          2143 => x"2e",
          2144 => x"08",
          2145 => x"a8",
          2146 => x"9e",
          2147 => x"c0",
          2148 => x"87",
          2149 => x"0c",
          2150 => x"c8",
          2151 => x"de",
          2152 => x"82",
          2153 => x"08",
          2154 => x"b8",
          2155 => x"9e",
          2156 => x"c0",
          2157 => x"87",
          2158 => x"0c",
          2159 => x"82",
          2160 => x"08",
          2161 => x"88",
          2162 => x"9e",
          2163 => x"0b",
          2164 => x"c0",
          2165 => x"06",
          2166 => x"38",
          2167 => x"80",
          2168 => x"88",
          2169 => x"80",
          2170 => x"de",
          2171 => x"90",
          2172 => x"52",
          2173 => x"52",
          2174 => x"87",
          2175 => x"80",
          2176 => x"83",
          2177 => x"34",
          2178 => x"70",
          2179 => x"70",
          2180 => x"82",
          2181 => x"9e",
          2182 => x"51",
          2183 => x"81",
          2184 => x"0b",
          2185 => x"80",
          2186 => x"2e",
          2187 => x"ff",
          2188 => x"08",
          2189 => x"52",
          2190 => x"71",
          2191 => x"c0",
          2192 => x"06",
          2193 => x"38",
          2194 => x"80",
          2195 => x"80",
          2196 => x"80",
          2197 => x"df",
          2198 => x"90",
          2199 => x"52",
          2200 => x"71",
          2201 => x"90",
          2202 => x"2a",
          2203 => x"34",
          2204 => x"70",
          2205 => x"80",
          2206 => x"df",
          2207 => x"70",
          2208 => x"51",
          2209 => x"0b",
          2210 => x"06",
          2211 => x"38",
          2212 => x"87",
          2213 => x"51",
          2214 => x"3d",
          2215 => x"9c",
          2216 => x"f8",
          2217 => x"82",
          2218 => x"82",
          2219 => x"82",
          2220 => x"94",
          2221 => x"d8",
          2222 => x"51",
          2223 => x"33",
          2224 => x"de",
          2225 => x"54",
          2226 => x"f9",
          2227 => x"80",
          2228 => x"82",
          2229 => x"c9",
          2230 => x"de",
          2231 => x"38",
          2232 => x"08",
          2233 => x"ff",
          2234 => x"54",
          2235 => x"c4",
          2236 => x"52",
          2237 => x"3f",
          2238 => x"2e",
          2239 => x"82",
          2240 => x"82",
          2241 => x"8e",
          2242 => x"ca",
          2243 => x"df",
          2244 => x"38",
          2245 => x"a8",
          2246 => x"f9",
          2247 => x"82",
          2248 => x"82",
          2249 => x"89",
          2250 => x"c4",
          2251 => x"80",
          2252 => x"ff",
          2253 => x"54",
          2254 => x"f4",
          2255 => x"82",
          2256 => x"82",
          2257 => x"82",
          2258 => x"82",
          2259 => x"51",
          2260 => x"08",
          2261 => x"e1",
          2262 => x"cb",
          2263 => x"cc",
          2264 => x"de",
          2265 => x"ff",
          2266 => x"56",
          2267 => x"b7",
          2268 => x"84",
          2269 => x"82",
          2270 => x"51",
          2271 => x"33",
          2272 => x"de",
          2273 => x"75",
          2274 => x"98",
          2275 => x"31",
          2276 => x"82",
          2277 => x"82",
          2278 => x"aa",
          2279 => x"84",
          2280 => x"3f",
          2281 => x"29",
          2282 => x"98",
          2283 => x"85",
          2284 => x"3f",
          2285 => x"02",
          2286 => x"84",
          2287 => x"b8",
          2288 => x"cd",
          2289 => x"51",
          2290 => x"39",
          2291 => x"cd",
          2292 => x"51",
          2293 => x"04",
          2294 => x"87",
          2295 => x"8c",
          2296 => x"fd",
          2297 => x"2c",
          2298 => x"10",
          2299 => x"54",
          2300 => x"12",
          2301 => x"38",
          2302 => x"84",
          2303 => x"52",
          2304 => x"83",
          2305 => x"0c",
          2306 => x"79",
          2307 => x"33",
          2308 => x"38",
          2309 => x"ff",
          2310 => x"52",
          2311 => x"fb",
          2312 => x"a3",
          2313 => x"74",
          2314 => x"39",
          2315 => x"74",
          2316 => x"0d",
          2317 => x"02",
          2318 => x"e8",
          2319 => x"05",
          2320 => x"59",
          2321 => x"9a",
          2322 => x"84",
          2323 => x"70",
          2324 => x"82",
          2325 => x"e8",
          2326 => x"05",
          2327 => x"2e",
          2328 => x"51",
          2329 => x"33",
          2330 => x"34",
          2331 => x"27",
          2332 => x"34",
          2333 => x"e4",
          2334 => x"82",
          2335 => x"8c",
          2336 => x"52",
          2337 => x"df",
          2338 => x"d6",
          2339 => x"ef",
          2340 => x"3d",
          2341 => x"72",
          2342 => x"71",
          2343 => x"ff",
          2344 => x"25",
          2345 => x"34",
          2346 => x"2e",
          2347 => x"3f",
          2348 => x"3f",
          2349 => x"3d",
          2350 => x"80",
          2351 => x"f5",
          2352 => x"d3",
          2353 => x"f8",
          2354 => x"9f",
          2355 => x"2e",
          2356 => x"3f",
          2357 => x"82",
          2358 => x"e0",
          2359 => x"55",
          2360 => x"81",
          2361 => x"80",
          2362 => x"06",
          2363 => x"d9",
          2364 => x"08",
          2365 => x"52",
          2366 => x"f2",
          2367 => x"38",
          2368 => x"55",
          2369 => x"56",
          2370 => x"08",
          2371 => x"a8",
          2372 => x"18",
          2373 => x"08",
          2374 => x"ff",
          2375 => x"34",
          2376 => x"9f",
          2377 => x"85",
          2378 => x"e4",
          2379 => x"f4",
          2380 => x"2e",
          2381 => x"ff",
          2382 => x"06",
          2383 => x"a8",
          2384 => x"3f",
          2385 => x"08",
          2386 => x"98",
          2387 => x"0d",
          2388 => x"57",
          2389 => x"81",
          2390 => x"56",
          2391 => x"70",
          2392 => x"73",
          2393 => x"75",
          2394 => x"88",
          2395 => x"52",
          2396 => x"98",
          2397 => x"ff",
          2398 => x"80",
          2399 => x"81",
          2400 => x"38",
          2401 => x"81",
          2402 => x"f8",
          2403 => x"98",
          2404 => x"53",
          2405 => x"82",
          2406 => x"74",
          2407 => x"14",
          2408 => x"74",
          2409 => x"82",
          2410 => x"d3",
          2411 => x"08",
          2412 => x"0b",
          2413 => x"82",
          2414 => x"cb",
          2415 => x"55",
          2416 => x"2e",
          2417 => x"55",
          2418 => x"a8",
          2419 => x"08",
          2420 => x"08",
          2421 => x"76",
          2422 => x"de",
          2423 => x"2e",
          2424 => x"98",
          2425 => x"98",
          2426 => x"80",
          2427 => x"81",
          2428 => x"56",
          2429 => x"81",
          2430 => x"08",
          2431 => x"98",
          2432 => x"08",
          2433 => x"ff",
          2434 => x"34",
          2435 => x"75",
          2436 => x"81",
          2437 => x"83",
          2438 => x"81",
          2439 => x"82",
          2440 => x"df",
          2441 => x"d6",
          2442 => x"a3",
          2443 => x"70",
          2444 => x"ec",
          2445 => x"d4",
          2446 => x"82",
          2447 => x"97",
          2448 => x"29",
          2449 => x"70",
          2450 => x"51",
          2451 => x"2e",
          2452 => x"38",
          2453 => x"0a",
          2454 => x"75",
          2455 => x"52",
          2456 => x"98",
          2457 => x"2e",
          2458 => x"81",
          2459 => x"29",
          2460 => x"70",
          2461 => x"95",
          2462 => x"77",
          2463 => x"08",
          2464 => x"d3",
          2465 => x"ca",
          2466 => x"d4",
          2467 => x"82",
          2468 => x"98",
          2469 => x"82",
          2470 => x"51",
          2471 => x"09",
          2472 => x"f0",
          2473 => x"f7",
          2474 => x"34",
          2475 => x"75",
          2476 => x"34",
          2477 => x"26",
          2478 => x"b8",
          2479 => x"f7",
          2480 => x"c9",
          2481 => x"75",
          2482 => x"98",
          2483 => x"38",
          2484 => x"34",
          2485 => x"0a",
          2486 => x"33",
          2487 => x"dc",
          2488 => x"f7",
          2489 => x"33",
          2490 => x"73",
          2491 => x"73",
          2492 => x"33",
          2493 => x"0a",
          2494 => x"33",
          2495 => x"a8",
          2496 => x"1a",
          2497 => x"3f",
          2498 => x"0a",
          2499 => x"33",
          2500 => x"38",
          2501 => x"70",
          2502 => x"51",
          2503 => x"38",
          2504 => x"ff",
          2505 => x"29",
          2506 => x"82",
          2507 => x"75",
          2508 => x"7a",
          2509 => x"f7",
          2510 => x"51",
          2511 => x"f7",
          2512 => x"55",
          2513 => x"f7",
          2514 => x"f7",
          2515 => x"f7",
          2516 => x"88",
          2517 => x"dc",
          2518 => x"82",
          2519 => x"74",
          2520 => x"81",
          2521 => x"08",
          2522 => x"3f",
          2523 => x"0a",
          2524 => x"33",
          2525 => x"38",
          2526 => x"ff",
          2527 => x"70",
          2528 => x"d8",
          2529 => x"24",
          2530 => x"52",
          2531 => x"81",
          2532 => x"70",
          2533 => x"51",
          2534 => x"99",
          2535 => x"54",
          2536 => x"52",
          2537 => x"f7",
          2538 => x"82",
          2539 => x"73",
          2540 => x"73",
          2541 => x"52",
          2542 => x"80",
          2543 => x"34",
          2544 => x"82",
          2545 => x"82",
          2546 => x"f9",
          2547 => x"88",
          2548 => x"dc",
          2549 => x"dc",
          2550 => x"39",
          2551 => x"33",
          2552 => x"38",
          2553 => x"34",
          2554 => x"81",
          2555 => x"25",
          2556 => x"33",
          2557 => x"73",
          2558 => x"81",
          2559 => x"70",
          2560 => x"51",
          2561 => x"fb",
          2562 => x"d3",
          2563 => x"2b",
          2564 => x"57",
          2565 => x"a1",
          2566 => x"51",
          2567 => x"0a",
          2568 => x"2c",
          2569 => x"75",
          2570 => x"82",
          2571 => x"82",
          2572 => x"77",
          2573 => x"08",
          2574 => x"dc",
          2575 => x"ff",
          2576 => x"70",
          2577 => x"58",
          2578 => x"f7",
          2579 => x"52",
          2580 => x"80",
          2581 => x"82",
          2582 => x"b0",
          2583 => x"80",
          2584 => x"f6",
          2585 => x"d8",
          2586 => x"06",
          2587 => x"ff",
          2588 => x"39",
          2589 => x"fc",
          2590 => x"a7",
          2591 => x"82",
          2592 => x"82",
          2593 => x"05",
          2594 => x"86",
          2595 => x"73",
          2596 => x"38",
          2597 => x"39",
          2598 => x"38",
          2599 => x"2e",
          2600 => x"3f",
          2601 => x"34",
          2602 => x"81",
          2603 => x"9b",
          2604 => x"29",
          2605 => x"54",
          2606 => x"ff",
          2607 => x"82",
          2608 => x"81",
          2609 => x"79",
          2610 => x"54",
          2611 => x"74",
          2612 => x"82",
          2613 => x"52",
          2614 => x"39",
          2615 => x"06",
          2616 => x"74",
          2617 => x"fc",
          2618 => x"f7",
          2619 => x"54",
          2620 => x"82",
          2621 => x"f4",
          2622 => x"88",
          2623 => x"dc",
          2624 => x"dc",
          2625 => x"84",
          2626 => x"a0",
          2627 => x"80",
          2628 => x"51",
          2629 => x"08",
          2630 => x"57",
          2631 => x"08",
          2632 => x"15",
          2633 => x"86",
          2634 => x"e0",
          2635 => x"05",
          2636 => x"ff",
          2637 => x"56",
          2638 => x"34",
          2639 => x"82",
          2640 => x"55",
          2641 => x"15",
          2642 => x"0d",
          2643 => x"8f",
          2644 => x"70",
          2645 => x"70",
          2646 => x"04",
          2647 => x"02",
          2648 => x"82",
          2649 => x"11",
          2650 => x"81",
          2651 => x"a4",
          2652 => x"ff",
          2653 => x"52",
          2654 => x"55",
          2655 => x"82",
          2656 => x"52",
          2657 => x"15",
          2658 => x"70",
          2659 => x"07",
          2660 => x"51",
          2661 => x"ff",
          2662 => x"51",
          2663 => x"06",
          2664 => x"88",
          2665 => x"81",
          2666 => x"3d",
          2667 => x"05",
          2668 => x"11",
          2669 => x"8b",
          2670 => x"59",
          2671 => x"33",
          2672 => x"70",
          2673 => x"84",
          2674 => x"e0",
          2675 => x"85",
          2676 => x"2b",
          2677 => x"86",
          2678 => x"2b",
          2679 => x"52",
          2680 => x"34",
          2681 => x"81",
          2682 => x"81",
          2683 => x"51",
          2684 => x"81",
          2685 => x"3d",
          2686 => x"88",
          2687 => x"33",
          2688 => x"70",
          2689 => x"33",
          2690 => x"53",
          2691 => x"53",
          2692 => x"72",
          2693 => x"08",
          2694 => x"71",
          2695 => x"11",
          2696 => x"2b",
          2697 => x"06",
          2698 => x"53",
          2699 => x"72",
          2700 => x"82",
          2701 => x"81",
          2702 => x"2b",
          2703 => x"70",
          2704 => x"07",
          2705 => x"2a",
          2706 => x"34",
          2707 => x"04",
          2708 => x"02",
          2709 => x"2b",
          2710 => x"33",
          2711 => x"59",
          2712 => x"71",
          2713 => x"07",
          2714 => x"07",
          2715 => x"53",
          2716 => x"82",
          2717 => x"81",
          2718 => x"2b",
          2719 => x"82",
          2720 => x"2b",
          2721 => x"52",
          2722 => x"34",
          2723 => x"33",
          2724 => x"82",
          2725 => x"0d",
          2726 => x"88",
          2727 => x"ff",
          2728 => x"3f",
          2729 => x"71",
          2730 => x"71",
          2731 => x"11",
          2732 => x"2b",
          2733 => x"51",
          2734 => x"80",
          2735 => x"75",
          2736 => x"84",
          2737 => x"2b",
          2738 => x"88",
          2739 => x"86",
          2740 => x"75",
          2741 => x"70",
          2742 => x"71",
          2743 => x"57",
          2744 => x"73",
          2745 => x"18",
          2746 => x"0b",
          2747 => x"53",
          2748 => x"34",
          2749 => x"81",
          2750 => x"82",
          2751 => x"51",
          2752 => x"81",
          2753 => x"3d",
          2754 => x"84",
          2755 => x"86",
          2756 => x"3d",
          2757 => x"52",
          2758 => x"08",
          2759 => x"08",
          2760 => x"88",
          2761 => x"5a",
          2762 => x"80",
          2763 => x"33",
          2764 => x"70",
          2765 => x"83",
          2766 => x"53",
          2767 => x"8a",
          2768 => x"78",
          2769 => x"33",
          2770 => x"c2",
          2771 => x"38",
          2772 => x"2b",
          2773 => x"81",
          2774 => x"81",
          2775 => x"5c",
          2776 => x"55",
          2777 => x"38",
          2778 => x"38",
          2779 => x"38",
          2780 => x"39",
          2781 => x"51",
          2782 => x"70",
          2783 => x"71",
          2784 => x"5a",
          2785 => x"83",
          2786 => x"59",
          2787 => x"81",
          2788 => x"82",
          2789 => x"11",
          2790 => x"33",
          2791 => x"53",
          2792 => x"86",
          2793 => x"e0",
          2794 => x"85",
          2795 => x"2b",
          2796 => x"54",
          2797 => x"34",
          2798 => x"1d",
          2799 => x"88",
          2800 => x"5f",
          2801 => x"75",
          2802 => x"1b",
          2803 => x"0c",
          2804 => x"74",
          2805 => x"f4",
          2806 => x"8b",
          2807 => x"e0",
          2808 => x"0c",
          2809 => x"64",
          2810 => x"82",
          2811 => x"06",
          2812 => x"38",
          2813 => x"98",
          2814 => x"38",
          2815 => x"83",
          2816 => x"82",
          2817 => x"82",
          2818 => x"2a",
          2819 => x"2b",
          2820 => x"71",
          2821 => x"83",
          2822 => x"05",
          2823 => x"12",
          2824 => x"2b",
          2825 => x"5c",
          2826 => x"73",
          2827 => x"ff",
          2828 => x"06",
          2829 => x"33",
          2830 => x"1c",
          2831 => x"2b",
          2832 => x"52",
          2833 => x"78",
          2834 => x"41",
          2835 => x"60",
          2836 => x"06",
          2837 => x"7a",
          2838 => x"39",
          2839 => x"38",
          2840 => x"39",
          2841 => x"c8",
          2842 => x"12",
          2843 => x"54",
          2844 => x"f7",
          2845 => x"ff",
          2846 => x"83",
          2847 => x"05",
          2848 => x"82",
          2849 => x"83",
          2850 => x"39",
          2851 => x"d4",
          2852 => x"e0",
          2853 => x"12",
          2854 => x"54",
          2855 => x"f6",
          2856 => x"ff",
          2857 => x"83",
          2858 => x"05",
          2859 => x"82",
          2860 => x"62",
          2861 => x"ff",
          2862 => x"54",
          2863 => x"5c",
          2864 => x"38",
          2865 => x"08",
          2866 => x"f7",
          2867 => x"99",
          2868 => x"f2",
          2869 => x"e0",
          2870 => x"f9",
          2871 => x"0c",
          2872 => x"77",
          2873 => x"3f",
          2874 => x"98",
          2875 => x"80",
          2876 => x"90",
          2877 => x"86",
          2878 => x"8f",
          2879 => x"26",
          2880 => x"52",
          2881 => x"0d",
          2882 => x"33",
          2883 => x"53",
          2884 => x"38",
          2885 => x"11",
          2886 => x"84",
          2887 => x"87",
          2888 => x"0c",
          2889 => x"70",
          2890 => x"51",
          2891 => x"98",
          2892 => x"08",
          2893 => x"38",
          2894 => x"80",
          2895 => x"14",
          2896 => x"70",
          2897 => x"04",
          2898 => x"8c",
          2899 => x"5b",
          2900 => x"82",
          2901 => x"52",
          2902 => x"84",
          2903 => x"c0",
          2904 => x"13",
          2905 => x"0b",
          2906 => x"0c",
          2907 => x"2a",
          2908 => x"80",
          2909 => x"7b",
          2910 => x"59",
          2911 => x"73",
          2912 => x"ff",
          2913 => x"38",
          2914 => x"c3",
          2915 => x"71",
          2916 => x"2e",
          2917 => x"92",
          2918 => x"06",
          2919 => x"5a",
          2920 => x"70",
          2921 => x"80",
          2922 => x"06",
          2923 => x"fe",
          2924 => x"52",
          2925 => x"71",
          2926 => x"3d",
          2927 => x"64",
          2928 => x"40",
          2929 => x"58",
          2930 => x"81",
          2931 => x"09",
          2932 => x"84",
          2933 => x"c0",
          2934 => x"13",
          2935 => x"87",
          2936 => x"82",
          2937 => x"84",
          2938 => x"71",
          2939 => x"05",
          2940 => x"73",
          2941 => x"71",
          2942 => x"8c",
          2943 => x"98",
          2944 => x"38",
          2945 => x"76",
          2946 => x"72",
          2947 => x"f7",
          2948 => x"1a",
          2949 => x"59",
          2950 => x"73",
          2951 => x"38",
          2952 => x"fc",
          2953 => x"83",
          2954 => x"e0",
          2955 => x"3d",
          2956 => x"33",
          2957 => x"54",
          2958 => x"e0",
          2959 => x"72",
          2960 => x"98",
          2961 => x"80",
          2962 => x"74",
          2963 => x"54",
          2964 => x"d4",
          2965 => x"80",
          2966 => x"70",
          2967 => x"2e",
          2968 => x"52",
          2969 => x"08",
          2970 => x"87",
          2971 => x"70",
          2972 => x"96",
          2973 => x"0a",
          2974 => x"0c",
          2975 => x"54",
          2976 => x"0d",
          2977 => x"33",
          2978 => x"e0",
          2979 => x"04",
          2980 => x"82",
          2981 => x"2b",
          2982 => x"88",
          2983 => x"98",
          2984 => x"85",
          2985 => x"02",
          2986 => x"70",
          2987 => x"88",
          2988 => x"0d",
          2989 => x"52",
          2990 => x"70",
          2991 => x"05",
          2992 => x"72",
          2993 => x"2a",
          2994 => x"04",
          2995 => x"54",
          2996 => x"70",
          2997 => x"05",
          2998 => x"84",
          2999 => x"77",
          3000 => x"81",
          3001 => x"f4",
          3002 => x"0d",
          3003 => x"70",
          3004 => x"05",
          3005 => x"56",
          3006 => x"38",
          3007 => x"e0",
          3008 => x"3d",
          3009 => x"71",
          3010 => x"70",
          3011 => x"82",
          3012 => x"80",
          3013 => x"3d",
          3014 => x"05",
          3015 => x"e7",
          3016 => x"a2",
          3017 => x"b5",
          3018 => x"82",
          3019 => x"53",
          3020 => x"0c",
          3021 => x"87",
          3022 => x"56",
          3023 => x"74",
          3024 => x"b4",
          3025 => x"81",
          3026 => x"82",
          3027 => x"06",
          3028 => x"17",
          3029 => x"08",
          3030 => x"74",
          3031 => x"55",
          3032 => x"38",
          3033 => x"81",
          3034 => x"39",
          3035 => x"8b",
          3036 => x"7a",
          3037 => x"08",
          3038 => x"3f",
          3039 => x"98",
          3040 => x"b8",
          3041 => x"80",
          3042 => x"85",
          3043 => x"17",
          3044 => x"3d",
          3045 => x"52",
          3046 => x"08",
          3047 => x"38",
          3048 => x"81",
          3049 => x"59",
          3050 => x"e3",
          3051 => x"08",
          3052 => x"d3",
          3053 => x"17",
          3054 => x"a4",
          3055 => x"86",
          3056 => x"17",
          3057 => x"52",
          3058 => x"90",
          3059 => x"fb",
          3060 => x"70",
          3061 => x"52",
          3062 => x"77",
          3063 => x"81",
          3064 => x"e0",
          3065 => x"58",
          3066 => x"0d",
          3067 => x"9c",
          3068 => x"80",
          3069 => x"14",
          3070 => x"05",
          3071 => x"87",
          3072 => x"7a",
          3073 => x"27",
          3074 => x"27",
          3075 => x"58",
          3076 => x"82",
          3077 => x"38",
          3078 => x"8e",
          3079 => x"17",
          3080 => x"53",
          3081 => x"e0",
          3082 => x"ff",
          3083 => x"70",
          3084 => x"76",
          3085 => x"82",
          3086 => x"83",
          3087 => x"88",
          3088 => x"84",
          3089 => x"80",
          3090 => x"80",
          3091 => x"08",
          3092 => x"82",
          3093 => x"10",
          3094 => x"51",
          3095 => x"83",
          3096 => x"87",
          3097 => x"51",
          3098 => x"9b",
          3099 => x"74",
          3100 => x"82",
          3101 => x"83",
          3102 => x"0c",
          3103 => x"7a",
          3104 => x"81",
          3105 => x"17",
          3106 => x"53",
          3107 => x"79",
          3108 => x"38",
          3109 => x"b8",
          3110 => x"17",
          3111 => x"53",
          3112 => x"e0",
          3113 => x"81",
          3114 => x"b8",
          3115 => x"56",
          3116 => x"38",
          3117 => x"33",
          3118 => x"74",
          3119 => x"89",
          3120 => x"51",
          3121 => x"59",
          3122 => x"74",
          3123 => x"84",
          3124 => x"88",
          3125 => x"8f",
          3126 => x"80",
          3127 => x"08",
          3128 => x"82",
          3129 => x"08",
          3130 => x"06",
          3131 => x"05",
          3132 => x"39",
          3133 => x"52",
          3134 => x"98",
          3135 => x"38",
          3136 => x"83",
          3137 => x"54",
          3138 => x"e0",
          3139 => x"52",
          3140 => x"83",
          3141 => x"8a",
          3142 => x"7c",
          3143 => x"81",
          3144 => x"08",
          3145 => x"38",
          3146 => x"a4",
          3147 => x"e0",
          3148 => x"82",
          3149 => x"e6",
          3150 => x"de",
          3151 => x"3f",
          3152 => x"98",
          3153 => x"e0",
          3154 => x"e0",
          3155 => x"53",
          3156 => x"82",
          3157 => x"08",
          3158 => x"57",
          3159 => x"94",
          3160 => x"54",
          3161 => x"78",
          3162 => x"82",
          3163 => x"f6",
          3164 => x"5b",
          3165 => x"58",
          3166 => x"08",
          3167 => x"39",
          3168 => x"81",
          3169 => x"82",
          3170 => x"82",
          3171 => x"38",
          3172 => x"26",
          3173 => x"08",
          3174 => x"b9",
          3175 => x"80",
          3176 => x"08",
          3177 => x"52",
          3178 => x"82",
          3179 => x"06",
          3180 => x"82",
          3181 => x"72",
          3182 => x"e0",
          3183 => x"73",
          3184 => x"80",
          3185 => x"81",
          3186 => x"08",
          3187 => x"75",
          3188 => x"56",
          3189 => x"82",
          3190 => x"75",
          3191 => x"e0",
          3192 => x"59",
          3193 => x"81",
          3194 => x"59",
          3195 => x"70",
          3196 => x"51",
          3197 => x"75",
          3198 => x"38",
          3199 => x"75",
          3200 => x"e0",
          3201 => x"70",
          3202 => x"51",
          3203 => x"73",
          3204 => x"52",
          3205 => x"98",
          3206 => x"18",
          3207 => x"18",
          3208 => x"38",
          3209 => x"33",
          3210 => x"97",
          3211 => x"38",
          3212 => x"e0",
          3213 => x"75",
          3214 => x"3d",
          3215 => x"52",
          3216 => x"08",
          3217 => x"80",
          3218 => x"c1",
          3219 => x"98",
          3220 => x"53",
          3221 => x"f2",
          3222 => x"16",
          3223 => x"27",
          3224 => x"76",
          3225 => x"3f",
          3226 => x"38",
          3227 => x"70",
          3228 => x"56",
          3229 => x"3d",
          3230 => x"71",
          3231 => x"0a",
          3232 => x"53",
          3233 => x"0c",
          3234 => x"75",
          3235 => x"ac",
          3236 => x"85",
          3237 => x"5a",
          3238 => x"ac",
          3239 => x"39",
          3240 => x"58",
          3241 => x"76",
          3242 => x"08",
          3243 => x"bd",
          3244 => x"27",
          3245 => x"98",
          3246 => x"39",
          3247 => x"52",
          3248 => x"98",
          3249 => x"0c",
          3250 => x"80",
          3251 => x"94",
          3252 => x"0c",
          3253 => x"9c",
          3254 => x"98",
          3255 => x"0d",
          3256 => x"05",
          3257 => x"27",
          3258 => x"98",
          3259 => x"2e",
          3260 => x"58",
          3261 => x"15",
          3262 => x"38",
          3263 => x"53",
          3264 => x"c0",
          3265 => x"89",
          3266 => x"74",
          3267 => x"e0",
          3268 => x"82",
          3269 => x"81",
          3270 => x"80",
          3271 => x"98",
          3272 => x"38",
          3273 => x"dd",
          3274 => x"f9",
          3275 => x"87",
          3276 => x"80",
          3277 => x"08",
          3278 => x"e0",
          3279 => x"e0",
          3280 => x"3f",
          3281 => x"94",
          3282 => x"c1",
          3283 => x"0c",
          3284 => x"05",
          3285 => x"e0",
          3286 => x"3d",
          3287 => x"57",
          3288 => x"82",
          3289 => x"08",
          3290 => x"56",
          3291 => x"83",
          3292 => x"e0",
          3293 => x"98",
          3294 => x"54",
          3295 => x"06",
          3296 => x"08",
          3297 => x"75",
          3298 => x"81",
          3299 => x"06",
          3300 => x"08",
          3301 => x"3f",
          3302 => x"98",
          3303 => x"84",
          3304 => x"54",
          3305 => x"0d",
          3306 => x"52",
          3307 => x"08",
          3308 => x"51",
          3309 => x"06",
          3310 => x"3f",
          3311 => x"07",
          3312 => x"3d",
          3313 => x"70",
          3314 => x"53",
          3315 => x"33",
          3316 => x"06",
          3317 => x"15",
          3318 => x"04",
          3319 => x"8b",
          3320 => x"29",
          3321 => x"71",
          3322 => x"56",
          3323 => x"82",
          3324 => x"f2",
          3325 => x"79",
          3326 => x"5d",
          3327 => x"38",
          3328 => x"db",
          3329 => x"e0",
          3330 => x"08",
          3331 => x"84",
          3332 => x"bf",
          3333 => x"72",
          3334 => x"56",
          3335 => x"83",
          3336 => x"53",
          3337 => x"38",
          3338 => x"99",
          3339 => x"06",
          3340 => x"06",
          3341 => x"87",
          3342 => x"76",
          3343 => x"38",
          3344 => x"53",
          3345 => x"33",
          3346 => x"08",
          3347 => x"7c",
          3348 => x"8d",
          3349 => x"81",
          3350 => x"9a",
          3351 => x"e0",
          3352 => x"72",
          3353 => x"bf",
          3354 => x"81",
          3355 => x"33",
          3356 => x"e0",
          3357 => x"77",
          3358 => x"26",
          3359 => x"59",
          3360 => x"8b",
          3361 => x"81",
          3362 => x"77",
          3363 => x"2a",
          3364 => x"80",
          3365 => x"92",
          3366 => x"23",
          3367 => x"53",
          3368 => x"9d",
          3369 => x"e8",
          3370 => x"06",
          3371 => x"0b",
          3372 => x"78",
          3373 => x"08",
          3374 => x"98",
          3375 => x"80",
          3376 => x"98",
          3377 => x"0d",
          3378 => x"78",
          3379 => x"08",
          3380 => x"38",
          3381 => x"ac",
          3382 => x"51",
          3383 => x"58",
          3384 => x"9c",
          3385 => x"86",
          3386 => x"17",
          3387 => x"56",
          3388 => x"e5",
          3389 => x"70",
          3390 => x"8e",
          3391 => x"2e",
          3392 => x"19",
          3393 => x"51",
          3394 => x"86",
          3395 => x"80",
          3396 => x"81",
          3397 => x"1d",
          3398 => x"09",
          3399 => x"33",
          3400 => x"81",
          3401 => x"52",
          3402 => x"08",
          3403 => x"95",
          3404 => x"29",
          3405 => x"5a",
          3406 => x"51",
          3407 => x"83",
          3408 => x"b1",
          3409 => x"38",
          3410 => x"e0",
          3411 => x"53",
          3412 => x"8d",
          3413 => x"09",
          3414 => x"8b",
          3415 => x"81",
          3416 => x"7b",
          3417 => x"86",
          3418 => x"79",
          3419 => x"8b",
          3420 => x"54",
          3421 => x"ff",
          3422 => x"54",
          3423 => x"76",
          3424 => x"08",
          3425 => x"bb",
          3426 => x"73",
          3427 => x"9c",
          3428 => x"e0",
          3429 => x"ff",
          3430 => x"52",
          3431 => x"98",
          3432 => x"2e",
          3433 => x"0c",
          3434 => x"64",
          3435 => x"06",
          3436 => x"b5",
          3437 => x"56",
          3438 => x"81",
          3439 => x"55",
          3440 => x"70",
          3441 => x"e4",
          3442 => x"81",
          3443 => x"38",
          3444 => x"5b",
          3445 => x"53",
          3446 => x"85",
          3447 => x"77",
          3448 => x"55",
          3449 => x"ff",
          3450 => x"57",
          3451 => x"81",
          3452 => x"51",
          3453 => x"38",
          3454 => x"17",
          3455 => x"39",
          3456 => x"05",
          3457 => x"54",
          3458 => x"54",
          3459 => x"76",
          3460 => x"38",
          3461 => x"fe",
          3462 => x"78",
          3463 => x"74",
          3464 => x"3f",
          3465 => x"38",
          3466 => x"38",
          3467 => x"77",
          3468 => x"51",
          3469 => x"eb",
          3470 => x"58",
          3471 => x"81",
          3472 => x"57",
          3473 => x"38",
          3474 => x"98",
          3475 => x"e3",
          3476 => x"7a",
          3477 => x"e0",
          3478 => x"84",
          3479 => x"02",
          3480 => x"02",
          3481 => x"70",
          3482 => x"73",
          3483 => x"1d",
          3484 => x"98",
          3485 => x"f3",
          3486 => x"82",
          3487 => x"19",
          3488 => x"78",
          3489 => x"53",
          3490 => x"e0",
          3491 => x"81",
          3492 => x"3f",
          3493 => x"5d",
          3494 => x"ab",
          3495 => x"e0",
          3496 => x"08",
          3497 => x"5a",
          3498 => x"0b",
          3499 => x"8c",
          3500 => x"9a",
          3501 => x"29",
          3502 => x"ff",
          3503 => x"70",
          3504 => x"52",
          3505 => x"51",
          3506 => x"ff",
          3507 => x"27",
          3508 => x"8b",
          3509 => x"54",
          3510 => x"58",
          3511 => x"34",
          3512 => x"82",
          3513 => x"08",
          3514 => x"fe",
          3515 => x"51",
          3516 => x"57",
          3517 => x"53",
          3518 => x"08",
          3519 => x"1a",
          3520 => x"3f",
          3521 => x"06",
          3522 => x"0b",
          3523 => x"e0",
          3524 => x"3d",
          3525 => x"ac",
          3526 => x"ff",
          3527 => x"ed",
          3528 => x"82",
          3529 => x"15",
          3530 => x"82",
          3531 => x"08",
          3532 => x"73",
          3533 => x"15",
          3534 => x"98",
          3535 => x"82",
          3536 => x"08",
          3537 => x"09",
          3538 => x"82",
          3539 => x"f4",
          3540 => x"59",
          3541 => x"1c",
          3542 => x"1c",
          3543 => x"70",
          3544 => x"57",
          3545 => x"81",
          3546 => x"81",
          3547 => x"80",
          3548 => x"06",
          3549 => x"38",
          3550 => x"96",
          3551 => x"54",
          3552 => x"07",
          3553 => x"98",
          3554 => x"ff",
          3555 => x"a5",
          3556 => x"34",
          3557 => x"39",
          3558 => x"80",
          3559 => x"54",
          3560 => x"9a",
          3561 => x"17",
          3562 => x"10",
          3563 => x"fe",
          3564 => x"70",
          3565 => x"17",
          3566 => x"34",
          3567 => x"9c",
          3568 => x"5b",
          3569 => x"74",
          3570 => x"81",
          3571 => x"70",
          3572 => x"76",
          3573 => x"8b",
          3574 => x"34",
          3575 => x"05",
          3576 => x"27",
          3577 => x"53",
          3578 => x"33",
          3579 => x"38",
          3580 => x"80",
          3581 => x"55",
          3582 => x"38",
          3583 => x"33",
          3584 => x"26",
          3585 => x"33",
          3586 => x"72",
          3587 => x"2a",
          3588 => x"2e",
          3589 => x"ff",
          3590 => x"05",
          3591 => x"19",
          3592 => x"ff",
          3593 => x"80",
          3594 => x"8c",
          3595 => x"72",
          3596 => x"8b",
          3597 => x"08",
          3598 => x"82",
          3599 => x"51",
          3600 => x"86",
          3601 => x"3f",
          3602 => x"8e",
          3603 => x"70",
          3604 => x"51",
          3605 => x"81",
          3606 => x"74",
          3607 => x"08",
          3608 => x"44",
          3609 => x"73",
          3610 => x"81",
          3611 => x"70",
          3612 => x"73",
          3613 => x"70",
          3614 => x"38",
          3615 => x"52",
          3616 => x"98",
          3617 => x"7d",
          3618 => x"59",
          3619 => x"3f",
          3620 => x"b1",
          3621 => x"98",
          3622 => x"82",
          3623 => x"73",
          3624 => x"98",
          3625 => x"32",
          3626 => x"25",
          3627 => x"38",
          3628 => x"80",
          3629 => x"d1",
          3630 => x"98",
          3631 => x"26",
          3632 => x"75",
          3633 => x"39",
          3634 => x"56",
          3635 => x"06",
          3636 => x"32",
          3637 => x"51",
          3638 => x"9f",
          3639 => x"2e",
          3640 => x"54",
          3641 => x"39",
          3642 => x"c9",
          3643 => x"2e",
          3644 => x"22",
          3645 => x"b6",
          3646 => x"23",
          3647 => x"54",
          3648 => x"73",
          3649 => x"18",
          3650 => x"a0",
          3651 => x"c4",
          3652 => x"10",
          3653 => x"16",
          3654 => x"9f",
          3655 => x"75",
          3656 => x"ff",
          3657 => x"7a",
          3658 => x"8d",
          3659 => x"83",
          3660 => x"22",
          3661 => x"5d",
          3662 => x"38",
          3663 => x"51",
          3664 => x"7c",
          3665 => x"54",
          3666 => x"38",
          3667 => x"aa",
          3668 => x"51",
          3669 => x"10",
          3670 => x"78",
          3671 => x"22",
          3672 => x"06",
          3673 => x"1e",
          3674 => x"5c",
          3675 => x"81",
          3676 => x"82",
          3677 => x"75",
          3678 => x"51",
          3679 => x"73",
          3680 => x"57",
          3681 => x"78",
          3682 => x"32",
          3683 => x"70",
          3684 => x"80",
          3685 => x"ae",
          3686 => x"83",
          3687 => x"38",
          3688 => x"2b",
          3689 => x"39",
          3690 => x"82",
          3691 => x"80",
          3692 => x"83",
          3693 => x"81",
          3694 => x"8c",
          3695 => x"b8",
          3696 => x"27",
          3697 => x"26",
          3698 => x"57",
          3699 => x"76",
          3700 => x"81",
          3701 => x"2e",
          3702 => x"51",
          3703 => x"80",
          3704 => x"07",
          3705 => x"54",
          3706 => x"07",
          3707 => x"26",
          3708 => x"70",
          3709 => x"7d",
          3710 => x"81",
          3711 => x"33",
          3712 => x"06",
          3713 => x"7e",
          3714 => x"7b",
          3715 => x"8c",
          3716 => x"7b",
          3717 => x"81",
          3718 => x"76",
          3719 => x"73",
          3720 => x"80",
          3721 => x"7b",
          3722 => x"73",
          3723 => x"57",
          3724 => x"a5",
          3725 => x"33",
          3726 => x"2e",
          3727 => x"2e",
          3728 => x"85",
          3729 => x"57",
          3730 => x"74",
          3731 => x"ed",
          3732 => x"80",
          3733 => x"54",
          3734 => x"74",
          3735 => x"73",
          3736 => x"2a",
          3737 => x"80",
          3738 => x"ff",
          3739 => x"51",
          3740 => x"88",
          3741 => x"e0",
          3742 => x"3d",
          3743 => x"71",
          3744 => x"80",
          3745 => x"05",
          3746 => x"71",
          3747 => x"71",
          3748 => x"38",
          3749 => x"06",
          3750 => x"38",
          3751 => x"05",
          3752 => x"38",
          3753 => x"77",
          3754 => x"05",
          3755 => x"33",
          3756 => x"99",
          3757 => x"ff",
          3758 => x"70",
          3759 => x"81",
          3760 => x"9f",
          3761 => x"81",
          3762 => x"72",
          3763 => x"72",
          3764 => x"53",
          3765 => x"38",
          3766 => x"75",
          3767 => x"83",
          3768 => x"59",
          3769 => x"33",
          3770 => x"3d",
          3771 => x"80",
          3772 => x"17",
          3773 => x"3f",
          3774 => x"80",
          3775 => x"3f",
          3776 => x"06",
          3777 => x"2e",
          3778 => x"0b",
          3779 => x"e9",
          3780 => x"57",
          3781 => x"80",
          3782 => x"8a",
          3783 => x"06",
          3784 => x"52",
          3785 => x"82",
          3786 => x"08",
          3787 => x"d1",
          3788 => x"ed",
          3789 => x"e0",
          3790 => x"55",
          3791 => x"0d",
          3792 => x"05",
          3793 => x"75",
          3794 => x"e0",
          3795 => x"82",
          3796 => x"82",
          3797 => x"e0",
          3798 => x"73",
          3799 => x"0c",
          3800 => x"57",
          3801 => x"33",
          3802 => x"08",
          3803 => x"55",
          3804 => x"83",
          3805 => x"51",
          3806 => x"86",
          3807 => x"59",
          3808 => x"34",
          3809 => x"81",
          3810 => x"06",
          3811 => x"72",
          3812 => x"38",
          3813 => x"53",
          3814 => x"70",
          3815 => x"82",
          3816 => x"76",
          3817 => x"81",
          3818 => x"53",
          3819 => x"3d",
          3820 => x"15",
          3821 => x"8d",
          3822 => x"3f",
          3823 => x"70",
          3824 => x"16",
          3825 => x"77",
          3826 => x"30",
          3827 => x"3d",
          3828 => x"53",
          3829 => x"83",
          3830 => x"52",
          3831 => x"98",
          3832 => x"82",
          3833 => x"78",
          3834 => x"58",
          3835 => x"2e",
          3836 => x"56",
          3837 => x"76",
          3838 => x"76",
          3839 => x"14",
          3840 => x"08",
          3841 => x"80",
          3842 => x"80",
          3843 => x"e0",
          3844 => x"77",
          3845 => x"f0",
          3846 => x"a0",
          3847 => x"15",
          3848 => x"70",
          3849 => x"56",
          3850 => x"81",
          3851 => x"16",
          3852 => x"23",
          3853 => x"73",
          3854 => x"8d",
          3855 => x"51",
          3856 => x"53",
          3857 => x"72",
          3858 => x"d5",
          3859 => x"3f",
          3860 => x"06",
          3861 => x"51",
          3862 => x"55",
          3863 => x"82",
          3864 => x"53",
          3865 => x"38",
          3866 => x"2a",
          3867 => x"8d",
          3868 => x"31",
          3869 => x"98",
          3870 => x"2e",
          3871 => x"80",
          3872 => x"83",
          3873 => x"38",
          3874 => x"38",
          3875 => x"80",
          3876 => x"9c",
          3877 => x"1c",
          3878 => x"17",
          3879 => x"81",
          3880 => x"c7",
          3881 => x"ff",
          3882 => x"95",
          3883 => x"14",
          3884 => x"08",
          3885 => x"a2",
          3886 => x"f5",
          3887 => x"15",
          3888 => x"10",
          3889 => x"05",
          3890 => x"53",
          3891 => x"81",
          3892 => x"ff",
          3893 => x"84",
          3894 => x"06",
          3895 => x"c6",
          3896 => x"ff",
          3897 => x"81",
          3898 => x"73",
          3899 => x"08",
          3900 => x"84",
          3901 => x"99",
          3902 => x"ff",
          3903 => x"09",
          3904 => x"51",
          3905 => x"84",
          3906 => x"06",
          3907 => x"80",
          3908 => x"85",
          3909 => x"38",
          3910 => x"82",
          3911 => x"a4",
          3912 => x"98",
          3913 => x"82",
          3914 => x"82",
          3915 => x"82",
          3916 => x"0b",
          3917 => x"e0",
          3918 => x"3d",
          3919 => x"2e",
          3920 => x"2e",
          3921 => x"2e",
          3922 => x"22",
          3923 => x"06",
          3924 => x"be",
          3925 => x"06",
          3926 => x"54",
          3927 => x"71",
          3928 => x"87",
          3929 => x"ab",
          3930 => x"05",
          3931 => x"80",
          3932 => x"38",
          3933 => x"f7",
          3934 => x"80",
          3935 => x"54",
          3936 => x"34",
          3937 => x"2e",
          3938 => x"53",
          3939 => x"e0",
          3940 => x"0c",
          3941 => x"68",
          3942 => x"59",
          3943 => x"c8",
          3944 => x"3d",
          3945 => x"52",
          3946 => x"08",
          3947 => x"38",
          3948 => x"52",
          3949 => x"08",
          3950 => x"02",
          3951 => x"55",
          3952 => x"55",
          3953 => x"81",
          3954 => x"74",
          3955 => x"75",
          3956 => x"08",
          3957 => x"91",
          3958 => x"82",
          3959 => x"80",
          3960 => x"39",
          3961 => x"38",
          3962 => x"54",
          3963 => x"52",
          3964 => x"98",
          3965 => x"62",
          3966 => x"54",
          3967 => x"62",
          3968 => x"52",
          3969 => x"7a",
          3970 => x"80",
          3971 => x"08",
          3972 => x"3d",
          3973 => x"e0",
          3974 => x"82",
          3975 => x"38",
          3976 => x"70",
          3977 => x"2e",
          3978 => x"77",
          3979 => x"73",
          3980 => x"54",
          3981 => x"82",
          3982 => x"eb",
          3983 => x"18",
          3984 => x"98",
          3985 => x"70",
          3986 => x"86",
          3987 => x"b4",
          3988 => x"1b",
          3989 => x"a1",
          3990 => x"98",
          3991 => x"52",
          3992 => x"08",
          3993 => x"77",
          3994 => x"1a",
          3995 => x"91",
          3996 => x"80",
          3997 => x"70",
          3998 => x"81",
          3999 => x"2e",
          4000 => x"94",
          4001 => x"2b",
          4002 => x"52",
          4003 => x"98",
          4004 => x"26",
          4005 => x"08",
          4006 => x"79",
          4007 => x"70",
          4008 => x"76",
          4009 => x"55",
          4010 => x"0c",
          4011 => x"54",
          4012 => x"7a",
          4013 => x"08",
          4014 => x"89",
          4015 => x"1a",
          4016 => x"54",
          4017 => x"0d",
          4018 => x"64",
          4019 => x"90",
          4020 => x"ce",
          4021 => x"e0",
          4022 => x"55",
          4023 => x"82",
          4024 => x"55",
          4025 => x"38",
          4026 => x"82",
          4027 => x"1a",
          4028 => x"19",
          4029 => x"7c",
          4030 => x"2e",
          4031 => x"83",
          4032 => x"38",
          4033 => x"89",
          4034 => x"75",
          4035 => x"39",
          4036 => x"db",
          4037 => x"75",
          4038 => x"ff",
          4039 => x"19",
          4040 => x"82",
          4041 => x"38",
          4042 => x"2a",
          4043 => x"38",
          4044 => x"5c",
          4045 => x"7a",
          4046 => x"52",
          4047 => x"3f",
          4048 => x"7e",
          4049 => x"2e",
          4050 => x"55",
          4051 => x"53",
          4052 => x"31",
          4053 => x"e8",
          4054 => x"76",
          4055 => x"ff",
          4056 => x"7b",
          4057 => x"19",
          4058 => x"82",
          4059 => x"53",
          4060 => x"b8",
          4061 => x"3f",
          4062 => x"0c",
          4063 => x"1c",
          4064 => x"56",
          4065 => x"0d",
          4066 => x"64",
          4067 => x"90",
          4068 => x"ce",
          4069 => x"e0",
          4070 => x"55",
          4071 => x"83",
          4072 => x"2a",
          4073 => x"56",
          4074 => x"39",
          4075 => x"83",
          4076 => x"81",
          4077 => x"7c",
          4078 => x"38",
          4079 => x"f3",
          4080 => x"06",
          4081 => x"8a",
          4082 => x"06",
          4083 => x"38",
          4084 => x"7a",
          4085 => x"77",
          4086 => x"08",
          4087 => x"82",
          4088 => x"38",
          4089 => x"98",
          4090 => x"74",
          4091 => x"08",
          4092 => x"8e",
          4093 => x"82",
          4094 => x"18",
          4095 => x"3f",
          4096 => x"d0",
          4097 => x"89",
          4098 => x"d7",
          4099 => x"58",
          4100 => x"75",
          4101 => x"7c",
          4102 => x"c2",
          4103 => x"38",
          4104 => x"56",
          4105 => x"53",
          4106 => x"7d",
          4107 => x"b8",
          4108 => x"34",
          4109 => x"8c",
          4110 => x"38",
          4111 => x"e0",
          4112 => x"b4",
          4113 => x"94",
          4114 => x"71",
          4115 => x"38",
          4116 => x"51",
          4117 => x"08",
          4118 => x"94",
          4119 => x"05",
          4120 => x"81",
          4121 => x"7e",
          4122 => x"1a",
          4123 => x"1b",
          4124 => x"27",
          4125 => x"0c",
          4126 => x"c0",
          4127 => x"56",
          4128 => x"0d",
          4129 => x"fc",
          4130 => x"3f",
          4131 => x"98",
          4132 => x"70",
          4133 => x"55",
          4134 => x"16",
          4135 => x"3f",
          4136 => x"98",
          4137 => x"8b",
          4138 => x"8b",
          4139 => x"52",
          4140 => x"16",
          4141 => x"f9",
          4142 => x"15",
          4143 => x"92",
          4144 => x"54",
          4145 => x"ff",
          4146 => x"90",
          4147 => x"73",
          4148 => x"0c",
          4149 => x"76",
          4150 => x"e0",
          4151 => x"9c",
          4152 => x"51",
          4153 => x"53",
          4154 => x"e0",
          4155 => x"98",
          4156 => x"0d",
          4157 => x"52",
          4158 => x"8b",
          4159 => x"f4",
          4160 => x"0c",
          4161 => x"80",
          4162 => x"3d",
          4163 => x"08",
          4164 => x"38",
          4165 => x"05",
          4166 => x"08",
          4167 => x"02",
          4168 => x"55",
          4169 => x"7a",
          4170 => x"a2",
          4171 => x"06",
          4172 => x"38",
          4173 => x"e1",
          4174 => x"0c",
          4175 => x"2e",
          4176 => x"74",
          4177 => x"04",
          4178 => x"08",
          4179 => x"7a",
          4180 => x"b4",
          4181 => x"d1",
          4182 => x"e0",
          4183 => x"d4",
          4184 => x"80",
          4185 => x"3d",
          4186 => x"38",
          4187 => x"55",
          4188 => x"57",
          4189 => x"80",
          4190 => x"b7",
          4191 => x"82",
          4192 => x"da",
          4193 => x"3f",
          4194 => x"0c",
          4195 => x"82",
          4196 => x"08",
          4197 => x"c9",
          4198 => x"82",
          4199 => x"3d",
          4200 => x"73",
          4201 => x"76",
          4202 => x"e0",
          4203 => x"80",
          4204 => x"81",
          4205 => x"39",
          4206 => x"fd",
          4207 => x"3f",
          4208 => x"33",
          4209 => x"92",
          4210 => x"16",
          4211 => x"73",
          4212 => x"26",
          4213 => x"38",
          4214 => x"80",
          4215 => x"18",
          4216 => x"34",
          4217 => x"3d",
          4218 => x"fd",
          4219 => x"06",
          4220 => x"08",
          4221 => x"0b",
          4222 => x"82",
          4223 => x"52",
          4224 => x"8d",
          4225 => x"51",
          4226 => x"54",
          4227 => x"74",
          4228 => x"73",
          4229 => x"81",
          4230 => x"81",
          4231 => x"81",
          4232 => x"80",
          4233 => x"54",
          4234 => x"34",
          4235 => x"34",
          4236 => x"3d",
          4237 => x"8d",
          4238 => x"55",
          4239 => x"53",
          4240 => x"91",
          4241 => x"8c",
          4242 => x"38",
          4243 => x"81",
          4244 => x"73",
          4245 => x"94",
          4246 => x"9b",
          4247 => x"2b",
          4248 => x"38",
          4249 => x"88",
          4250 => x"78",
          4251 => x"f8",
          4252 => x"96",
          4253 => x"94",
          4254 => x"08",
          4255 => x"15",
          4256 => x"74",
          4257 => x"98",
          4258 => x"2e",
          4259 => x"ff",
          4260 => x"08",
          4261 => x"73",
          4262 => x"27",
          4263 => x"16",
          4264 => x"33",
          4265 => x"55",
          4266 => x"73",
          4267 => x"82",
          4268 => x"08",
          4269 => x"a8",
          4270 => x"8b",
          4271 => x"ff",
          4272 => x"38",
          4273 => x"a7",
          4274 => x"39",
          4275 => x"75",
          4276 => x"ab",
          4277 => x"a9",
          4278 => x"82",
          4279 => x"c4",
          4280 => x"53",
          4281 => x"98",
          4282 => x"8c",
          4283 => x"8c",
          4284 => x"07",
          4285 => x"ff",
          4286 => x"77",
          4287 => x"9c",
          4288 => x"98",
          4289 => x"0d",
          4290 => x"81",
          4291 => x"05",
          4292 => x"d9",
          4293 => x"e0",
          4294 => x"0c",
          4295 => x"82",
          4296 => x"08",
          4297 => x"98",
          4298 => x"38",
          4299 => x"81",
          4300 => x"ae",
          4301 => x"c1",
          4302 => x"17",
          4303 => x"17",
          4304 => x"ea",
          4305 => x"84",
          4306 => x"55",
          4307 => x"80",
          4308 => x"98",
          4309 => x"0d",
          4310 => x"52",
          4311 => x"08",
          4312 => x"0c",
          4313 => x"77",
          4314 => x"53",
          4315 => x"98",
          4316 => x"e1",
          4317 => x"08",
          4318 => x"82",
          4319 => x"82",
          4320 => x"df",
          4321 => x"e0",
          4322 => x"85",
          4323 => x"98",
          4324 => x"ce",
          4325 => x"bd",
          4326 => x"32",
          4327 => x"70",
          4328 => x"54",
          4329 => x"3d",
          4330 => x"80",
          4331 => x"52",
          4332 => x"08",
          4333 => x"65",
          4334 => x"e0",
          4335 => x"a0",
          4336 => x"98",
          4337 => x"38",
          4338 => x"88",
          4339 => x"3f",
          4340 => x"0d",
          4341 => x"5c",
          4342 => x"93",
          4343 => x"98",
          4344 => x"82",
          4345 => x"11",
          4346 => x"56",
          4347 => x"75",
          4348 => x"81",
          4349 => x"82",
          4350 => x"73",
          4351 => x"38",
          4352 => x"3d",
          4353 => x"82",
          4354 => x"82",
          4355 => x"82",
          4356 => x"98",
          4357 => x"19",
          4358 => x"08",
          4359 => x"a8",
          4360 => x"58",
          4361 => x"7d",
          4362 => x"e0",
          4363 => x"80",
          4364 => x"ff",
          4365 => x"2e",
          4366 => x"51",
          4367 => x"08",
          4368 => x"80",
          4369 => x"54",
          4370 => x"88",
          4371 => x"06",
          4372 => x"19",
          4373 => x"06",
          4374 => x"78",
          4375 => x"84",
          4376 => x"84",
          4377 => x"92",
          4378 => x"8a",
          4379 => x"e3",
          4380 => x"82",
          4381 => x"17",
          4382 => x"17",
          4383 => x"51",
          4384 => x"81",
          4385 => x"8c",
          4386 => x"9c",
          4387 => x"17",
          4388 => x"3f",
          4389 => x"0c",
          4390 => x"52",
          4391 => x"e0",
          4392 => x"83",
          4393 => x"81",
          4394 => x"56",
          4395 => x"82",
          4396 => x"95",
          4397 => x"98",
          4398 => x"3f",
          4399 => x"08",
          4400 => x"c0",
          4401 => x"80",
          4402 => x"75",
          4403 => x"3d",
          4404 => x"a2",
          4405 => x"51",
          4406 => x"55",
          4407 => x"78",
          4408 => x"70",
          4409 => x"98",
          4410 => x"df",
          4411 => x"85",
          4412 => x"86",
          4413 => x"2b",
          4414 => x"02",
          4415 => x"58",
          4416 => x"6c",
          4417 => x"82",
          4418 => x"81",
          4419 => x"80",
          4420 => x"08",
          4421 => x"73",
          4422 => x"52",
          4423 => x"b2",
          4424 => x"e0",
          4425 => x"98",
          4426 => x"3f",
          4427 => x"98",
          4428 => x"39",
          4429 => x"38",
          4430 => x"77",
          4431 => x"08",
          4432 => x"e0",
          4433 => x"55",
          4434 => x"2e",
          4435 => x"51",
          4436 => x"08",
          4437 => x"a8",
          4438 => x"74",
          4439 => x"04",
          4440 => x"ff",
          4441 => x"b1",
          4442 => x"e0",
          4443 => x"6a",
          4444 => x"b3",
          4445 => x"e0",
          4446 => x"9b",
          4447 => x"09",
          4448 => x"df",
          4449 => x"51",
          4450 => x"78",
          4451 => x"57",
          4452 => x"08",
          4453 => x"83",
          4454 => x"81",
          4455 => x"54",
          4456 => x"81",
          4457 => x"39",
          4458 => x"08",
          4459 => x"82",
          4460 => x"08",
          4461 => x"b8",
          4462 => x"54",
          4463 => x"90",
          4464 => x"b2",
          4465 => x"a3",
          4466 => x"53",
          4467 => x"78",
          4468 => x"ff",
          4469 => x"80",
          4470 => x"d8",
          4471 => x"78",
          4472 => x"51",
          4473 => x"08",
          4474 => x"82",
          4475 => x"51",
          4476 => x"52",
          4477 => x"54",
          4478 => x"81",
          4479 => x"a6",
          4480 => x"8b",
          4481 => x"ff",
          4482 => x"0c",
          4483 => x"ab",
          4484 => x"82",
          4485 => x"ab",
          4486 => x"98",
          4487 => x"d8",
          4488 => x"9e",
          4489 => x"82",
          4490 => x"08",
          4491 => x"33",
          4492 => x"82",
          4493 => x"52",
          4494 => x"a2",
          4495 => x"3d",
          4496 => x"ac",
          4497 => x"3f",
          4498 => x"98",
          4499 => x"2e",
          4500 => x"3d",
          4501 => x"e8",
          4502 => x"09",
          4503 => x"ff",
          4504 => x"55",
          4505 => x"68",
          4506 => x"05",
          4507 => x"3f",
          4508 => x"8b",
          4509 => x"06",
          4510 => x"a0",
          4511 => x"54",
          4512 => x"33",
          4513 => x"55",
          4514 => x"6f",
          4515 => x"78",
          4516 => x"98",
          4517 => x"3f",
          4518 => x"2e",
          4519 => x"52",
          4520 => x"e0",
          4521 => x"58",
          4522 => x"38",
          4523 => x"09",
          4524 => x"52",
          4525 => x"54",
          4526 => x"82",
          4527 => x"c1",
          4528 => x"82",
          4529 => x"ff",
          4530 => x"55",
          4531 => x"0d",
          4532 => x"05",
          4533 => x"33",
          4534 => x"05",
          4535 => x"82",
          4536 => x"08",
          4537 => x"96",
          4538 => x"82",
          4539 => x"08",
          4540 => x"81",
          4541 => x"38",
          4542 => x"12",
          4543 => x"51",
          4544 => x"78",
          4545 => x"51",
          4546 => x"08",
          4547 => x"3d",
          4548 => x"82",
          4549 => x"3d",
          4550 => x"08",
          4551 => x"38",
          4552 => x"05",
          4553 => x"08",
          4554 => x"02",
          4555 => x"54",
          4556 => x"22",
          4557 => x"53",
          4558 => x"3f",
          4559 => x"76",
          4560 => x"98",
          4561 => x"94",
          4562 => x"6c",
          4563 => x"05",
          4564 => x"82",
          4565 => x"30",
          4566 => x"25",
          4567 => x"86",
          4568 => x"73",
          4569 => x"80",
          4570 => x"54",
          4571 => x"08",
          4572 => x"38",
          4573 => x"3f",
          4574 => x"98",
          4575 => x"82",
          4576 => x"78",
          4577 => x"55",
          4578 => x"8a",
          4579 => x"1a",
          4580 => x"9e",
          4581 => x"51",
          4582 => x"8e",
          4583 => x"86",
          4584 => x"30",
          4585 => x"7a",
          4586 => x"2e",
          4587 => x"51",
          4588 => x"08",
          4589 => x"7b",
          4590 => x"73",
          4591 => x"73",
          4592 => x"15",
          4593 => x"82",
          4594 => x"e0",
          4595 => x"3d",
          4596 => x"05",
          4597 => x"82",
          4598 => x"56",
          4599 => x"38",
          4600 => x"52",
          4601 => x"70",
          4602 => x"81",
          4603 => x"ff",
          4604 => x"83",
          4605 => x"e0",
          4606 => x"b5",
          4607 => x"90",
          4608 => x"ff",
          4609 => x"74",
          4610 => x"ee",
          4611 => x"81",
          4612 => x"26",
          4613 => x"86",
          4614 => x"ff",
          4615 => x"54",
          4616 => x"81",
          4617 => x"59",
          4618 => x"55",
          4619 => x"8a",
          4620 => x"e5",
          4621 => x"99",
          4622 => x"70",
          4623 => x"81",
          4624 => x"ed",
          4625 => x"90",
          4626 => x"3f",
          4627 => x"98",
          4628 => x"51",
          4629 => x"08",
          4630 => x"75",
          4631 => x"34",
          4632 => x"84",
          4633 => x"80",
          4634 => x"81",
          4635 => x"82",
          4636 => x"08",
          4637 => x"08",
          4638 => x"66",
          4639 => x"53",
          4640 => x"3f",
          4641 => x"78",
          4642 => x"98",
          4643 => x"98",
          4644 => x"0d",
          4645 => x"05",
          4646 => x"54",
          4647 => x"e0",
          4648 => x"82",
          4649 => x"82",
          4650 => x"8c",
          4651 => x"1a",
          4652 => x"51",
          4653 => x"82",
          4654 => x"81",
          4655 => x"22",
          4656 => x"56",
          4657 => x"14",
          4658 => x"9f",
          4659 => x"19",
          4660 => x"81",
          4661 => x"77",
          4662 => x"56",
          4663 => x"ff",
          4664 => x"55",
          4665 => x"82",
          4666 => x"ff",
          4667 => x"2e",
          4668 => x"8e",
          4669 => x"09",
          4670 => x"59",
          4671 => x"06",
          4672 => x"39",
          4673 => x"55",
          4674 => x"15",
          4675 => x"83",
          4676 => x"7e",
          4677 => x"98",
          4678 => x"ce",
          4679 => x"56",
          4680 => x"19",
          4681 => x"7d",
          4682 => x"0c",
          4683 => x"80",
          4684 => x"9c",
          4685 => x"57",
          4686 => x"7b",
          4687 => x"81",
          4688 => x"54",
          4689 => x"0d",
          4690 => x"88",
          4691 => x"54",
          4692 => x"56",
          4693 => x"8d",
          4694 => x"29",
          4695 => x"55",
          4696 => x"34",
          4697 => x"08",
          4698 => x"e0",
          4699 => x"52",
          4700 => x"e0",
          4701 => x"06",
          4702 => x"38",
          4703 => x"55",
          4704 => x"3d",
          4705 => x"ff",
          4706 => x"99",
          4707 => x"38",
          4708 => x"ff",
          4709 => x"83",
          4710 => x"38",
          4711 => x"81",
          4712 => x"79",
          4713 => x"93",
          4714 => x"6f",
          4715 => x"49",
          4716 => x"61",
          4717 => x"55",
          4718 => x"80",
          4719 => x"53",
          4720 => x"3f",
          4721 => x"c1",
          4722 => x"f1",
          4723 => x"ff",
          4724 => x"d5",
          4725 => x"64",
          4726 => x"56",
          4727 => x"83",
          4728 => x"82",
          4729 => x"5f",
          4730 => x"08",
          4731 => x"53",
          4732 => x"3f",
          4733 => x"e1",
          4734 => x"82",
          4735 => x"83",
          4736 => x"7e",
          4737 => x"31",
          4738 => x"8a",
          4739 => x"26",
          4740 => x"81",
          4741 => x"38",
          4742 => x"83",
          4743 => x"80",
          4744 => x"55",
          4745 => x"8a",
          4746 => x"09",
          4747 => x"38",
          4748 => x"d3",
          4749 => x"9d",
          4750 => x"d3",
          4751 => x"22",
          4752 => x"38",
          4753 => x"67",
          4754 => x"98",
          4755 => x"89",
          4756 => x"82",
          4757 => x"56",
          4758 => x"80",
          4759 => x"38",
          4760 => x"d3",
          4761 => x"9d",
          4762 => x"d3",
          4763 => x"22",
          4764 => x"38",
          4765 => x"67",
          4766 => x"98",
          4767 => x"98",
          4768 => x"0b",
          4769 => x"98",
          4770 => x"05",
          4771 => x"2a",
          4772 => x"7d",
          4773 => x"05",
          4774 => x"5c",
          4775 => x"2e",
          4776 => x"61",
          4777 => x"5d",
          4778 => x"69",
          4779 => x"e4",
          4780 => x"53",
          4781 => x"e8",
          4782 => x"83",
          4783 => x"e0",
          4784 => x"dd",
          4785 => x"2a",
          4786 => x"39",
          4787 => x"c5",
          4788 => x"98",
          4789 => x"79",
          4790 => x"38",
          4791 => x"06",
          4792 => x"5e",
          4793 => x"9f",
          4794 => x"38",
          4795 => x"fc",
          4796 => x"7d",
          4797 => x"7d",
          4798 => x"74",
          4799 => x"d1",
          4800 => x"51",
          4801 => x"d1",
          4802 => x"3f",
          4803 => x"8e",
          4804 => x"83",
          4805 => x"ff",
          4806 => x"34",
          4807 => x"2a",
          4808 => x"1b",
          4809 => x"74",
          4810 => x"83",
          4811 => x"ff",
          4812 => x"a0",
          4813 => x"0b",
          4814 => x"51",
          4815 => x"9a",
          4816 => x"52",
          4817 => x"7d",
          4818 => x"38",
          4819 => x"1b",
          4820 => x"a4",
          4821 => x"52",
          4822 => x"81",
          4823 => x"3f",
          4824 => x"83",
          4825 => x"34",
          4826 => x"53",
          4827 => x"51",
          4828 => x"a7",
          4829 => x"83",
          4830 => x"ff",
          4831 => x"1c",
          4832 => x"53",
          4833 => x"ff",
          4834 => x"83",
          4835 => x"ab",
          4836 => x"7f",
          4837 => x"82",
          4838 => x"83",
          4839 => x"75",
          4840 => x"51",
          4841 => x"80",
          4842 => x"84",
          4843 => x"ff",
          4844 => x"f2",
          4845 => x"f9",
          4846 => x"51",
          4847 => x"ec",
          4848 => x"d4",
          4849 => x"3f",
          4850 => x"7f",
          4851 => x"75",
          4852 => x"87",
          4853 => x"51",
          4854 => x"58",
          4855 => x"38",
          4856 => x"3f",
          4857 => x"99",
          4858 => x"91",
          4859 => x"81",
          4860 => x"7a",
          4861 => x"61",
          4862 => x"57",
          4863 => x"51",
          4864 => x"08",
          4865 => x"e0",
          4866 => x"a3",
          4867 => x"56",
          4868 => x"80",
          4869 => x"83",
          4870 => x"74",
          4871 => x"54",
          4872 => x"86",
          4873 => x"f8",
          4874 => x"56",
          4875 => x"2e",
          4876 => x"ff",
          4877 => x"2e",
          4878 => x"b2",
          4879 => x"7f",
          4880 => x"82",
          4881 => x"90",
          4882 => x"34",
          4883 => x"7a",
          4884 => x"81",
          4885 => x"58",
          4886 => x"77",
          4887 => x"82",
          4888 => x"83",
          4889 => x"34",
          4890 => x"82",
          4891 => x"84",
          4892 => x"c1",
          4893 => x"fe",
          4894 => x"08",
          4895 => x"16",
          4896 => x"34",
          4897 => x"88",
          4898 => x"51",
          4899 => x"53",
          4900 => x"3f",
          4901 => x"38",
          4902 => x"86",
          4903 => x"08",
          4904 => x"39",
          4905 => x"08",
          4906 => x"3d",
          4907 => x"5b",
          4908 => x"57",
          4909 => x"3d",
          4910 => x"15",
          4911 => x"81",
          4912 => x"3d",
          4913 => x"74",
          4914 => x"17",
          4915 => x"c9",
          4916 => x"83",
          4917 => x"0c",
          4918 => x"7b",
          4919 => x"57",
          4920 => x"38",
          4921 => x"17",
          4922 => x"88",
          4923 => x"59",
          4924 => x"76",
          4925 => x"54",
          4926 => x"51",
          4927 => x"30",
          4928 => x"53",
          4929 => x"81",
          4930 => x"04",
          4931 => x"56",
          4932 => x"3d",
          4933 => x"52",
          4934 => x"e0",
          4935 => x"78",
          4936 => x"16",
          4937 => x"82",
          4938 => x"fd",
          4939 => x"80",
          4940 => x"76",
          4941 => x"3d",
          4942 => x"53",
          4943 => x"3f",
          4944 => x"72",
          4945 => x"04",
          4946 => x"9a",
          4947 => x"80",
          4948 => x"ff",
          4949 => x"ff",
          4950 => x"09",
          4951 => x"af",
          4952 => x"71",
          4953 => x"ff",
          4954 => x"26",
          4955 => x"05",
          4956 => x"80",
          4957 => x"71",
          4958 => x"04",
          4959 => x"02",
          4960 => x"80",
          4961 => x"70",
          4962 => x"09",
          4963 => x"26",
          4964 => x"05",
          4965 => x"98",
          4966 => x"0d",
          4967 => x"81",
          4968 => x"82",
          4969 => x"27",
          4970 => x"70",
          4971 => x"80",
          4972 => x"55",
          4973 => x"05",
          4974 => x"ff",
          4975 => x"71",
          4976 => x"26",
          4977 => x"b9",
          4978 => x"75",
          4979 => x"51",
          4980 => x"81",
          4981 => x"39",
          4982 => x"51",
          4983 => x"e6",
          4984 => x"8b",
          4985 => x"c7",
          4986 => x"06",
          4987 => x"72",
          4988 => x"51",
          4989 => x"0d",
          4990 => x"ff",
          4991 => x"ff",
          4992 => x"30",
          4993 => x"30",
          4994 => x"30",
          4995 => x"30",
          4996 => x"30",
          4997 => x"30",
          4998 => x"30",
          4999 => x"30",
          5000 => x"30",
          5001 => x"30",
          5002 => x"47",
          5003 => x"47",
          5004 => x"4d",
          5005 => x"4f",
          5006 => x"4e",
          5007 => x"50",
          5008 => x"50",
          5009 => x"50",
          5010 => x"4c",
          5011 => x"4f",
          5012 => x"4c",
          5013 => x"50",
          5014 => x"51",
          5015 => x"9b",
          5016 => x"9b",
          5017 => x"9b",
          5018 => x"9b",
          5019 => x"9b",
          5020 => x"17",
          5021 => x"0e",
          5022 => x"17",
          5023 => x"17",
          5024 => x"17",
          5025 => x"0e",
          5026 => x"0e",
          5027 => x"17",
          5028 => x"17",
          5029 => x"17",
          5030 => x"17",
          5031 => x"17",
          5032 => x"17",
          5033 => x"17",
          5034 => x"17",
          5035 => x"17",
          5036 => x"17",
          5037 => x"17",
          5038 => x"17",
          5039 => x"17",
          5040 => x"17",
          5041 => x"17",
          5042 => x"17",
          5043 => x"17",
          5044 => x"17",
          5045 => x"0f",
          5046 => x"17",
          5047 => x"17",
          5048 => x"17",
          5049 => x"17",
          5050 => x"17",
          5051 => x"17",
          5052 => x"17",
          5053 => x"0f",
          5054 => x"0e",
          5055 => x"0e",
          5056 => x"10",
          5057 => x"17",
          5058 => x"17",
          5059 => x"11",
          5060 => x"17",
          5061 => x"0f",
          5062 => x"11",
          5063 => x"17",
          5064 => x"6e",
          5065 => x"6f",
          5066 => x"6e",
          5067 => x"6f",
          5068 => x"78",
          5069 => x"6c",
          5070 => x"6f",
          5071 => x"69",
          5072 => x"75",
          5073 => x"62",
          5074 => x"77",
          5075 => x"65",
          5076 => x"65",
          5077 => x"00",
          5078 => x"73",
          5079 => x"73",
          5080 => x"66",
          5081 => x"61",
          5082 => x"61",
          5083 => x"6c",
          5084 => x"00",
          5085 => x"72",
          5086 => x"74",
          5087 => x"72",
          5088 => x"73",
          5089 => x"65",
          5090 => x"20",
          5091 => x"75",
          5092 => x"20",
          5093 => x"75",
          5094 => x"76",
          5095 => x"6c",
          5096 => x"00",
          5097 => x"20",
          5098 => x"00",
          5099 => x"6c",
          5100 => x"78",
          5101 => x"00",
          5102 => x"61",
          5103 => x"76",
          5104 => x"00",
          5105 => x"77",
          5106 => x"6f",
          5107 => x"00",
          5108 => x"6e",
          5109 => x"73",
          5110 => x"64",
          5111 => x"73",
          5112 => x"6e",
          5113 => x"00",
          5114 => x"70",
          5115 => x"66",
          5116 => x"65",
          5117 => x"20",
          5118 => x"2e",
          5119 => x"20",
          5120 => x"2e",
          5121 => x"74",
          5122 => x"74",
          5123 => x"63",
          5124 => x"00",
          5125 => x"73",
          5126 => x"2e",
          5127 => x"69",
          5128 => x"65",
          5129 => x"00",
          5130 => x"6e",
          5131 => x"66",
          5132 => x"00",
          5133 => x"74",
          5134 => x"6f",
          5135 => x"00",
          5136 => x"73",
          5137 => x"6b",
          5138 => x"72",
          5139 => x"6c",
          5140 => x"20",
          5141 => x"6c",
          5142 => x"2f",
          5143 => x"00",
          5144 => x"00",
          5145 => x"00",
          5146 => x"34",
          5147 => x"20",
          5148 => x"00",
          5149 => x"00",
          5150 => x"00",
          5151 => x"53",
          5152 => x"28",
          5153 => x"32",
          5154 => x"2e",
          5155 => x"50",
          5156 => x"25",
          5157 => x"20",
          5158 => x"00",
          5159 => x"74",
          5160 => x"48",
          5161 => x"00",
          5162 => x"69",
          5163 => x"74",
          5164 => x"74",
          5165 => x"00",
          5166 => x"52",
          5167 => x"72",
          5168 => x"43",
          5169 => x"6e",
          5170 => x"00",
          5171 => x"52",
          5172 => x"72",
          5173 => x"52",
          5174 => x"6e",
          5175 => x"00",
          5176 => x"52",
          5177 => x"72",
          5178 => x"52",
          5179 => x"6e",
          5180 => x"00",
          5181 => x"67",
          5182 => x"65",
          5183 => x"61",
          5184 => x"69",
          5185 => x"00",
          5186 => x"65",
          5187 => x"00",
          5188 => x"75",
          5189 => x"00",
          5190 => x"20",
          5191 => x"69",
          5192 => x"64",
          5193 => x"2c",
          5194 => x"20",
          5195 => x"6e",
          5196 => x"00",
          5197 => x"65",
          5198 => x"2e",
          5199 => x"70",
          5200 => x"00",
          5201 => x"69",
          5202 => x"00",
          5203 => x"25",
          5204 => x"30",
          5205 => x"78",
          5206 => x"6d",
          5207 => x"79",
          5208 => x"65",
          5209 => x"38",
          5210 => x"2d",
          5211 => x"38",
          5212 => x"2d",
          5213 => x"25",
          5214 => x"00",
          5215 => x"69",
          5216 => x"20",
          5217 => x"20",
          5218 => x"6c",
          5219 => x"64",
          5220 => x"6c",
          5221 => x"00",
          5222 => x"65",
          5223 => x"63",
          5224 => x"29",
          5225 => x"73",
          5226 => x"20",
          5227 => x"74",
          5228 => x"00",
          5229 => x"65",
          5230 => x"2e",
          5231 => x"55",
          5232 => x"3a",
          5233 => x"25",
          5234 => x"3a",
          5235 => x"00",
          5236 => x"00",
          5237 => x"6d",
          5238 => x"00",
          5239 => x"20",
          5240 => x"65",
          5241 => x"6f",
          5242 => x"73",
          5243 => x"6e",
          5244 => x"6e",
          5245 => x"00",
          5246 => x"6e",
          5247 => x"72",
          5248 => x"00",
          5249 => x"25",
          5250 => x"3a",
          5251 => x"0a",
          5252 => x"6e",
          5253 => x"69",
          5254 => x"66",
          5255 => x"20",
          5256 => x"00",
          5257 => x"63",
          5258 => x"65",
          5259 => x"00",
          5260 => x"20",
          5261 => x"28",
          5262 => x"38",
          5263 => x"20",
          5264 => x"20",
          5265 => x"58",
          5266 => x"0a",
          5267 => x"53",
          5268 => x"28",
          5269 => x"38",
          5270 => x"20",
          5271 => x"20",
          5272 => x"58",
          5273 => x"0a",
          5274 => x"4d",
          5275 => x"28",
          5276 => x"38",
          5277 => x"20",
          5278 => x"44",
          5279 => x"69",
          5280 => x"32",
          5281 => x"20",
          5282 => x"20",
          5283 => x"65",
          5284 => x"32",
          5285 => x"20",
          5286 => x"54",
          5287 => x"6e",
          5288 => x"32",
          5289 => x"20",
          5290 => x"4e",
          5291 => x"00",
          5292 => x"20",
          5293 => x"20",
          5294 => x"00",
          5295 => x"32",
          5296 => x"49",
          5297 => x"73",
          5298 => x"20",
          5299 => x"73",
          5300 => x"6f",
          5301 => x"73",
          5302 => x"58",
          5303 => x"20",
          5304 => x"6d",
          5305 => x"72",
          5306 => x"73",
          5307 => x"58",
          5308 => x"20",
          5309 => x"53",
          5310 => x"64",
          5311 => x"20",
          5312 => x"58",
          5313 => x"73",
          5314 => x"20",
          5315 => x"20",
          5316 => x"20",
          5317 => x"20",
          5318 => x"58",
          5319 => x"20",
          5320 => x"20",
          5321 => x"72",
          5322 => x"20",
          5323 => x"25",
          5324 => x"00",
          5325 => x"52",
          5326 => x"6b",
          5327 => x"20",
          5328 => x"20",
          5329 => x"4d",
          5330 => x"20",
          5331 => x"6e",
          5332 => x"20",
          5333 => x"72",
          5334 => x"25",
          5335 => x"00",
          5336 => x"00",
          5337 => x"00",
          5338 => x"00",
          5339 => x"4f",
          5340 => x"6b",
          5341 => x"a8",
          5342 => x"00",
          5343 => x"00",
          5344 => x"a8",
          5345 => x"00",
          5346 => x"00",
          5347 => x"a8",
          5348 => x"00",
          5349 => x"00",
          5350 => x"a8",
          5351 => x"00",
          5352 => x"00",
          5353 => x"a8",
          5354 => x"00",
          5355 => x"00",
          5356 => x"a8",
          5357 => x"00",
          5358 => x"00",
          5359 => x"a8",
          5360 => x"00",
          5361 => x"00",
          5362 => x"a8",
          5363 => x"00",
          5364 => x"00",
          5365 => x"a8",
          5366 => x"00",
          5367 => x"00",
          5368 => x"a7",
          5369 => x"00",
          5370 => x"00",
          5371 => x"a7",
          5372 => x"00",
          5373 => x"00",
          5374 => x"44",
          5375 => x"42",
          5376 => x"36",
          5377 => x"34",
          5378 => x"33",
          5379 => x"31",
          5380 => x"00",
          5381 => x"00",
          5382 => x"00",
          5383 => x"00",
          5384 => x"00",
          5385 => x"73",
          5386 => x"73",
          5387 => x"00",
          5388 => x"20",
          5389 => x"69",
          5390 => x"72",
          5391 => x"65",
          5392 => x"79",
          5393 => x"6f",
          5394 => x"00",
          5395 => x"20",
          5396 => x"65",
          5397 => x"74",
          5398 => x"65",
          5399 => x"6c",
          5400 => x"00",
          5401 => x"7c",
          5402 => x"3b",
          5403 => x"54",
          5404 => x"00",
          5405 => x"4f",
          5406 => x"20",
          5407 => x"20",
          5408 => x"20",
          5409 => x"45",
          5410 => x"20",
          5411 => x"a8",
          5412 => x"00",
          5413 => x"05",
          5414 => x"18",
          5415 => x"45",
          5416 => x"45",
          5417 => x"92",
          5418 => x"9a",
          5419 => x"4f",
          5420 => x"aa",
          5421 => x"b2",
          5422 => x"ba",
          5423 => x"c2",
          5424 => x"ca",
          5425 => x"d2",
          5426 => x"da",
          5427 => x"e2",
          5428 => x"ea",
          5429 => x"f2",
          5430 => x"fa",
          5431 => x"2c",
          5432 => x"2a",
          5433 => x"00",
          5434 => x"00",
          5435 => x"00",
          5436 => x"00",
          5437 => x"00",
          5438 => x"00",
          5439 => x"00",
          5440 => x"00",
          5441 => x"00",
          5442 => x"00",
          5443 => x"00",
          5444 => x"00",
          5445 => x"01",
          5446 => x"00",
          5447 => x"00",
          5448 => x"00",
          5449 => x"00",
          5450 => x"25",
          5451 => x"25",
          5452 => x"25",
          5453 => x"25",
          5454 => x"25",
          5455 => x"25",
          5456 => x"25",
          5457 => x"25",
          5458 => x"25",
          5459 => x"25",
          5460 => x"25",
          5461 => x"25",
          5462 => x"03",
          5463 => x"03",
          5464 => x"03",
          5465 => x"22",
          5466 => x"22",
          5467 => x"22",
          5468 => x"22",
          5469 => x"00",
          5470 => x"03",
          5471 => x"00",
          5472 => x"01",
          5473 => x"01",
          5474 => x"01",
          5475 => x"01",
          5476 => x"01",
          5477 => x"01",
          5478 => x"01",
          5479 => x"01",
          5480 => x"01",
          5481 => x"02",
          5482 => x"02",
          5483 => x"01",
          5484 => x"01",
          5485 => x"01",
          5486 => x"01",
          5487 => x"01",
          5488 => x"01",
          5489 => x"01",
          5490 => x"01",
          5491 => x"01",
          5492 => x"01",
          5493 => x"01",
          5494 => x"01",
          5495 => x"01",
          5496 => x"01",
          5497 => x"01",
          5498 => x"00",
          5499 => x"02",
          5500 => x"02",
          5501 => x"02",
          5502 => x"02",
          5503 => x"01",
          5504 => x"02",
          5505 => x"02",
          5506 => x"02",
          5507 => x"01",
          5508 => x"02",
          5509 => x"02",
          5510 => x"01",
          5511 => x"02",
          5512 => x"2c",
          5513 => x"02",
          5514 => x"02",
          5515 => x"02",
          5516 => x"02",
          5517 => x"02",
          5518 => x"03",
          5519 => x"00",
          5520 => x"03",
          5521 => x"00",
          5522 => x"03",
          5523 => x"03",
          5524 => x"03",
          5525 => x"03",
          5526 => x"03",
          5527 => x"04",
          5528 => x"04",
          5529 => x"04",
          5530 => x"04",
          5531 => x"04",
          5532 => x"00",
          5533 => x"1e",
          5534 => x"1f",
          5535 => x"1f",
          5536 => x"1f",
          5537 => x"1f",
          5538 => x"1f",
          5539 => x"00",
          5540 => x"1f",
          5541 => x"1f",
          5542 => x"1f",
          5543 => x"06",
          5544 => x"06",
          5545 => x"1f",
          5546 => x"00",
          5547 => x"1f",
          5548 => x"1f",
          5549 => x"21",
          5550 => x"02",
          5551 => x"24",
          5552 => x"2c",
          5553 => x"2c",
          5554 => x"2d",
          5555 => x"00",
          5556 => x"9e",
          5557 => x"00",
          5558 => x"9e",
          5559 => x"00",
          5560 => x"9e",
          5561 => x"00",
          5562 => x"9e",
          5563 => x"00",
          5564 => x"9e",
          5565 => x"00",
          5566 => x"9e",
          5567 => x"00",
          5568 => x"9e",
          5569 => x"00",
          5570 => x"9e",
          5571 => x"00",
          5572 => x"9e",
          5573 => x"00",
          5574 => x"9e",
          5575 => x"00",
          5576 => x"9e",
          5577 => x"00",
          5578 => x"9e",
          5579 => x"00",
          5580 => x"9e",
          5581 => x"00",
          5582 => x"9e",
          5583 => x"00",
          5584 => x"9e",
          5585 => x"00",
          5586 => x"9e",
          5587 => x"00",
          5588 => x"9e",
          5589 => x"00",
          5590 => x"9e",
          5591 => x"00",
          5592 => x"9e",
          5593 => x"00",
          5594 => x"9e",
          5595 => x"00",
          5596 => x"9e",
          5597 => x"00",
          5598 => x"9e",
          5599 => x"00",
          5600 => x"9e",
          5601 => x"00",
          5602 => x"9e",
          5603 => x"00",
          5604 => x"9e",
          5605 => x"00",
          5606 => x"00",
          5607 => x"7f",
          5608 => x"7f",
          5609 => x"7f",
          5610 => x"00",
          5611 => x"ff",
          5612 => x"00",
          5613 => x"00",
          5614 => x"e1",
          5615 => x"00",
          5616 => x"01",
          5617 => x"00",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"00",
          5630 => x"00",
          5631 => x"00",
          5632 => x"00",
          5633 => x"00",
          5634 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"93",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"2d",
             6 => x"00",
             7 => x"00",
             8 => x"fd",
             9 => x"05",
            10 => x"ff",
            11 => x"00",
            12 => x"fd",
            13 => x"06",
            14 => x"2b",
            15 => x"0b",
            16 => x"09",
            17 => x"06",
            18 => x"0a",
            19 => x"00",
            20 => x"72",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"73",
            25 => x"81",
            26 => x"10",
            27 => x"51",
            28 => x"72",
            29 => x"04",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"74",
            50 => x"07",
            51 => x"00",
            52 => x"71",
            53 => x"09",
            54 => x"2b",
            55 => x"04",
            56 => x"09",
            57 => x"05",
            58 => x"04",
            59 => x"00",
            60 => x"09",
            61 => x"05",
            62 => x"51",
            63 => x"00",
            64 => x"09",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"53",
            74 => x"00",
            75 => x"00",
            76 => x"fc",
            77 => x"05",
            78 => x"ff",
            79 => x"00",
            80 => x"fc",
            81 => x"73",
            82 => x"0b",
            83 => x"00",
            84 => x"08",
            85 => x"0b",
            86 => x"08",
            87 => x"51",
            88 => x"08",
            89 => x"0b",
            90 => x"08",
            91 => x"51",
            92 => x"09",
            93 => x"06",
            94 => x"09",
            95 => x"51",
            96 => x"09",
            97 => x"81",
            98 => x"73",
            99 => x"07",
           100 => x"ff",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"81",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"84",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"0d",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"92",
           173 => x"04",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"00",
           193 => x"81",
           194 => x"80",
           195 => x"0c",
           196 => x"80",
           197 => x"0c",
           198 => x"80",
           199 => x"0c",
           200 => x"80",
           201 => x"0c",
           202 => x"80",
           203 => x"0c",
           204 => x"80",
           205 => x"0c",
           206 => x"08",
           207 => x"a4",
           208 => x"a4",
           209 => x"e0",
           210 => x"a4",
           211 => x"e0",
           212 => x"a4",
           213 => x"e0",
           214 => x"a4",
           215 => x"e0",
           216 => x"e0",
           217 => x"82",
           218 => x"82",
           219 => x"04",
           220 => x"2d",
           221 => x"90",
           222 => x"b2",
           223 => x"80",
           224 => x"fe",
           225 => x"c0",
           226 => x"81",
           227 => x"80",
           228 => x"0c",
           229 => x"08",
           230 => x"a4",
           231 => x"a4",
           232 => x"e0",
           233 => x"e0",
           234 => x"82",
           235 => x"82",
           236 => x"04",
           237 => x"2d",
           238 => x"90",
           239 => x"84",
           240 => x"80",
           241 => x"8c",
           242 => x"c0",
           243 => x"82",
           244 => x"80",
           245 => x"0c",
           246 => x"08",
           247 => x"a4",
           248 => x"a4",
           249 => x"e0",
           250 => x"e0",
           251 => x"82",
           252 => x"82",
           253 => x"04",
           254 => x"2d",
           255 => x"90",
           256 => x"9c",
           257 => x"80",
           258 => x"9c",
           259 => x"c0",
           260 => x"82",
           261 => x"80",
           262 => x"0c",
           263 => x"08",
           264 => x"a4",
           265 => x"a4",
           266 => x"e0",
           267 => x"e0",
           268 => x"82",
           269 => x"82",
           270 => x"04",
           271 => x"2d",
           272 => x"90",
           273 => x"a0",
           274 => x"80",
           275 => x"f5",
           276 => x"c0",
           277 => x"82",
           278 => x"80",
           279 => x"0c",
           280 => x"08",
           281 => x"a4",
           282 => x"a4",
           283 => x"e0",
           284 => x"e0",
           285 => x"82",
           286 => x"82",
           287 => x"04",
           288 => x"2d",
           289 => x"90",
           290 => x"e4",
           291 => x"80",
           292 => x"fd",
           293 => x"c0",
           294 => x"81",
           295 => x"80",
           296 => x"0c",
           297 => x"08",
           298 => x"a4",
           299 => x"a4",
           300 => x"e0",
           301 => x"e0",
           302 => x"82",
           303 => x"82",
           304 => x"04",
           305 => x"2d",
           306 => x"90",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"10",
           311 => x"73",
           312 => x"81",
           313 => x"07",
           314 => x"72",
           315 => x"09",
           316 => x"0a",
           317 => x"51",
           318 => x"82",
           319 => x"70",
           320 => x"93",
           321 => x"a7",
           322 => x"82",
           323 => x"e0",
           324 => x"a4",
           325 => x"08",
           326 => x"08",
           327 => x"08",
           328 => x"98",
           329 => x"05",
           330 => x"08",
           331 => x"87",
           332 => x"82",
           333 => x"0c",
           334 => x"90",
           335 => x"32",
           336 => x"71",
           337 => x"08",
           338 => x"39",
           339 => x"05",
           340 => x"08",
           341 => x"a4",
           342 => x"e0",
           343 => x"a4",
           344 => x"08",
           345 => x"f8",
           346 => x"80",
           347 => x"08",
           348 => x"08",
           349 => x"82",
           350 => x"08",
           351 => x"08",
           352 => x"06",
           353 => x"08",
           354 => x"e0",
           355 => x"a4",
           356 => x"73",
           357 => x"08",
           358 => x"05",
           359 => x"08",
           360 => x"05",
           361 => x"08",
           362 => x"82",
           363 => x"82",
           364 => x"82",
           365 => x"e0",
           366 => x"a4",
           367 => x"82",
           368 => x"0b",
           369 => x"82",
           370 => x"e0",
           371 => x"0b",
           372 => x"82",
           373 => x"e0",
           374 => x"a4",
           375 => x"a4",
           376 => x"a4",
           377 => x"81",
           378 => x"82",
           379 => x"e0",
           380 => x"a4",
           381 => x"80",
           382 => x"05",
           383 => x"8e",
           384 => x"82",
           385 => x"0c",
           386 => x"90",
           387 => x"05",
           388 => x"08",
           389 => x"08",
           390 => x"08",
           391 => x"08",
           392 => x"0c",
           393 => x"70",
           394 => x"3d",
           395 => x"e0",
           396 => x"ed",
           397 => x"08",
           398 => x"88",
           399 => x"0c",
           400 => x"85",
           401 => x"32",
           402 => x"53",
           403 => x"82",
           404 => x"ac",
           405 => x"08",
           406 => x"a4",
           407 => x"06",
           408 => x"82",
           409 => x"05",
           410 => x"82",
           411 => x"81",
           412 => x"8b",
           413 => x"33",
           414 => x"82",
           415 => x"72",
           416 => x"a4",
           417 => x"2e",
           418 => x"e0",
           419 => x"2b",
           420 => x"b2",
           421 => x"22",
           422 => x"81",
           423 => x"2e",
           424 => x"05",
           425 => x"72",
           426 => x"fe",
           427 => x"05",
           428 => x"70",
           429 => x"51",
           430 => x"82",
           431 => x"e0",
           432 => x"e0",
           433 => x"d0",
           434 => x"a4",
           435 => x"08",
           436 => x"98",
           437 => x"8b",
           438 => x"08",
           439 => x"e4",
           440 => x"06",
           441 => x"82",
           442 => x"88",
           443 => x"70",
           444 => x"72",
           445 => x"fd",
           446 => x"05",
           447 => x"51",
           448 => x"82",
           449 => x"98",
           450 => x"72",
           451 => x"08",
           452 => x"f8",
           453 => x"08",
           454 => x"08",
           455 => x"94",
           456 => x"08",
           457 => x"70",
           458 => x"82",
           459 => x"90",
           460 => x"08",
           461 => x"e4",
           462 => x"72",
           463 => x"fc",
           464 => x"05",
           465 => x"72",
           466 => x"fc",
           467 => x"05",
           468 => x"72",
           469 => x"fb",
           470 => x"05",
           471 => x"82",
           472 => x"0b",
           473 => x"fb",
           474 => x"05",
           475 => x"82",
           476 => x"c1",
           477 => x"fc",
           478 => x"05",
           479 => x"e0",
           480 => x"0b",
           481 => x"8d",
           482 => x"05",
           483 => x"08",
           484 => x"05",
           485 => x"e0",
           486 => x"a4",
           487 => x"53",
           488 => x"23",
           489 => x"90",
           490 => x"05",
           491 => x"90",
           492 => x"08",
           493 => x"e4",
           494 => x"06",
           495 => x"ab",
           496 => x"33",
           497 => x"53",
           498 => x"52",
           499 => x"08",
           500 => x"05",
           501 => x"fc",
           502 => x"e0",
           503 => x"08",
           504 => x"ec",
           505 => x"f4",
           506 => x"72",
           507 => x"8b",
           508 => x"05",
           509 => x"08",
           510 => x"05",
           511 => x"fc",
           512 => x"05",
           513 => x"51",
           514 => x"38",
           515 => x"70",
           516 => x"82",
           517 => x"53",
           518 => x"53",
           519 => x"23",
           520 => x"05",
           521 => x"98",
           522 => x"f4",
           523 => x"05",
           524 => x"05",
           525 => x"82",
           526 => x"c1",
           527 => x"22",
           528 => x"51",
           529 => x"e0",
           530 => x"a4",
           531 => x"e0",
           532 => x"82",
           533 => x"a2",
           534 => x"08",
           535 => x"84",
           536 => x"0c",
           537 => x"05",
           538 => x"05",
           539 => x"0c",
           540 => x"80",
           541 => x"e4",
           542 => x"72",
           543 => x"82",
           544 => x"82",
           545 => x"e0",
           546 => x"bf",
           547 => x"08",
           548 => x"0b",
           549 => x"a9",
           550 => x"22",
           551 => x"82",
           552 => x"f8",
           553 => x"34",
           554 => x"05",
           555 => x"22",
           556 => x"51",
           557 => x"e0",
           558 => x"a4",
           559 => x"e0",
           560 => x"82",
           561 => x"a2",
           562 => x"08",
           563 => x"84",
           564 => x"0c",
           565 => x"05",
           566 => x"05",
           567 => x"0c",
           568 => x"70",
           569 => x"a4",
           570 => x"0b",
           571 => x"82",
           572 => x"e0",
           573 => x"a4",
           574 => x"54",
           575 => x"e0",
           576 => x"e0",
           577 => x"a4",
           578 => x"08",
           579 => x"89",
           580 => x"08",
           581 => x"82",
           582 => x"15",
           583 => x"e0",
           584 => x"82",
           585 => x"72",
           586 => x"e0",
           587 => x"a4",
           588 => x"a4",
           589 => x"e0",
           590 => x"82",
           591 => x"e0",
           592 => x"82",
           593 => x"53",
           594 => x"70",
           595 => x"53",
           596 => x"80",
           597 => x"e0",
           598 => x"a8",
           599 => x"31",
           600 => x"fc",
           601 => x"05",
           602 => x"80",
           603 => x"ec",
           604 => x"82",
           605 => x"e0",
           606 => x"2a",
           607 => x"80",
           608 => x"08",
           609 => x"e0",
           610 => x"a4",
           611 => x"e0",
           612 => x"a4",
           613 => x"90",
           614 => x"e0",
           615 => x"53",
           616 => x"23",
           617 => x"05",
           618 => x"a4",
           619 => x"08",
           620 => x"ec",
           621 => x"05",
           622 => x"51",
           623 => x"38",
           624 => x"70",
           625 => x"a4",
           626 => x"53",
           627 => x"a4",
           628 => x"51",
           629 => x"05",
           630 => x"e8",
           631 => x"fc",
           632 => x"72",
           633 => x"82",
           634 => x"83",
           635 => x"72",
           636 => x"08",
           637 => x"90",
           638 => x"51",
           639 => x"e0",
           640 => x"31",
           641 => x"ec",
           642 => x"08",
           643 => x"90",
           644 => x"51",
           645 => x"e0",
           646 => x"31",
           647 => x"ec",
           648 => x"05",
           649 => x"72",
           650 => x"05",
           651 => x"e0",
           652 => x"2b",
           653 => x"25",
           654 => x"05",
           655 => x"d2",
           656 => x"22",
           657 => x"51",
           658 => x"e0",
           659 => x"51",
           660 => x"e0",
           661 => x"2a",
           662 => x"80",
           663 => x"88",
           664 => x"3f",
           665 => x"05",
           666 => x"51",
           667 => x"82",
           668 => x"a0",
           669 => x"08",
           670 => x"81",
           671 => x"b1",
           672 => x"08",
           673 => x"e0",
           674 => x"90",
           675 => x"e0",
           676 => x"e0",
           677 => x"bc",
           678 => x"22",
           679 => x"51",
           680 => x"e0",
           681 => x"54",
           682 => x"05",
           683 => x"51",
           684 => x"e0",
           685 => x"51",
           686 => x"a4",
           687 => x"70",
           688 => x"2e",
           689 => x"05",
           690 => x"e0",
           691 => x"2b",
           692 => x"25",
           693 => x"05",
           694 => x"d2",
           695 => x"22",
           696 => x"51",
           697 => x"08",
           698 => x"72",
           699 => x"73",
           700 => x"80",
           701 => x"08",
           702 => x"f4",
           703 => x"f8",
           704 => x"09",
           705 => x"08",
           706 => x"08",
           707 => x"81",
           708 => x"05",
           709 => x"81",
           710 => x"08",
           711 => x"72",
           712 => x"72",
           713 => x"ff",
           714 => x"a4",
           715 => x"a4",
           716 => x"82",
           717 => x"05",
           718 => x"53",
           719 => x"e0",
           720 => x"80",
           721 => x"38",
           722 => x"ff",
           723 => x"08",
           724 => x"06",
           725 => x"df",
           726 => x"08",
           727 => x"08",
           728 => x"82",
           729 => x"05",
           730 => x"ff",
           731 => x"05",
           732 => x"82",
           733 => x"82",
           734 => x"05",
           735 => x"82",
           736 => x"33",
           737 => x"82",
           738 => x"87",
           739 => x"72",
           740 => x"a4",
           741 => x"54",
           742 => x"23",
           743 => x"53",
           744 => x"a4",
           745 => x"85",
           746 => x"08",
           747 => x"08",
           748 => x"80",
           749 => x"23",
           750 => x"f8",
           751 => x"81",
           752 => x"a4",
           753 => x"e0",
           754 => x"82",
           755 => x"0b",
           756 => x"ea",
           757 => x"05",
           758 => x"05",
           759 => x"39",
           760 => x"8c",
           761 => x"e0",
           762 => x"08",
           763 => x"95",
           764 => x"82",
           765 => x"0c",
           766 => x"53",
           767 => x"52",
           768 => x"51",
           769 => x"70",
           770 => x"0d",
           771 => x"a4",
           772 => x"3d",
           773 => x"f8",
           774 => x"11",
           775 => x"70",
           776 => x"72",
           777 => x"e0",
           778 => x"39",
           779 => x"53",
           780 => x"05",
           781 => x"88",
           782 => x"08",
           783 => x"53",
           784 => x"fc",
           785 => x"e0",
           786 => x"11",
           787 => x"98",
           788 => x"38",
           789 => x"05",
           790 => x"08",
           791 => x"51",
           792 => x"e0",
           793 => x"38",
           794 => x"05",
           795 => x"08",
           796 => x"0c",
           797 => x"08",
           798 => x"82",
           799 => x"08",
           800 => x"0d",
           801 => x"05",
           802 => x"08",
           803 => x"81",
           804 => x"51",
           805 => x"0b",
           806 => x"80",
           807 => x"05",
           808 => x"08",
           809 => x"a4",
           810 => x"e0",
           811 => x"ff",
           812 => x"82",
           813 => x"e0",
           814 => x"e0",
           815 => x"11",
           816 => x"98",
           817 => x"38",
           818 => x"05",
           819 => x"08",
           820 => x"08",
           821 => x"08",
           822 => x"87",
           823 => x"82",
           824 => x"0c",
           825 => x"52",
           826 => x"51",
           827 => x"82",
           828 => x"82",
           829 => x"08",
           830 => x"0d",
           831 => x"85",
           832 => x"32",
           833 => x"53",
           834 => x"82",
           835 => x"cb",
           836 => x"08",
           837 => x"81",
           838 => x"2e",
           839 => x"8c",
           840 => x"05",
           841 => x"14",
           842 => x"08",
           843 => x"e0",
           844 => x"54",
           845 => x"05",
           846 => x"05",
           847 => x"12",
           848 => x"08",
           849 => x"0c",
           850 => x"a4",
           851 => x"08",
           852 => x"08",
           853 => x"53",
           854 => x"2d",
           855 => x"38",
           856 => x"8c",
           857 => x"82",
           858 => x"82",
           859 => x"53",
           860 => x"08",
           861 => x"fc",
           862 => x"3d",
           863 => x"e0",
           864 => x"f9",
           865 => x"05",
           866 => x"70",
           867 => x"80",
           868 => x"a4",
           869 => x"82",
           870 => x"11",
           871 => x"51",
           872 => x"c5",
           873 => x"08",
           874 => x"53",
           875 => x"06",
           876 => x"e0",
           877 => x"08",
           878 => x"a4",
           879 => x"70",
           880 => x"51",
           881 => x"a4",
           882 => x"70",
           883 => x"51",
           884 => x"82",
           885 => x"08",
           886 => x"05",
           887 => x"fc",
           888 => x"08",
           889 => x"88",
           890 => x"70",
           891 => x"34",
           892 => x"05",
           893 => x"08",
           894 => x"71",
           895 => x"a4",
           896 => x"08",
           897 => x"51",
           898 => x"70",
           899 => x"52",
           900 => x"80",
           901 => x"08",
           902 => x"f4",
           903 => x"05",
           904 => x"08",
           905 => x"08",
           906 => x"06",
           907 => x"05",
           908 => x"a4",
           909 => x"e0",
           910 => x"52",
           911 => x"34",
           912 => x"52",
           913 => x"85",
           914 => x"08",
           915 => x"a4",
           916 => x"81",
           917 => x"08",
           918 => x"70",
           919 => x"51",
           920 => x"05",
           921 => x"0d",
           922 => x"a4",
           923 => x"3d",
           924 => x"08",
           925 => x"82",
           926 => x"e0",
           927 => x"a4",
           928 => x"a2",
           929 => x"08",
           930 => x"26",
           931 => x"f8",
           932 => x"05",
           933 => x"fc",
           934 => x"82",
           935 => x"e0",
           936 => x"e0",
           937 => x"a4",
           938 => x"08",
           939 => x"08",
           940 => x"90",
           941 => x"08",
           942 => x"90",
           943 => x"08",
           944 => x"90",
           945 => x"82",
           946 => x"05",
           947 => x"82",
           948 => x"05",
           949 => x"82",
           950 => x"e0",
           951 => x"71",
           952 => x"e0",
           953 => x"82",
           954 => x"e0",
           955 => x"82",
           956 => x"e0",
           957 => x"ba",
           958 => x"08",
           959 => x"f8",
           960 => x"08",
           961 => x"fc",
           962 => x"82",
           963 => x"05",
           964 => x"ff",
           965 => x"05",
           966 => x"85",
           967 => x"82",
           968 => x"0c",
           969 => x"88",
           970 => x"05",
           971 => x"08",
           972 => x"fc",
           973 => x"08",
           974 => x"51",
           975 => x"39",
           976 => x"ff",
           977 => x"0c",
           978 => x"82",
           979 => x"70",
           980 => x"0d",
           981 => x"a4",
           982 => x"3d",
           983 => x"08",
           984 => x"82",
           985 => x"71",
           986 => x"08",
           987 => x"05",
           988 => x"08",
           989 => x"a4",
           990 => x"e0",
           991 => x"ff",
           992 => x"ff",
           993 => x"05",
           994 => x"84",
           995 => x"82",
           996 => x"0c",
           997 => x"88",
           998 => x"05",
           999 => x"08",
          1000 => x"82",
          1001 => x"2e",
          1002 => x"90",
          1003 => x"08",
          1004 => x"90",
          1005 => x"08",
          1006 => x"90",
          1007 => x"e0",
          1008 => x"33",
          1009 => x"81",
          1010 => x"0c",
          1011 => x"52",
          1012 => x"08",
          1013 => x"a4",
          1014 => x"82",
          1015 => x"82",
          1016 => x"82",
          1017 => x"08",
          1018 => x"0d",
          1019 => x"80",
          1020 => x"08",
          1021 => x"e0",
          1022 => x"82",
          1023 => x"e0",
          1024 => x"72",
          1025 => x"71",
          1026 => x"82",
          1027 => x"71",
          1028 => x"08",
          1029 => x"05",
          1030 => x"70",
          1031 => x"08",
          1032 => x"e0",
          1033 => x"82",
          1034 => x"e0",
          1035 => x"84",
          1036 => x"08",
          1037 => x"38",
          1038 => x"70",
          1039 => x"0b",
          1040 => x"80",
          1041 => x"05",
          1042 => x"8c",
          1043 => x"05",
          1044 => x"38",
          1045 => x"05",
          1046 => x"88",
          1047 => x"08",
          1048 => x"31",
          1049 => x"0c",
          1050 => x"80",
          1051 => x"0c",
          1052 => x"82",
          1053 => x"e0",
          1054 => x"02",
          1055 => x"82",
          1056 => x"82",
          1057 => x"81",
          1058 => x"82",
          1059 => x"e0",
          1060 => x"70",
          1061 => x"82",
          1062 => x"08",
          1063 => x"08",
          1064 => x"82",
          1065 => x"39",
          1066 => x"82",
          1067 => x"54",
          1068 => x"f8",
          1069 => x"88",
          1070 => x"fc",
          1071 => x"e0",
          1072 => x"f4",
          1073 => x"f4",
          1074 => x"3d",
          1075 => x"e0",
          1076 => x"fd",
          1077 => x"05",
          1078 => x"0c",
          1079 => x"8d",
          1080 => x"fc",
          1081 => x"a4",
          1082 => x"82",
          1083 => x"05",
          1084 => x"70",
          1085 => x"2e",
          1086 => x"05",
          1087 => x"8c",
          1088 => x"05",
          1089 => x"39",
          1090 => x"ff",
          1091 => x"0c",
          1092 => x"82",
          1093 => x"70",
          1094 => x"51",
          1095 => x"82",
          1096 => x"e0",
          1097 => x"02",
          1098 => x"82",
          1099 => x"e0",
          1100 => x"a4",
          1101 => x"d4",
          1102 => x"08",
          1103 => x"05",
          1104 => x"08",
          1105 => x"05",
          1106 => x"08",
          1107 => x"08",
          1108 => x"a4",
          1109 => x"71",
          1110 => x"08",
          1111 => x"05",
          1112 => x"08",
          1113 => x"0c",
          1114 => x"0c",
          1115 => x"e0",
          1116 => x"a4",
          1117 => x"a4",
          1118 => x"82",
          1119 => x"0c",
          1120 => x"0c",
          1121 => x"e0",
          1122 => x"82",
          1123 => x"e0",
          1124 => x"9b",
          1125 => x"08",
          1126 => x"08",
          1127 => x"0c",
          1128 => x"fc",
          1129 => x"05",
          1130 => x"08",
          1131 => x"08",
          1132 => x"82",
          1133 => x"e4",
          1134 => x"08",
          1135 => x"e0",
          1136 => x"a4",
          1137 => x"a4",
          1138 => x"08",
          1139 => x"f8",
          1140 => x"05",
          1141 => x"a4",
          1142 => x"80",
          1143 => x"0c",
          1144 => x"fc",
          1145 => x"e0",
          1146 => x"81",
          1147 => x"88",
          1148 => x"e8",
          1149 => x"e0",
          1150 => x"82",
          1151 => x"e0",
          1152 => x"a4",
          1153 => x"a4",
          1154 => x"08",
          1155 => x"f8",
          1156 => x"88",
          1157 => x"08",
          1158 => x"e0",
          1159 => x"a4",
          1160 => x"ab",
          1161 => x"08",
          1162 => x"08",
          1163 => x"05",
          1164 => x"e0",
          1165 => x"a4",
          1166 => x"e0",
          1167 => x"e0",
          1168 => x"a4",
          1169 => x"08",
          1170 => x"e0",
          1171 => x"71",
          1172 => x"05",
          1173 => x"08",
          1174 => x"05",
          1175 => x"08",
          1176 => x"06",
          1177 => x"71",
          1178 => x"0c",
          1179 => x"ff",
          1180 => x"0c",
          1181 => x"53",
          1182 => x"88",
          1183 => x"08",
          1184 => x"08",
          1185 => x"88",
          1186 => x"e8",
          1187 => x"08",
          1188 => x"8c",
          1189 => x"82",
          1190 => x"0c",
          1191 => x"88",
          1192 => x"05",
          1193 => x"08",
          1194 => x"38",
          1195 => x"05",
          1196 => x"a4",
          1197 => x"08",
          1198 => x"f8",
          1199 => x"08",
          1200 => x"08",
          1201 => x"a4",
          1202 => x"08",
          1203 => x"f4",
          1204 => x"05",
          1205 => x"70",
          1206 => x"08",
          1207 => x"82",
          1208 => x"e0",
          1209 => x"a4",
          1210 => x"e0",
          1211 => x"e0",
          1212 => x"82",
          1213 => x"e0",
          1214 => x"a4",
          1215 => x"a4",
          1216 => x"08",
          1217 => x"51",
          1218 => x"a4",
          1219 => x"0b",
          1220 => x"82",
          1221 => x"e0",
          1222 => x"82",
          1223 => x"82",
          1224 => x"2a",
          1225 => x"82",
          1226 => x"e0",
          1227 => x"e0",
          1228 => x"a4",
          1229 => x"51",
          1230 => x"a4",
          1231 => x"0b",
          1232 => x"82",
          1233 => x"e0",
          1234 => x"82",
          1235 => x"82",
          1236 => x"2a",
          1237 => x"82",
          1238 => x"e0",
          1239 => x"e0",
          1240 => x"82",
          1241 => x"82",
          1242 => x"2a",
          1243 => x"30",
          1244 => x"f4",
          1245 => x"98",
          1246 => x"52",
          1247 => x"a4",
          1248 => x"82",
          1249 => x"e0",
          1250 => x"e0",
          1251 => x"e4",
          1252 => x"e0",
          1253 => x"e0",
          1254 => x"70",
          1255 => x"84",
          1256 => x"82",
          1257 => x"0c",
          1258 => x"8c",
          1259 => x"88",
          1260 => x"98",
          1261 => x"84",
          1262 => x"82",
          1263 => x"0c",
          1264 => x"a4",
          1265 => x"08",
          1266 => x"82",
          1267 => x"fb",
          1268 => x"82",
          1269 => x"8f",
          1270 => x"08",
          1271 => x"82",
          1272 => x"2e",
          1273 => x"05",
          1274 => x"98",
          1275 => x"08",
          1276 => x"05",
          1277 => x"08",
          1278 => x"fc",
          1279 => x"e0",
          1280 => x"05",
          1281 => x"0c",
          1282 => x"ff",
          1283 => x"f8",
          1284 => x"a4",
          1285 => x"a4",
          1286 => x"39",
          1287 => x"ff",
          1288 => x"f8",
          1289 => x"38",
          1290 => x"05",
          1291 => x"08",
          1292 => x"a4",
          1293 => x"08",
          1294 => x"f8",
          1295 => x"f4",
          1296 => x"05",
          1297 => x"08",
          1298 => x"08",
          1299 => x"05",
          1300 => x"08",
          1301 => x"f8",
          1302 => x"82",
          1303 => x"82",
          1304 => x"05",
          1305 => x"71",
          1306 => x"08",
          1307 => x"88",
          1308 => x"08",
          1309 => x"08",
          1310 => x"8c",
          1311 => x"05",
          1312 => x"08",
          1313 => x"2c",
          1314 => x"82",
          1315 => x"06",
          1316 => x"82",
          1317 => x"e0",
          1318 => x"e0",
          1319 => x"82",
          1320 => x"e0",
          1321 => x"82",
          1322 => x"52",
          1323 => x"cb",
          1324 => x"08",
          1325 => x"0c",
          1326 => x"08",
          1327 => x"82",
          1328 => x"08",
          1329 => x"0d",
          1330 => x"05",
          1331 => x"08",
          1332 => x"2c",
          1333 => x"82",
          1334 => x"e0",
          1335 => x"e0",
          1336 => x"a4",
          1337 => x"08",
          1338 => x"a4",
          1339 => x"a4",
          1340 => x"08",
          1341 => x"f4",
          1342 => x"08",
          1343 => x"08",
          1344 => x"f8",
          1345 => x"05",
          1346 => x"05",
          1347 => x"08",
          1348 => x"08",
          1349 => x"e0",
          1350 => x"f8",
          1351 => x"08",
          1352 => x"98",
          1353 => x"82",
          1354 => x"08",
          1355 => x"0d",
          1356 => x"05",
          1357 => x"08",
          1358 => x"08",
          1359 => x"72",
          1360 => x"f8",
          1361 => x"72",
          1362 => x"82",
          1363 => x"08",
          1364 => x"82",
          1365 => x"72",
          1366 => x"81",
          1367 => x"34",
          1368 => x"70",
          1369 => x"51",
          1370 => x"f8",
          1371 => x"05",
          1372 => x"06",
          1373 => x"88",
          1374 => x"0c",
          1375 => x"e0",
          1376 => x"a4",
          1377 => x"08",
          1378 => x"e8",
          1379 => x"82",
          1380 => x"f8",
          1381 => x"0b",
          1382 => x"82",
          1383 => x"08",
          1384 => x"53",
          1385 => x"05",
          1386 => x"e0",
          1387 => x"a4",
          1388 => x"05",
          1389 => x"33",
          1390 => x"80",
          1391 => x"05",
          1392 => x"81",
          1393 => x"0c",
          1394 => x"f8",
          1395 => x"38",
          1396 => x"53",
          1397 => x"80",
          1398 => x"0c",
          1399 => x"a4",
          1400 => x"e0",
          1401 => x"73",
          1402 => x"f8",
          1403 => x"38",
          1404 => x"08",
          1405 => x"0b",
          1406 => x"80",
          1407 => x"0c",
          1408 => x"53",
          1409 => x"e0",
          1410 => x"e0",
          1411 => x"08",
          1412 => x"72",
          1413 => x"82",
          1414 => x"11",
          1415 => x"f8",
          1416 => x"05",
          1417 => x"82",
          1418 => x"11",
          1419 => x"f8",
          1420 => x"05",
          1421 => x"80",
          1422 => x"0c",
          1423 => x"f8",
          1424 => x"05",
          1425 => x"38",
          1426 => x"05",
          1427 => x"08",
          1428 => x"08",
          1429 => x"08",
          1430 => x"a4",
          1431 => x"08",
          1432 => x"71",
          1433 => x"53",
          1434 => x"05",
          1435 => x"08",
          1436 => x"90",
          1437 => x"08",
          1438 => x"0c",
          1439 => x"82",
          1440 => x"0c",
          1441 => x"ec",
          1442 => x"05",
          1443 => x"0d",
          1444 => x"a4",
          1445 => x"3d",
          1446 => x"f0",
          1447 => x"05",
          1448 => x"a4",
          1449 => x"53",
          1450 => x"08",
          1451 => x"53",
          1452 => x"38",
          1453 => x"70",
          1454 => x"39",
          1455 => x"53",
          1456 => x"38",
          1457 => x"05",
          1458 => x"08",
          1459 => x"08",
          1460 => x"08",
          1461 => x"f8",
          1462 => x"81",
          1463 => x"08",
          1464 => x"71",
          1465 => x"82",
          1466 => x"e0",
          1467 => x"a4",
          1468 => x"08",
          1469 => x"38",
          1470 => x"80",
          1471 => x"90",
          1472 => x"34",
          1473 => x"70",
          1474 => x"51",
          1475 => x"f8",
          1476 => x"82",
          1477 => x"e0",
          1478 => x"81",
          1479 => x"72",
          1480 => x"34",
          1481 => x"f8",
          1482 => x"38",
          1483 => x"05",
          1484 => x"08",
          1485 => x"90",
          1486 => x"33",
          1487 => x"39",
          1488 => x"05",
          1489 => x"e0",
          1490 => x"82",
          1491 => x"af",
          1492 => x"08",
          1493 => x"83",
          1494 => x"a4",
          1495 => x"8a",
          1496 => x"34",
          1497 => x"05",
          1498 => x"33",
          1499 => x"82",
          1500 => x"80",
          1501 => x"a4",
          1502 => x"53",
          1503 => x"34",
          1504 => x"d0",
          1505 => x"08",
          1506 => x"f8",
          1507 => x"38",
          1508 => x"f9",
          1509 => x"08",
          1510 => x"f8",
          1511 => x"38",
          1512 => x"05",
          1513 => x"08",
          1514 => x"f4",
          1515 => x"8d",
          1516 => x"ec",
          1517 => x"a4",
          1518 => x"a4",
          1519 => x"a4",
          1520 => x"e0",
          1521 => x"a4",
          1522 => x"05",
          1523 => x"55",
          1524 => x"f8",
          1525 => x"a4",
          1526 => x"2e",
          1527 => x"05",
          1528 => x"05",
          1529 => x"08",
          1530 => x"71",
          1531 => x"08",
          1532 => x"ec",
          1533 => x"3d",
          1534 => x"3d",
          1535 => x"59",
          1536 => x"39",
          1537 => x"54",
          1538 => x"a0",
          1539 => x"15",
          1540 => x"29",
          1541 => x"56",
          1542 => x"82",
          1543 => x"08",
          1544 => x"98",
          1545 => x"73",
          1546 => x"70",
          1547 => x"27",
          1548 => x"98",
          1549 => x"0b",
          1550 => x"0d",
          1551 => x"38",
          1552 => x"52",
          1553 => x"81",
          1554 => x"f9",
          1555 => x"39",
          1556 => x"82",
          1557 => x"be",
          1558 => x"c4",
          1559 => x"51",
          1560 => x"80",
          1561 => x"c1",
          1562 => x"82",
          1563 => x"cc",
          1564 => x"a9",
          1565 => x"82",
          1566 => x"b4",
          1567 => x"91",
          1568 => x"82",
          1569 => x"88",
          1570 => x"04",
          1571 => x"74",
          1572 => x"75",
          1573 => x"e8",
          1574 => x"e0",
          1575 => x"3f",
          1576 => x"75",
          1577 => x"c2",
          1578 => x"0d",
          1579 => x"33",
          1580 => x"7a",
          1581 => x"78",
          1582 => x"81",
          1583 => x"06",
          1584 => x"38",
          1585 => x"52",
          1586 => x"98",
          1587 => x"38",
          1588 => x"88",
          1589 => x"3d",
          1590 => x"52",
          1591 => x"e0",
          1592 => x"90",
          1593 => x"38",
          1594 => x"39",
          1595 => x"cd",
          1596 => x"25",
          1597 => x"51",
          1598 => x"38",
          1599 => x"88",
          1600 => x"76",
          1601 => x"3d",
          1602 => x"84",
          1603 => x"58",
          1604 => x"ad",
          1605 => x"76",
          1606 => x"9c",
          1607 => x"61",
          1608 => x"7f",
          1609 => x"98",
          1610 => x"82",
          1611 => x"f3",
          1612 => x"05",
          1613 => x"68",
          1614 => x"77",
          1615 => x"98",
          1616 => x"72",
          1617 => x"80",
          1618 => x"53",
          1619 => x"82",
          1620 => x"82",
          1621 => x"80",
          1622 => x"7b",
          1623 => x"a7",
          1624 => x"72",
          1625 => x"82",
          1626 => x"89",
          1627 => x"b2",
          1628 => x"74",
          1629 => x"72",
          1630 => x"ae",
          1631 => x"51",
          1632 => x"a1",
          1633 => x"8e",
          1634 => x"51",
          1635 => x"c1",
          1636 => x"15",
          1637 => x"51",
          1638 => x"c1",
          1639 => x"55",
          1640 => x"19",
          1641 => x"7a",
          1642 => x"9f",
          1643 => x"73",
          1644 => x"72",
          1645 => x"26",
          1646 => x"73",
          1647 => x"52",
          1648 => x"55",
          1649 => x"c9",
          1650 => x"59",
          1651 => x"98",
          1652 => x"57",
          1653 => x"38",
          1654 => x"98",
          1655 => x"a0",
          1656 => x"30",
          1657 => x"51",
          1658 => x"73",
          1659 => x"b6",
          1660 => x"fd",
          1661 => x"98",
          1662 => x"0d",
          1663 => x"cb",
          1664 => x"c1",
          1665 => x"de",
          1666 => x"c2",
          1667 => x"de",
          1668 => x"ff",
          1669 => x"38",
          1670 => x"fe",
          1671 => x"53",
          1672 => x"3f",
          1673 => x"80",
          1674 => x"70",
          1675 => x"92",
          1676 => x"c2",
          1677 => x"99",
          1678 => x"06",
          1679 => x"81",
          1680 => x"51",
          1681 => x"3f",
          1682 => x"52",
          1683 => x"98",
          1684 => x"fa",
          1685 => x"84",
          1686 => x"80",
          1687 => x"3f",
          1688 => x"80",
          1689 => x"70",
          1690 => x"92",
          1691 => x"c3",
          1692 => x"98",
          1693 => x"06",
          1694 => x"81",
          1695 => x"51",
          1696 => x"3f",
          1697 => x"52",
          1698 => x"97",
          1699 => x"82",
          1700 => x"88",
          1701 => x"80",
          1702 => x"3f",
          1703 => x"80",
          1704 => x"84",
          1705 => x"02",
          1706 => x"56",
          1707 => x"3f",
          1708 => x"73",
          1709 => x"52",
          1710 => x"3f",
          1711 => x"e0",
          1712 => x"31",
          1713 => x"db",
          1714 => x"33",
          1715 => x"af",
          1716 => x"75",
          1717 => x"98",
          1718 => x"98",
          1719 => x"82",
          1720 => x"82",
          1721 => x"0b",
          1722 => x"82",
          1723 => x"c4",
          1724 => x"f0",
          1725 => x"87",
          1726 => x"70",
          1727 => x"0c",
          1728 => x"8a",
          1729 => x"06",
          1730 => x"a3",
          1731 => x"c4",
          1732 => x"7d",
          1733 => x"81",
          1734 => x"7e",
          1735 => x"8d",
          1736 => x"c4",
          1737 => x"3d",
          1738 => x"51",
          1739 => x"05",
          1740 => x"08",
          1741 => x"78",
          1742 => x"80",
          1743 => x"81",
          1744 => x"78",
          1745 => x"2e",
          1746 => x"80",
          1747 => x"c0",
          1748 => x"82",
          1749 => x"f9",
          1750 => x"24",
          1751 => x"8d",
          1752 => x"38",
          1753 => x"8a",
          1754 => x"38",
          1755 => x"8a",
          1756 => x"83",
          1757 => x"80",
          1758 => x"ad",
          1759 => x"fe",
          1760 => x"53",
          1761 => x"82",
          1762 => x"38",
          1763 => x"84",
          1764 => x"98",
          1765 => x"43",
          1766 => x"3f",
          1767 => x"81",
          1768 => x"84",
          1769 => x"38",
          1770 => x"11",
          1771 => x"3f",
          1772 => x"de",
          1773 => x"ff",
          1774 => x"e0",
          1775 => x"b5",
          1776 => x"05",
          1777 => x"08",
          1778 => x"f8",
          1779 => x"79",
          1780 => x"79",
          1781 => x"62",
          1782 => x"ff",
          1783 => x"ea",
          1784 => x"2e",
          1785 => x"11",
          1786 => x"3f",
          1787 => x"e6",
          1788 => x"ff",
          1789 => x"e0",
          1790 => x"82",
          1791 => x"64",
          1792 => x"70",
          1793 => x"7c",
          1794 => x"79",
          1795 => x"51",
          1796 => x"81",
          1797 => x"c3",
          1798 => x"ff",
          1799 => x"e9",
          1800 => x"df",
          1801 => x"80",
          1802 => x"45",
          1803 => x"59",
          1804 => x"bc",
          1805 => x"33",
          1806 => x"de",
          1807 => x"ff",
          1808 => x"82",
          1809 => x"de",
          1810 => x"38",
          1811 => x"82",
          1812 => x"b5",
          1813 => x"05",
          1814 => x"08",
          1815 => x"59",
          1816 => x"b8",
          1817 => x"fd",
          1818 => x"82",
          1819 => x"de",
          1820 => x"38",
          1821 => x"82",
          1822 => x"88",
          1823 => x"39",
          1824 => x"2e",
          1825 => x"88",
          1826 => x"44",
          1827 => x"84",
          1828 => x"98",
          1829 => x"5c",
          1830 => x"5c",
          1831 => x"07",
          1832 => x"5a",
          1833 => x"a0",
          1834 => x"b0",
          1835 => x"64",
          1836 => x"f1",
          1837 => x"b6",
          1838 => x"ff",
          1839 => x"e0",
          1840 => x"b5",
          1841 => x"05",
          1842 => x"08",
          1843 => x"80",
          1844 => x"05",
          1845 => x"ff",
          1846 => x"e0",
          1847 => x"64",
          1848 => x"51",
          1849 => x"08",
          1850 => x"a1",
          1851 => x"78",
          1852 => x"27",
          1853 => x"53",
          1854 => x"82",
          1855 => x"64",
          1856 => x"34",
          1857 => x"82",
          1858 => x"ff",
          1859 => x"53",
          1860 => x"82",
          1861 => x"38",
          1862 => x"84",
          1863 => x"98",
          1864 => x"02",
          1865 => x"05",
          1866 => x"f0",
          1867 => x"f4",
          1868 => x"f7",
          1869 => x"82",
          1870 => x"82",
          1871 => x"79",
          1872 => x"79",
          1873 => x"38",
          1874 => x"05",
          1875 => x"11",
          1876 => x"3f",
          1877 => x"38",
          1878 => x"79",
          1879 => x"ff",
          1880 => x"ba",
          1881 => x"fe",
          1882 => x"de",
          1883 => x"2e",
          1884 => x"11",
          1885 => x"3f",
          1886 => x"38",
          1887 => x"05",
          1888 => x"ff",
          1889 => x"e0",
          1890 => x"61",
          1891 => x"51",
          1892 => x"08",
          1893 => x"9e",
          1894 => x"78",
          1895 => x"27",
          1896 => x"53",
          1897 => x"82",
          1898 => x"61",
          1899 => x"42",
          1900 => x"ff",
          1901 => x"3d",
          1902 => x"51",
          1903 => x"80",
          1904 => x"c5",
          1905 => x"59",
          1906 => x"53",
          1907 => x"82",
          1908 => x"38",
          1909 => x"9c",
          1910 => x"e0",
          1911 => x"82",
          1912 => x"51",
          1913 => x"82",
          1914 => x"ff",
          1915 => x"c6",
          1916 => x"59",
          1917 => x"d6",
          1918 => x"2e",
          1919 => x"51",
          1920 => x"5d",
          1921 => x"92",
          1922 => x"3d",
          1923 => x"82",
          1924 => x"5c",
          1925 => x"e0",
          1926 => x"e0",
          1927 => x"81",
          1928 => x"82",
          1929 => x"38",
          1930 => x"38",
          1931 => x"7b",
          1932 => x"82",
          1933 => x"05",
          1934 => x"7b",
          1935 => x"c4",
          1936 => x"c6",
          1937 => x"52",
          1938 => x"9d",
          1939 => x"53",
          1940 => x"b0",
          1941 => x"de",
          1942 => x"56",
          1943 => x"53",
          1944 => x"b0",
          1945 => x"98",
          1946 => x"30",
          1947 => x"5b",
          1948 => x"38",
          1949 => x"80",
          1950 => x"ff",
          1951 => x"7f",
          1952 => x"78",
          1953 => x"06",
          1954 => x"b6",
          1955 => x"f2",
          1956 => x"b5",
          1957 => x"0d",
          1958 => x"c0",
          1959 => x"84",
          1960 => x"82",
          1961 => x"55",
          1962 => x"cb",
          1963 => x"07",
          1964 => x"08",
          1965 => x"51",
          1966 => x"90",
          1967 => x"80",
          1968 => x"82",
          1969 => x"80",
          1970 => x"8c",
          1971 => x"0c",
          1972 => x"5b",
          1973 => x"80",
          1974 => x"70",
          1975 => x"fb",
          1976 => x"ee",
          1977 => x"cd",
          1978 => x"c5",
          1979 => x"3f",
          1980 => x"3f",
          1981 => x"08",
          1982 => x"74",
          1983 => x"70",
          1984 => x"81",
          1985 => x"70",
          1986 => x"81",
          1987 => x"81",
          1988 => x"39",
          1989 => x"54",
          1990 => x"70",
          1991 => x"98",
          1992 => x"52",
          1993 => x"54",
          1994 => x"38",
          1995 => x"2e",
          1996 => x"70",
          1997 => x"76",
          1998 => x"88",
          1999 => x"34",
          2000 => x"e0",
          2001 => x"3d",
          2002 => x"91",
          2003 => x"51",
          2004 => x"85",
          2005 => x"72",
          2006 => x"04",
          2007 => x"ff",
          2008 => x"26",
          2009 => x"05",
          2010 => x"8a",
          2011 => x"70",
          2012 => x"33",
          2013 => x"f2",
          2014 => x"70",
          2015 => x"22",
          2016 => x"80",
          2017 => x"52",
          2018 => x"81",
          2019 => x"22",
          2020 => x"33",
          2021 => x"33",
          2022 => x"33",
          2023 => x"33",
          2024 => x"33",
          2025 => x"c0",
          2026 => x"a0",
          2027 => x"0c",
          2028 => x"86",
          2029 => x"5b",
          2030 => x"0c",
          2031 => x"7b",
          2032 => x"79",
          2033 => x"08",
          2034 => x"98",
          2035 => x"87",
          2036 => x"1c",
          2037 => x"79",
          2038 => x"08",
          2039 => x"98",
          2040 => x"80",
          2041 => x"59",
          2042 => x"1b",
          2043 => x"1b",
          2044 => x"1b",
          2045 => x"52",
          2046 => x"3f",
          2047 => x"02",
          2048 => x"81",
          2049 => x"52",
          2050 => x"25",
          2051 => x"2e",
          2052 => x"84",
          2053 => x"2b",
          2054 => x"2e",
          2055 => x"72",
          2056 => x"72",
          2057 => x"80",
          2058 => x"ff",
          2059 => x"85",
          2060 => x"53",
          2061 => x"51",
          2062 => x"98",
          2063 => x"16",
          2064 => x"38",
          2065 => x"0d",
          2066 => x"33",
          2067 => x"06",
          2068 => x"51",
          2069 => x"94",
          2070 => x"70",
          2071 => x"2e",
          2072 => x"06",
          2073 => x"32",
          2074 => x"2e",
          2075 => x"06",
          2076 => x"81",
          2077 => x"52",
          2078 => x"94",
          2079 => x"e0",
          2080 => x"3d",
          2081 => x"70",
          2082 => x"de",
          2083 => x"3d",
          2084 => x"8a",
          2085 => x"52",
          2086 => x"33",
          2087 => x"c0",
          2088 => x"38",
          2089 => x"70",
          2090 => x"54",
          2091 => x"2a",
          2092 => x"38",
          2093 => x"53",
          2094 => x"2a",
          2095 => x"be",
          2096 => x"c0",
          2097 => x"38",
          2098 => x"0c",
          2099 => x"3d",
          2100 => x"80",
          2101 => x"53",
          2102 => x"71",
          2103 => x"b0",
          2104 => x"55",
          2105 => x"80",
          2106 => x"51",
          2107 => x"06",
          2108 => x"38",
          2109 => x"51",
          2110 => x"81",
          2111 => x"38",
          2112 => x"51",
          2113 => x"06",
          2114 => x"80",
          2115 => x"52",
          2116 => x"70",
          2117 => x"ff",
          2118 => x"89",
          2119 => x"de",
          2120 => x"52",
          2121 => x"2e",
          2122 => x"70",
          2123 => x"51",
          2124 => x"71",
          2125 => x"80",
          2126 => x"c0",
          2127 => x"ff",
          2128 => x"3d",
          2129 => x"98",
          2130 => x"0c",
          2131 => x"33",
          2132 => x"c0",
          2133 => x"38",
          2134 => x"70",
          2135 => x"51",
          2136 => x"72",
          2137 => x"80",
          2138 => x"c0",
          2139 => x"2b",
          2140 => x"82",
          2141 => x"ff",
          2142 => x"70",
          2143 => x"80",
          2144 => x"a4",
          2145 => x"9e",
          2146 => x"c0",
          2147 => x"87",
          2148 => x"0c",
          2149 => x"c4",
          2150 => x"de",
          2151 => x"82",
          2152 => x"08",
          2153 => x"b4",
          2154 => x"9e",
          2155 => x"c0",
          2156 => x"87",
          2157 => x"0c",
          2158 => x"e4",
          2159 => x"70",
          2160 => x"84",
          2161 => x"9e",
          2162 => x"c0",
          2163 => x"81",
          2164 => x"87",
          2165 => x"0a",
          2166 => x"83",
          2167 => x"34",
          2168 => x"70",
          2169 => x"70",
          2170 => x"82",
          2171 => x"9e",
          2172 => x"51",
          2173 => x"81",
          2174 => x"0b",
          2175 => x"80",
          2176 => x"2e",
          2177 => x"fc",
          2178 => x"08",
          2179 => x"52",
          2180 => x"71",
          2181 => x"c0",
          2182 => x"06",
          2183 => x"38",
          2184 => x"80",
          2185 => x"84",
          2186 => x"80",
          2187 => x"de",
          2188 => x"90",
          2189 => x"52",
          2190 => x"52",
          2191 => x"87",
          2192 => x"80",
          2193 => x"83",
          2194 => x"34",
          2195 => x"70",
          2196 => x"70",
          2197 => x"82",
          2198 => x"9e",
          2199 => x"52",
          2200 => x"52",
          2201 => x"9e",
          2202 => x"8a",
          2203 => x"84",
          2204 => x"08",
          2205 => x"70",
          2206 => x"82",
          2207 => x"08",
          2208 => x"51",
          2209 => x"80",
          2210 => x"88",
          2211 => x"83",
          2212 => x"34",
          2213 => x"06",
          2214 => x"83",
          2215 => x"c8",
          2216 => x"de",
          2217 => x"38",
          2218 => x"3f",
          2219 => x"3f",
          2220 => x"2e",
          2221 => x"de",
          2222 => x"dc",
          2223 => x"ff",
          2224 => x"82",
          2225 => x"11",
          2226 => x"88",
          2227 => x"73",
          2228 => x"08",
          2229 => x"82",
          2230 => x"82",
          2231 => x"94",
          2232 => x"c0",
          2233 => x"51",
          2234 => x"33",
          2235 => x"de",
          2236 => x"54",
          2237 => x"a2",
          2238 => x"80",
          2239 => x"52",
          2240 => x"3f",
          2241 => x"2e",
          2242 => x"82",
          2243 => x"82",
          2244 => x"8e",
          2245 => x"ca",
          2246 => x"de",
          2247 => x"38",
          2248 => x"3f",
          2249 => x"2e",
          2250 => x"a3",
          2251 => x"73",
          2252 => x"51",
          2253 => x"33",
          2254 => x"ca",
          2255 => x"df",
          2256 => x"38",
          2257 => x"3f",
          2258 => x"3f",
          2259 => x"90",
          2260 => x"e0",
          2261 => x"86",
          2262 => x"82",
          2263 => x"82",
          2264 => x"82",
          2265 => x"51",
          2266 => x"08",
          2267 => x"ff",
          2268 => x"bd",
          2269 => x"54",
          2270 => x"b8",
          2271 => x"ff",
          2272 => x"82",
          2273 => x"52",
          2274 => x"e0",
          2275 => x"71",
          2276 => x"52",
          2277 => x"3f",
          2278 => x"2e",
          2279 => x"bd",
          2280 => x"91",
          2281 => x"c0",
          2282 => x"e0",
          2283 => x"ff",
          2284 => x"d7",
          2285 => x"0d",
          2286 => x"71",
          2287 => x"82",
          2288 => x"82",
          2289 => x"c4",
          2290 => x"91",
          2291 => x"82",
          2292 => x"e0",
          2293 => x"0d",
          2294 => x"0b",
          2295 => x"df",
          2296 => x"04",
          2297 => x"98",
          2298 => x"72",
          2299 => x"51",
          2300 => x"ec",
          2301 => x"9c",
          2302 => x"02",
          2303 => x"52",
          2304 => x"06",
          2305 => x"98",
          2306 => x"0d",
          2307 => x"71",
          2308 => x"b1",
          2309 => x"51",
          2310 => x"08",
          2311 => x"82",
          2312 => x"a3",
          2313 => x"72",
          2314 => x"cc",
          2315 => x"74",
          2316 => x"3d",
          2317 => x"33",
          2318 => x"df",
          2319 => x"90",
          2320 => x"58",
          2321 => x"51",
          2322 => x"70",
          2323 => x"19",
          2324 => x"3f",
          2325 => x"df",
          2326 => x"90",
          2327 => x"80",
          2328 => x"74",
          2329 => x"e8",
          2330 => x"e8",
          2331 => x"75",
          2332 => x"e8",
          2333 => x"df",
          2334 => x"38",
          2335 => x"38",
          2336 => x"78",
          2337 => x"82",
          2338 => x"a2",
          2339 => x"80",
          2340 => x"fd",
          2341 => x"54",
          2342 => x"38",
          2343 => x"0c",
          2344 => x"80",
          2345 => x"e8",
          2346 => x"80",
          2347 => x"cd",
          2348 => x"a7",
          2349 => x"85",
          2350 => x"57",
          2351 => x"80",
          2352 => x"80",
          2353 => x"80",
          2354 => x"81",
          2355 => x"80",
          2356 => x"97",
          2357 => x"0b",
          2358 => x"82",
          2359 => x"55",
          2360 => x"52",
          2361 => x"ff",
          2362 => x"81",
          2363 => x"04",
          2364 => x"3d",
          2365 => x"80",
          2366 => x"f4",
          2367 => x"95",
          2368 => x"54",
          2369 => x"52",
          2370 => x"98",
          2371 => x"ff",
          2372 => x"81",
          2373 => x"98",
          2374 => x"08",
          2375 => x"74",
          2376 => x"07",
          2377 => x"2e",
          2378 => x"df",
          2379 => x"80",
          2380 => x"80",
          2381 => x"fe",
          2382 => x"81",
          2383 => x"ff",
          2384 => x"b7",
          2385 => x"98",
          2386 => x"e0",
          2387 => x"3d",
          2388 => x"33",
          2389 => x"09",
          2390 => x"05",
          2391 => x"17",
          2392 => x"55",
          2393 => x"38",
          2394 => x"73",
          2395 => x"08",
          2396 => x"e0",
          2397 => x"51",
          2398 => x"08",
          2399 => x"74",
          2400 => x"88",
          2401 => x"39",
          2402 => x"53",
          2403 => x"e0",
          2404 => x"1b",
          2405 => x"3f",
          2406 => x"55",
          2407 => x"81",
          2408 => x"82",
          2409 => x"73",
          2410 => x"04",
          2411 => x"3d",
          2412 => x"80",
          2413 => x"33",
          2414 => x"81",
          2415 => x"55",
          2416 => x"80",
          2417 => x"06",
          2418 => x"38",
          2419 => x"98",
          2420 => x"98",
          2421 => x"53",
          2422 => x"80",
          2423 => x"80",
          2424 => x"ff",
          2425 => x"e0",
          2426 => x"53",
          2427 => x"54",
          2428 => x"08",
          2429 => x"09",
          2430 => x"98",
          2431 => x"e0",
          2432 => x"98",
          2433 => x"08",
          2434 => x"74",
          2435 => x"52",
          2436 => x"70",
          2437 => x"27",
          2438 => x"09",
          2439 => x"75",
          2440 => x"82",
          2441 => x"f9",
          2442 => x"e7",
          2443 => x"2b",
          2444 => x"2e",
          2445 => x"f7",
          2446 => x"2c",
          2447 => x"70",
          2448 => x"84",
          2449 => x"15",
          2450 => x"59",
          2451 => x"78",
          2452 => x"b4",
          2453 => x"ff",
          2454 => x"80",
          2455 => x"74",
          2456 => x"e0",
          2457 => x"80",
          2458 => x"34",
          2459 => x"0a",
          2460 => x"2c",
          2461 => x"73",
          2462 => x"52",
          2463 => x"98",
          2464 => x"38",
          2465 => x"80",
          2466 => x"f7",
          2467 => x"2c",
          2468 => x"70",
          2469 => x"2b",
          2470 => x"51",
          2471 => x"2e",
          2472 => x"cd",
          2473 => x"82",
          2474 => x"d0",
          2475 => x"34",
          2476 => x"3d",
          2477 => x"95",
          2478 => x"82",
          2479 => x"82",
          2480 => x"fd",
          2481 => x"73",
          2482 => x"70",
          2483 => x"9e",
          2484 => x"15",
          2485 => x"ff",
          2486 => x"dc",
          2487 => x"f7",
          2488 => x"82",
          2489 => x"3d",
          2490 => x"54",
          2491 => x"54",
          2492 => x"dc",
          2493 => x"ff",
          2494 => x"d8",
          2495 => x"25",
          2496 => x"74",
          2497 => x"dc",
          2498 => x"80",
          2499 => x"d8",
          2500 => x"da",
          2501 => x"2b",
          2502 => x"5a",
          2503 => x"92",
          2504 => x"51",
          2505 => x"0a",
          2506 => x"2c",
          2507 => x"73",
          2508 => x"83",
          2509 => x"82",
          2510 => x"b8",
          2511 => x"82",
          2512 => x"55",
          2513 => x"82",
          2514 => x"82",
          2515 => x"82",
          2516 => x"52",
          2517 => x"f7",
          2518 => x"2c",
          2519 => x"57",
          2520 => x"54",
          2521 => x"fc",
          2522 => x"94",
          2523 => x"80",
          2524 => x"d8",
          2525 => x"d5",
          2526 => x"51",
          2527 => x"33",
          2528 => x"f7",
          2529 => x"74",
          2530 => x"08",
          2531 => x"74",
          2532 => x"05",
          2533 => x"58",
          2534 => x"fa",
          2535 => x"05",
          2536 => x"08",
          2537 => x"82",
          2538 => x"3f",
          2539 => x"54",
          2540 => x"54",
          2541 => x"73",
          2542 => x"39",
          2543 => x"dc",
          2544 => x"79",
          2545 => x"04",
          2546 => x"2e",
          2547 => x"52",
          2548 => x"f7",
          2549 => x"f7",
          2550 => x"dd",
          2551 => x"d8",
          2552 => x"8a",
          2553 => x"d8",
          2554 => x"75",
          2555 => x"74",
          2556 => x"14",
          2557 => x"52",
          2558 => x"74",
          2559 => x"05",
          2560 => x"58",
          2561 => x"82",
          2562 => x"93",
          2563 => x"98",
          2564 => x"33",
          2565 => x"f8",
          2566 => x"88",
          2567 => x"80",
          2568 => x"98",
          2569 => x"55",
          2570 => x"39",
          2571 => x"06",
          2572 => x"74",
          2573 => x"fc",
          2574 => x"f7",
          2575 => x"54",
          2576 => x"33",
          2577 => x"33",
          2578 => x"38",
          2579 => x"80",
          2580 => x"3f",
          2581 => x"0b",
          2582 => x"7a",
          2583 => x"74",
          2584 => x"9a",
          2585 => x"f7",
          2586 => x"ff",
          2587 => x"51",
          2588 => x"c0",
          2589 => x"05",
          2590 => x"2e",
          2591 => x"3f",
          2592 => x"34",
          2593 => x"81",
          2594 => x"9c",
          2595 => x"39",
          2596 => x"aa",
          2597 => x"99",
          2598 => x"ae",
          2599 => x"80",
          2600 => x"f7",
          2601 => x"d8",
          2602 => x"06",
          2603 => x"ff",
          2604 => x"84",
          2605 => x"56",
          2606 => x"51",
          2607 => x"08",
          2608 => x"08",
          2609 => x"52",
          2610 => x"1b",
          2611 => x"39",
          2612 => x"34",
          2613 => x"33",
          2614 => x"9a",
          2615 => x"ff",
          2616 => x"54",
          2617 => x"fb",
          2618 => x"82",
          2619 => x"52",
          2620 => x"39",
          2621 => x"2e",
          2622 => x"52",
          2623 => x"f7",
          2624 => x"f7",
          2625 => x"0d",
          2626 => x"0c",
          2627 => x"82",
          2628 => x"f4",
          2629 => x"88",
          2630 => x"81",
          2631 => x"88",
          2632 => x"85",
          2633 => x"77",
          2634 => x"82",
          2635 => x"ff",
          2636 => x"ff",
          2637 => x"55",
          2638 => x"17",
          2639 => x"29",
          2640 => x"51",
          2641 => x"83",
          2642 => x"3d",
          2643 => x"27",
          2644 => x"11",
          2645 => x"51",
          2646 => x"0d",
          2647 => x"22",
          2648 => x"05",
          2649 => x"71",
          2650 => x"33",
          2651 => x"02",
          2652 => x"ff",
          2653 => x"51",
          2654 => x"54",
          2655 => x"34",
          2656 => x"2a",
          2657 => x"83",
          2658 => x"17",
          2659 => x"2b",
          2660 => x"06",
          2661 => x"83",
          2662 => x"54",
          2663 => x"ff",
          2664 => x"e0",
          2665 => x"72",
          2666 => x"fb",
          2667 => x"84",
          2668 => x"72",
          2669 => x"71",
          2670 => x"5b",
          2671 => x"12",
          2672 => x"07",
          2673 => x"70",
          2674 => x"82",
          2675 => x"33",
          2676 => x"83",
          2677 => x"05",
          2678 => x"88",
          2679 => x"56",
          2680 => x"13",
          2681 => x"33",
          2682 => x"70",
          2683 => x"53",
          2684 => x"70",
          2685 => x"fa",
          2686 => x"e0",
          2687 => x"70",
          2688 => x"07",
          2689 => x"12",
          2690 => x"07",
          2691 => x"57",
          2692 => x"38",
          2693 => x"88",
          2694 => x"33",
          2695 => x"74",
          2696 => x"88",
          2697 => x"f8",
          2698 => x"58",
          2699 => x"52",
          2700 => x"34",
          2701 => x"33",
          2702 => x"83",
          2703 => x"05",
          2704 => x"2b",
          2705 => x"88",
          2706 => x"74",
          2707 => x"0d",
          2708 => x"08",
          2709 => x"83",
          2710 => x"12",
          2711 => x"07",
          2712 => x"05",
          2713 => x"2b",
          2714 => x"71",
          2715 => x"53",
          2716 => x"34",
          2717 => x"33",
          2718 => x"83",
          2719 => x"05",
          2720 => x"88",
          2721 => x"56",
          2722 => x"13",
          2723 => x"11",
          2724 => x"07",
          2725 => x"3d",
          2726 => x"e0",
          2727 => x"ff",
          2728 => x"a7",
          2729 => x"2b",
          2730 => x"33",
          2731 => x"75",
          2732 => x"98",
          2733 => x"40",
          2734 => x"72",
          2735 => x"52",
          2736 => x"39",
          2737 => x"8b",
          2738 => x"79",
          2739 => x"76",
          2740 => x"56",
          2741 => x"08",
          2742 => x"33",
          2743 => x"54",
          2744 => x"34",
          2745 => x"08",
          2746 => x"80",
          2747 => x"08",
          2748 => x"14",
          2749 => x"33",
          2750 => x"70",
          2751 => x"53",
          2752 => x"72",
          2753 => x"ff",
          2754 => x"08",
          2755 => x"2e",
          2756 => x"83",
          2757 => x"7e",
          2758 => x"98",
          2759 => x"88",
          2760 => x"71",
          2761 => x"58",
          2762 => x"2e",
          2763 => x"70",
          2764 => x"07",
          2765 => x"70",
          2766 => x"52",
          2767 => x"27",
          2768 => x"75",
          2769 => x"16",
          2770 => x"75",
          2771 => x"85",
          2772 => x"83",
          2773 => x"33",
          2774 => x"70",
          2775 => x"56",
          2776 => x"81",
          2777 => x"cc",
          2778 => x"c4",
          2779 => x"89",
          2780 => x"ac",
          2781 => x"75",
          2782 => x"08",
          2783 => x"33",
          2784 => x"53",
          2785 => x"70",
          2786 => x"5c",
          2787 => x"76",
          2788 => x"34",
          2789 => x"71",
          2790 => x"12",
          2791 => x"2a",
          2792 => x"73",
          2793 => x"82",
          2794 => x"33",
          2795 => x"83",
          2796 => x"05",
          2797 => x"15",
          2798 => x"71",
          2799 => x"71",
          2800 => x"5a",
          2801 => x"34",
          2802 => x"08",
          2803 => x"98",
          2804 => x"0d",
          2805 => x"38",
          2806 => x"2e",
          2807 => x"82",
          2808 => x"98",
          2809 => x"0d",
          2810 => x"40",
          2811 => x"81",
          2812 => x"8e",
          2813 => x"e0",
          2814 => x"8b",
          2815 => x"54",
          2816 => x"3f",
          2817 => x"06",
          2818 => x"83",
          2819 => x"83",
          2820 => x"33",
          2821 => x"70",
          2822 => x"fc",
          2823 => x"81",
          2824 => x"90",
          2825 => x"52",
          2826 => x"5b",
          2827 => x"ff",
          2828 => x"ff",
          2829 => x"17",
          2830 => x"29",
          2831 => x"98",
          2832 => x"45",
          2833 => x"38",
          2834 => x"06",
          2835 => x"38",
          2836 => x"81",
          2837 => x"3f",
          2838 => x"e5",
          2839 => x"89",
          2840 => x"a5",
          2841 => x"80",
          2842 => x"83",
          2843 => x"57",
          2844 => x"51",
          2845 => x"83",
          2846 => x"70",
          2847 => x"84",
          2848 => x"3f",
          2849 => x"75",
          2850 => x"85",
          2851 => x"80",
          2852 => x"82",
          2853 => x"83",
          2854 => x"43",
          2855 => x"51",
          2856 => x"83",
          2857 => x"70",
          2858 => x"84",
          2859 => x"3f",
          2860 => x"60",
          2861 => x"ff",
          2862 => x"52",
          2863 => x"08",
          2864 => x"93",
          2865 => x"98",
          2866 => x"51",
          2867 => x"27",
          2868 => x"51",
          2869 => x"82",
          2870 => x"f6",
          2871 => x"98",
          2872 => x"0d",
          2873 => x"d5",
          2874 => x"e0",
          2875 => x"53",
          2876 => x"ff",
          2877 => x"0c",
          2878 => x"02",
          2879 => x"72",
          2880 => x"33",
          2881 => x"3d",
          2882 => x"05",
          2883 => x"56",
          2884 => x"e0",
          2885 => x"8c",
          2886 => x"2e",
          2887 => x"0c",
          2888 => x"71",
          2889 => x"0c",
          2890 => x"51",
          2891 => x"c0",
          2892 => x"71",
          2893 => x"92",
          2894 => x"70",
          2895 => x"94",
          2896 => x"51",
          2897 => x"0d",
          2898 => x"02",
          2899 => x"58",
          2900 => x"3f",
          2901 => x"54",
          2902 => x"75",
          2903 => x"87",
          2904 => x"84",
          2905 => x"85",
          2906 => x"7d",
          2907 => x"85",
          2908 => x"71",
          2909 => x"71",
          2910 => x"19",
          2911 => x"71",
          2912 => x"83",
          2913 => x"8a",
          2914 => x"71",
          2915 => x"52",
          2916 => x"80",
          2917 => x"c0",
          2918 => x"82",
          2919 => x"1a",
          2920 => x"19",
          2921 => x"79",
          2922 => x"80",
          2923 => x"26",
          2924 => x"06",
          2925 => x"52",
          2926 => x"8f",
          2927 => x"62",
          2928 => x"57",
          2929 => x"52",
          2930 => x"08",
          2931 => x"2e",
          2932 => x"74",
          2933 => x"87",
          2934 => x"84",
          2935 => x"0b",
          2936 => x"0c",
          2937 => x"70",
          2938 => x"54",
          2939 => x"81",
          2940 => x"58",
          2941 => x"52",
          2942 => x"98",
          2943 => x"c0",
          2944 => x"87",
          2945 => x"81",
          2946 => x"53",
          2947 => x"71",
          2948 => x"81",
          2949 => x"19",
          2950 => x"38",
          2951 => x"87",
          2952 => x"73",
          2953 => x"2e",
          2954 => x"82",
          2955 => x"fa",
          2956 => x"05",
          2957 => x"71",
          2958 => x"82",
          2959 => x"54",
          2960 => x"c0",
          2961 => x"2e",
          2962 => x"38",
          2963 => x"11",
          2964 => x"80",
          2965 => x"38",
          2966 => x"2a",
          2967 => x"80",
          2968 => x"08",
          2969 => x"8c",
          2970 => x"0c",
          2971 => x"08",
          2972 => x"38",
          2973 => x"80",
          2974 => x"77",
          2975 => x"75",
          2976 => x"3d",
          2977 => x"11",
          2978 => x"82",
          2979 => x"0d",
          2980 => x"33",
          2981 => x"88",
          2982 => x"07",
          2983 => x"e0",
          2984 => x"52",
          2985 => x"73",
          2986 => x"52",
          2987 => x"70",
          2988 => x"3d",
          2989 => x"52",
          2990 => x"34",
          2991 => x"81",
          2992 => x"70",
          2993 => x"88",
          2994 => x"0d",
          2995 => x"54",
          2996 => x"71",
          2997 => x"81",
          2998 => x"39",
          2999 => x"75",
          3000 => x"70",
          3001 => x"70",
          3002 => x"3d",
          3003 => x"74",
          3004 => x"81",
          3005 => x"16",
          3006 => x"86",
          3007 => x"82",
          3008 => x"fe",
          3009 => x"39",
          3010 => x"51",
          3011 => x"33",
          3012 => x"04",
          3013 => x"fb",
          3014 => x"81",
          3015 => x"56",
          3016 => x"08",
          3017 => x"83",
          3018 => x"3f",
          3019 => x"06",
          3020 => x"76",
          3021 => x"0c",
          3022 => x"7b",
          3023 => x"5a",
          3024 => x"54",
          3025 => x"53",
          3026 => x"3f",
          3027 => x"81",
          3028 => x"83",
          3029 => x"18",
          3030 => x"58",
          3031 => x"33",
          3032 => x"93",
          3033 => x"52",
          3034 => x"83",
          3035 => x"0c",
          3036 => x"78",
          3037 => x"17",
          3038 => x"fc",
          3039 => x"e0",
          3040 => x"53",
          3041 => x"f7",
          3042 => x"2e",
          3043 => x"b4",
          3044 => x"88",
          3045 => x"70",
          3046 => x"98",
          3047 => x"91",
          3048 => x"09",
          3049 => x"33",
          3050 => x"80",
          3051 => x"98",
          3052 => x"fc",
          3053 => x"b6",
          3054 => x"85",
          3055 => x"3f",
          3056 => x"9c",
          3057 => x"08",
          3058 => x"3f",
          3059 => x"51",
          3060 => x"05",
          3061 => x"75",
          3062 => x"3f",
          3063 => x"52",
          3064 => x"82",
          3065 => x"81",
          3066 => x"3d",
          3067 => x"1a",
          3068 => x"54",
          3069 => x"8a",
          3070 => x"08",
          3071 => x"0c",
          3072 => x"7a",
          3073 => x"77",
          3074 => x"08",
          3075 => x"54",
          3076 => x"72",
          3077 => x"8d",
          3078 => x"81",
          3079 => x"2a",
          3080 => x"05",
          3081 => x"82",
          3082 => x"83",
          3083 => x"17",
          3084 => x"55",
          3085 => x"3f",
          3086 => x"74",
          3087 => x"70",
          3088 => x"71",
          3089 => x"72",
          3090 => x"58",
          3091 => x"15",
          3092 => x"3f",
          3093 => x"76",
          3094 => x"05",
          3095 => x"08",
          3096 => x"76",
          3097 => x"73",
          3098 => x"08",
          3099 => x"06",
          3100 => x"3f",
          3101 => x"58",
          3102 => x"98",
          3103 => x"0d",
          3104 => x"59",
          3105 => x"9c",
          3106 => x"33",
          3107 => x"72",
          3108 => x"8d",
          3109 => x"81",
          3110 => x"2a",
          3111 => x"05",
          3112 => x"82",
          3113 => x"08",
          3114 => x"16",
          3115 => x"59",
          3116 => x"8f",
          3117 => x"74",
          3118 => x"72",
          3119 => x"74",
          3120 => x"75",
          3121 => x"08",
          3122 => x"38",
          3123 => x"78",
          3124 => x"77",
          3125 => x"71",
          3126 => x"34",
          3127 => x"17",
          3128 => x"3f",
          3129 => x"98",
          3130 => x"ff",
          3131 => x"76",
          3132 => x"be",
          3133 => x"05",
          3134 => x"e0",
          3135 => x"ab",
          3136 => x"2b",
          3137 => x"70",
          3138 => x"82",
          3139 => x"07",
          3140 => x"0b",
          3141 => x"0c",
          3142 => x"7a",
          3143 => x"59",
          3144 => x"17",
          3145 => x"aa",
          3146 => x"fd",
          3147 => x"82",
          3148 => x"39",
          3149 => x"80",
          3150 => x"80",
          3151 => x"84",
          3152 => x"e0",
          3153 => x"82",
          3154 => x"82",
          3155 => x"80",
          3156 => x"3f",
          3157 => x"16",
          3158 => x"55",
          3159 => x"15",
          3160 => x"07",
          3161 => x"76",
          3162 => x"73",
          3163 => x"04",
          3164 => x"59",
          3165 => x"08",
          3166 => x"17",
          3167 => x"ae",
          3168 => x"3f",
          3169 => x"27",
          3170 => x"55",
          3171 => x"d2",
          3172 => x"08",
          3173 => x"17",
          3174 => x"82",
          3175 => x"06",
          3176 => x"17",
          3177 => x"75",
          3178 => x"59",
          3179 => x"81",
          3180 => x"59",
          3181 => x"70",
          3182 => x"82",
          3183 => x"55",
          3184 => x"08",
          3185 => x"54",
          3186 => x"18",
          3187 => x"39",
          3188 => x"16",
          3189 => x"38",
          3190 => x"38",
          3191 => x"82",
          3192 => x"80",
          3193 => x"09",
          3194 => x"08",
          3195 => x"30",
          3196 => x"07",
          3197 => x"38",
          3198 => x"ae",
          3199 => x"53",
          3200 => x"82",
          3201 => x"30",
          3202 => x"25",
          3203 => x"38",
          3204 => x"79",
          3205 => x"e0",
          3206 => x"90",
          3207 => x"94",
          3208 => x"86",
          3209 => x"17",
          3210 => x"34",
          3211 => x"90",
          3212 => x"82",
          3213 => x"56",
          3214 => x"8c",
          3215 => x"70",
          3216 => x"98",
          3217 => x"08",
          3218 => x"f6",
          3219 => x"e0",
          3220 => x"80",
          3221 => x"57",
          3222 => x"81",
          3223 => x"78",
          3224 => x"53",
          3225 => x"ab",
          3226 => x"df",
          3227 => x"30",
          3228 => x"51",
          3229 => x"8a",
          3230 => x"7c",
          3231 => x"80",
          3232 => x"06",
          3233 => x"18",
          3234 => x"38",
          3235 => x"38",
          3236 => x"74",
          3237 => x"22",
          3238 => x"38",
          3239 => x"cd",
          3240 => x"54",
          3241 => x"52",
          3242 => x"98",
          3243 => x"2e",
          3244 => x"08",
          3245 => x"e0",
          3246 => x"bd",
          3247 => x"73",
          3248 => x"e0",
          3249 => x"18",
          3250 => x"72",
          3251 => x"58",
          3252 => x"18",
          3253 => x"05",
          3254 => x"e0",
          3255 => x"3d",
          3256 => x"a0",
          3257 => x"77",
          3258 => x"0c",
          3259 => x"80",
          3260 => x"06",
          3261 => x"98",
          3262 => x"92",
          3263 => x"56",
          3264 => x"80",
          3265 => x"77",
          3266 => x"38",
          3267 => x"82",
          3268 => x"0b",
          3269 => x"38",
          3270 => x"2e",
          3271 => x"e0",
          3272 => x"8a",
          3273 => x"80",
          3274 => x"51",
          3275 => x"53",
          3276 => x"2e",
          3277 => x"98",
          3278 => x"82",
          3279 => x"82",
          3280 => x"f3",
          3281 => x"72",
          3282 => x"f2",
          3283 => x"15",
          3284 => x"b8",
          3285 => x"82",
          3286 => x"f7",
          3287 => x"5b",
          3288 => x"3f",
          3289 => x"98",
          3290 => x"08",
          3291 => x"f0",
          3292 => x"82",
          3293 => x"e0",
          3294 => x"51",
          3295 => x"81",
          3296 => x"98",
          3297 => x"77",
          3298 => x"38",
          3299 => x"81",
          3300 => x"98",
          3301 => x"8e",
          3302 => x"e0",
          3303 => x"73",
          3304 => x"87",
          3305 => x"3d",
          3306 => x"11",
          3307 => x"98",
          3308 => x"33",
          3309 => x"81",
          3310 => x"92",
          3311 => x"73",
          3312 => x"85",
          3313 => x"79",
          3314 => x"12",
          3315 => x"70",
          3316 => x"81",
          3317 => x"94",
          3318 => x"0d",
          3319 => x"51",
          3320 => x"80",
          3321 => x"33",
          3322 => x"16",
          3323 => x"70",
          3324 => x"04",
          3325 => x"84",
          3326 => x"5d",
          3327 => x"80",
          3328 => x"ed",
          3329 => x"82",
          3330 => x"19",
          3331 => x"38",
          3332 => x"33",
          3333 => x"53",
          3334 => x"08",
          3335 => x"06",
          3336 => x"08",
          3337 => x"83",
          3338 => x"72",
          3339 => x"df",
          3340 => x"81",
          3341 => x"2e",
          3342 => x"39",
          3343 => x"ca",
          3344 => x"51",
          3345 => x"15",
          3346 => x"1c",
          3347 => x"73",
          3348 => x"38",
          3349 => x"09",
          3350 => x"08",
          3351 => x"82",
          3352 => x"53",
          3353 => x"81",
          3354 => x"54",
          3355 => x"17",
          3356 => x"82",
          3357 => x"56",
          3358 => x"fe",
          3359 => x"76",
          3360 => x"54",
          3361 => x"09",
          3362 => x"8c",
          3363 => x"86",
          3364 => x"72",
          3365 => x"26",
          3366 => x"73",
          3367 => x"51",
          3368 => x"5c",
          3369 => x"fc",
          3370 => x"ff",
          3371 => x"ff",
          3372 => x"52",
          3373 => x"98",
          3374 => x"38",
          3375 => x"39",
          3376 => x"e0",
          3377 => x"3d",
          3378 => x"52",
          3379 => x"98",
          3380 => x"a4",
          3381 => x"0b",
          3382 => x"7e",
          3383 => x"08",
          3384 => x"38",
          3385 => x"75",
          3386 => x"8b",
          3387 => x"06",
          3388 => x"81",
          3389 => x"2a",
          3390 => x"2e",
          3391 => x"8f",
          3392 => x"ab",
          3393 => x"06",
          3394 => x"75",
          3395 => x"73",
          3396 => x"76",
          3397 => x"ac",
          3398 => x"2e",
          3399 => x"17",
          3400 => x"06",
          3401 => x"18",
          3402 => x"98",
          3403 => x"81",
          3404 => x"8d",
          3405 => x"5c",
          3406 => x"05",
          3407 => x"08",
          3408 => x"2e",
          3409 => x"e6",
          3410 => x"82",
          3411 => x"22",
          3412 => x"e1",
          3413 => x"2e",
          3414 => x"5a",
          3415 => x"09",
          3416 => x"8c",
          3417 => x"70",
          3418 => x"57",
          3419 => x"2e",
          3420 => x"51",
          3421 => x"81",
          3422 => x"ff",
          3423 => x"38",
          3424 => x"98",
          3425 => x"2e",
          3426 => x"54",
          3427 => x"52",
          3428 => x"82",
          3429 => x"81",
          3430 => x"80",
          3431 => x"e0",
          3432 => x"80",
          3433 => x"98",
          3434 => x"0d",
          3435 => x"a0",
          3436 => x"85",
          3437 => x"22",
          3438 => x"38",
          3439 => x"51",
          3440 => x"1a",
          3441 => x"59",
          3442 => x"33",
          3443 => x"a8",
          3444 => x"81",
          3445 => x"8b",
          3446 => x"3f",
          3447 => x"56",
          3448 => x"55",
          3449 => x"83",
          3450 => x"8f",
          3451 => x"75",
          3452 => x"06",
          3453 => x"87",
          3454 => x"ff",
          3455 => x"c0",
          3456 => x"bf",
          3457 => x"06",
          3458 => x"14",
          3459 => x"18",
          3460 => x"e3",
          3461 => x"80",
          3462 => x"38",
          3463 => x"38",
          3464 => x"e0",
          3465 => x"8c",
          3466 => x"94",
          3467 => x"74",
          3468 => x"33",
          3469 => x"05",
          3470 => x"56",
          3471 => x"38",
          3472 => x"55",
          3473 => x"e3",
          3474 => x"e0",
          3475 => x"80",
          3476 => x"55",
          3477 => x"82",
          3478 => x"08",
          3479 => x"38",
          3480 => x"34",
          3481 => x"2a",
          3482 => x"59",
          3483 => x"8c",
          3484 => x"e0",
          3485 => x"51",
          3486 => x"57",
          3487 => x"ff",
          3488 => x"38",
          3489 => x"31",
          3490 => x"82",
          3491 => x"08",
          3492 => x"91",
          3493 => x"06",
          3494 => x"e3",
          3495 => x"82",
          3496 => x"1c",
          3497 => x"06",
          3498 => x"8f",
          3499 => x"08",
          3500 => x"52",
          3501 => x"8d",
          3502 => x"83",
          3503 => x"1b",
          3504 => x"73",
          3505 => x"05",
          3506 => x"83",
          3507 => x"77",
          3508 => x"2e",
          3509 => x"51",
          3510 => x"07",
          3511 => x"1d",
          3512 => x"3f",
          3513 => x"98",
          3514 => x"78",
          3515 => x"7b",
          3516 => x"08",
          3517 => x"a0",
          3518 => x"1a",
          3519 => x"a0",
          3520 => x"91",
          3521 => x"98",
          3522 => x"81",
          3523 => x"82",
          3524 => x"fa",
          3525 => x"08",
          3526 => x"72",
          3527 => x"51",
          3528 => x"54",
          3529 => x"98",
          3530 => x"3f",
          3531 => x"98",
          3532 => x"e5",
          3533 => x"90",
          3534 => x"e0",
          3535 => x"3f",
          3536 => x"98",
          3537 => x"2e",
          3538 => x"73",
          3539 => x"04",
          3540 => x"5f",
          3541 => x"98",
          3542 => x"ac",
          3543 => x"80",
          3544 => x"22",
          3545 => x"2e",
          3546 => x"22",
          3547 => x"38",
          3548 => x"ff",
          3549 => x"86",
          3550 => x"18",
          3551 => x"5b",
          3552 => x"75",
          3553 => x"e0",
          3554 => x"81",
          3555 => x"27",
          3556 => x"7a",
          3557 => x"9f",
          3558 => x"07",
          3559 => x"54",
          3560 => x"57",
          3561 => x"74",
          3562 => x"79",
          3563 => x"72",
          3564 => x"25",
          3565 => x"77",
          3566 => x"14",
          3567 => x"57",
          3568 => x"1b",
          3569 => x"38",
          3570 => x"38",
          3571 => x"30",
          3572 => x"54",
          3573 => x"2e",
          3574 => x"58",
          3575 => x"81",
          3576 => x"79",
          3577 => x"05",
          3578 => x"18",
          3579 => x"8b",
          3580 => x"57",
          3581 => x"33",
          3582 => x"d3",
          3583 => x"73",
          3584 => x"99",
          3585 => x"11",
          3586 => x"38",
          3587 => x"83",
          3588 => x"80",
          3589 => x"ff",
          3590 => x"81",
          3591 => x"81",
          3592 => x"72",
          3593 => x"53",
          3594 => x"08",
          3595 => x"38",
          3596 => x"53",
          3597 => x"1c",
          3598 => x"3f",
          3599 => x"13",
          3600 => x"08",
          3601 => x"fa",
          3602 => x"23",
          3603 => x"62",
          3604 => x"33",
          3605 => x"38",
          3606 => x"38",
          3607 => x"05",
          3608 => x"15",
          3609 => x"56",
          3610 => x"38",
          3611 => x"30",
          3612 => x"54",
          3613 => x"63",
          3614 => x"96",
          3615 => x"80",
          3616 => x"e0",
          3617 => x"41",
          3618 => x"80",
          3619 => x"8f",
          3620 => x"82",
          3621 => x"e0",
          3622 => x"1a",
          3623 => x"55",
          3624 => x"e0",
          3625 => x"af",
          3626 => x"80",
          3627 => x"b4",
          3628 => x"75",
          3629 => x"82",
          3630 => x"e0",
          3631 => x"fe",
          3632 => x"54",
          3633 => x"89",
          3634 => x"33",
          3635 => x"81",
          3636 => x"dc",
          3637 => x"07",
          3638 => x"44",
          3639 => x"81",
          3640 => x"22",
          3641 => x"d2",
          3642 => x"80",
          3643 => x"ae",
          3644 => x"79",
          3645 => x"06",
          3646 => x"74",
          3647 => x"ae",
          3648 => x"54",
          3649 => x"81",
          3650 => x"76",
          3651 => x"84",
          3652 => x"78",
          3653 => x"fe",
          3654 => x"70",
          3655 => x"54",
          3656 => x"38",
          3657 => x"19",
          3658 => x"78",
          3659 => x"76",
          3660 => x"7a",
          3661 => x"56",
          3662 => x"93",
          3663 => x"22",
          3664 => x"38",
          3665 => x"06",
          3666 => x"85",
          3667 => x"2e",
          3668 => x"22",
          3669 => x"78",
          3670 => x"59",
          3671 => x"70",
          3672 => x"81",
          3673 => x"a0",
          3674 => x"59",
          3675 => x"22",
          3676 => x"2e",
          3677 => x"38",
          3678 => x"25",
          3679 => x"38",
          3680 => x"07",
          3681 => x"7e",
          3682 => x"79",
          3683 => x"25",
          3684 => x"73",
          3685 => x"fe",
          3686 => x"76",
          3687 => x"be",
          3688 => x"82",
          3689 => x"8b",
          3690 => x"76",
          3691 => x"51",
          3692 => x"08",
          3693 => x"70",
          3694 => x"2e",
          3695 => x"d2",
          3696 => x"76",
          3697 => x"78",
          3698 => x"59",
          3699 => x"05",
          3700 => x"34",
          3701 => x"80",
          3702 => x"d0",
          3703 => x"08",
          3704 => x"83",
          3705 => x"16",
          3706 => x"82",
          3707 => x"99",
          3708 => x"17",
          3709 => x"5c",
          3710 => x"34",
          3711 => x"1e",
          3712 => x"81",
          3713 => x"34",
          3714 => x"38",
          3715 => x"7b",
          3716 => x"38",
          3717 => x"09",
          3718 => x"57",
          3719 => x"54",
          3720 => x"73",
          3721 => x"57",
          3722 => x"54",
          3723 => x"07",
          3724 => x"ea",
          3725 => x"1f",
          3726 => x"80",
          3727 => x"84",
          3728 => x"74",
          3729 => x"2a",
          3730 => x"38",
          3731 => x"f8",
          3732 => x"34",
          3733 => x"06",
          3734 => x"39",
          3735 => x"54",
          3736 => x"84",
          3737 => x"73",
          3738 => x"83",
          3739 => x"7f",
          3740 => x"08",
          3741 => x"82",
          3742 => x"f6",
          3743 => x"70",
          3744 => x"73",
          3745 => x"81",
          3746 => x"52",
          3747 => x"38",
          3748 => x"a5",
          3749 => x"ff",
          3750 => x"91",
          3751 => x"d0",
          3752 => x"f7",
          3753 => x"55",
          3754 => x"81",
          3755 => x"56",
          3756 => x"70",
          3757 => x"81",
          3758 => x"51",
          3759 => x"70",
          3760 => x"70",
          3761 => x"09",
          3762 => x"38",
          3763 => x"70",
          3764 => x"07",
          3765 => x"8f",
          3766 => x"83",
          3767 => x"74",
          3768 => x"0c",
          3769 => x"f4",
          3770 => x"8c",
          3771 => x"56",
          3772 => x"b4",
          3773 => x"f4",
          3774 => x"81",
          3775 => x"8a",
          3776 => x"ff",
          3777 => x"d5",
          3778 => x"80",
          3779 => x"81",
          3780 => x"81",
          3781 => x"70",
          3782 => x"73",
          3783 => x"81",
          3784 => x"d8",
          3785 => x"3f",
          3786 => x"98",
          3787 => x"82",
          3788 => x"ce",
          3789 => x"82",
          3790 => x"82",
          3791 => x"3d",
          3792 => x"84",
          3793 => x"80",
          3794 => x"82",
          3795 => x"0b",
          3796 => x"38",
          3797 => x"f7",
          3798 => x"56",
          3799 => x"75",
          3800 => x"54",
          3801 => x"14",
          3802 => x"98",
          3803 => x"54",
          3804 => x"87",
          3805 => x"06",
          3806 => x"38",
          3807 => x"18",
          3808 => x"15",
          3809 => x"c6",
          3810 => x"ff",
          3811 => x"56",
          3812 => x"8f",
          3813 => x"51",
          3814 => x"80",
          3815 => x"3f",
          3816 => x"57",
          3817 => x"26",
          3818 => x"33",
          3819 => x"8c",
          3820 => x"fa",
          3821 => x"2e",
          3822 => x"a9",
          3823 => x"79",
          3824 => x"90",
          3825 => x"38",
          3826 => x"70",
          3827 => x"95",
          3828 => x"5a",
          3829 => x"5b",
          3830 => x"7a",
          3831 => x"e0",
          3832 => x"0b",
          3833 => x"72",
          3834 => x"81",
          3835 => x"80",
          3836 => x"56",
          3837 => x"56",
          3838 => x"56",
          3839 => x"c3",
          3840 => x"98",
          3841 => x"84",
          3842 => x"38",
          3843 => x"82",
          3844 => x"58",
          3845 => x"c9",
          3846 => x"77",
          3847 => x"82",
          3848 => x"11",
          3849 => x"8d",
          3850 => x"74",
          3851 => x"c5",
          3852 => x"15",
          3853 => x"13",
          3854 => x"38",
          3855 => x"14",
          3856 => x"08",
          3857 => x"23",
          3858 => x"83",
          3859 => x"ea",
          3860 => x"ff",
          3861 => x"14",
          3862 => x"08",
          3863 => x"3f",
          3864 => x"06",
          3865 => x"9e",
          3866 => x"84",
          3867 => x"83",
          3868 => x"79",
          3869 => x"e0",
          3870 => x"80",
          3871 => x"08",
          3872 => x"38",
          3873 => x"83",
          3874 => x"85",
          3875 => x"76",
          3876 => x"70",
          3877 => x"73",
          3878 => x"b0",
          3879 => x"09",
          3880 => x"51",
          3881 => x"83",
          3882 => x"82",
          3883 => x"e4",
          3884 => x"98",
          3885 => x"53",
          3886 => x"81",
          3887 => x"74",
          3888 => x"74",
          3889 => x"06",
          3890 => x"2a",
          3891 => x"26",
          3892 => x"0c",
          3893 => x"0b",
          3894 => x"81",
          3895 => x"51",
          3896 => x"83",
          3897 => x"09",
          3898 => x"52",
          3899 => x"98",
          3900 => x"08",
          3901 => x"c6",
          3902 => x"ff",
          3903 => x"2e",
          3904 => x"14",
          3905 => x"08",
          3906 => x"81",
          3907 => x"c6",
          3908 => x"8a",
          3909 => x"9d",
          3910 => x"3f",
          3911 => x"84",
          3912 => x"e0",
          3913 => x"34",
          3914 => x"72",
          3915 => x"23",
          3916 => x"80",
          3917 => x"82",
          3918 => x"fb",
          3919 => x"80",
          3920 => x"80",
          3921 => x"80",
          3922 => x"15",
          3923 => x"81",
          3924 => x"ff",
          3925 => x"81",
          3926 => x"08",
          3927 => x"73",
          3928 => x"0c",
          3929 => x"02",
          3930 => x"fc",
          3931 => x"54",
          3932 => x"bc",
          3933 => x"82",
          3934 => x"73",
          3935 => x"78",
          3936 => x"74",
          3937 => x"80",
          3938 => x"70",
          3939 => x"82",
          3940 => x"98",
          3941 => x"0d",
          3942 => x"33",
          3943 => x"84",
          3944 => x"99",
          3945 => x"05",
          3946 => x"98",
          3947 => x"a4",
          3948 => x"70",
          3949 => x"98",
          3950 => x"38",
          3951 => x"2b",
          3952 => x"86",
          3953 => x"2e",
          3954 => x"38",
          3955 => x"38",
          3956 => x"98",
          3957 => x"33",
          3958 => x"77",
          3959 => x"73",
          3960 => x"bc",
          3961 => x"b4",
          3962 => x"51",
          3963 => x"62",
          3964 => x"e0",
          3965 => x"52",
          3966 => x"62",
          3967 => x"53",
          3968 => x"80",
          3969 => x"3f",
          3970 => x"75",
          3971 => x"11",
          3972 => x"98",
          3973 => x"82",
          3974 => x"08",
          3975 => x"c4",
          3976 => x"2a",
          3977 => x"80",
          3978 => x"39",
          3979 => x"54",
          3980 => x"06",
          3981 => x"55",
          3982 => x"c4",
          3983 => x"ff",
          3984 => x"e0",
          3985 => x"2a",
          3986 => x"2e",
          3987 => x"7a",
          3988 => x"a4",
          3989 => x"d5",
          3990 => x"e0",
          3991 => x"05",
          3992 => x"98",
          3993 => x"0c",
          3994 => x"84",
          3995 => x"0b",
          3996 => x"0c",
          3997 => x"2a",
          3998 => x"2e",
          3999 => x"80",
          4000 => x"08",
          4001 => x"89",
          4002 => x"76",
          4003 => x"e0",
          4004 => x"81",
          4005 => x"98",
          4006 => x"38",
          4007 => x"30",
          4008 => x"77",
          4009 => x"06",
          4010 => x"1a",
          4011 => x"06",
          4012 => x"52",
          4013 => x"98",
          4014 => x"75",
          4015 => x"9c",
          4016 => x"74",
          4017 => x"3d",
          4018 => x"65",
          4019 => x"0c",
          4020 => x"f9",
          4021 => x"82",
          4022 => x"33",
          4023 => x"56",
          4024 => x"06",
          4025 => x"b9",
          4026 => x"34",
          4027 => x"91",
          4028 => x"8c",
          4029 => x"74",
          4030 => x"80",
          4031 => x"70",
          4032 => x"b4",
          4033 => x"77",
          4034 => x"38",
          4035 => x"8f",
          4036 => x"c3",
          4037 => x"81",
          4038 => x"2e",
          4039 => x"98",
          4040 => x"3f",
          4041 => x"83",
          4042 => x"89",
          4043 => x"d8",
          4044 => x"58",
          4045 => x"75",
          4046 => x"7c",
          4047 => x"91",
          4048 => x"38",
          4049 => x"80",
          4050 => x"31",
          4051 => x"80",
          4052 => x"77",
          4053 => x"bd",
          4054 => x"39",
          4055 => x"83",
          4056 => x"55",
          4057 => x"9c",
          4058 => x"3f",
          4059 => x"75",
          4060 => x"1f",
          4061 => x"a9",
          4062 => x"7f",
          4063 => x"94",
          4064 => x"80",
          4065 => x"3d",
          4066 => x"65",
          4067 => x"0c",
          4068 => x"f6",
          4069 => x"82",
          4070 => x"33",
          4071 => x"56",
          4072 => x"81",
          4073 => x"87",
          4074 => x"95",
          4075 => x"56",
          4076 => x"34",
          4077 => x"08",
          4078 => x"84",
          4079 => x"82",
          4080 => x"ff",
          4081 => x"7e",
          4082 => x"2a",
          4083 => x"8c",
          4084 => x"38",
          4085 => x"52",
          4086 => x"98",
          4087 => x"2e",
          4088 => x"91",
          4089 => x"74",
          4090 => x"38",
          4091 => x"15",
          4092 => x"06",
          4093 => x"3f",
          4094 => x"98",
          4095 => x"da",
          4096 => x"fe",
          4097 => x"7c",
          4098 => x"80",
          4099 => x"22",
          4100 => x"38",
          4101 => x"53",
          4102 => x"b6",
          4103 => x"a3",
          4104 => x"56",
          4105 => x"80",
          4106 => x"2b",
          4107 => x"ba",
          4108 => x"16",
          4109 => x"39",
          4110 => x"94",
          4111 => x"82",
          4112 => x"77",
          4113 => x"0c",
          4114 => x"80",
          4115 => x"83",
          4116 => x"7e",
          4117 => x"98",
          4118 => x"52",
          4119 => x"b8",
          4120 => x"55",
          4121 => x"31",
          4122 => x"94",
          4123 => x"8c",
          4124 => x"76",
          4125 => x"19",
          4126 => x"80",
          4127 => x"80",
          4128 => x"3d",
          4129 => x"3d",
          4130 => x"df",
          4131 => x"e0",
          4132 => x"33",
          4133 => x"55",
          4134 => x"a0",
          4135 => x"a4",
          4136 => x"e0",
          4137 => x"08",
          4138 => x"73",
          4139 => x"74",
          4140 => x"8c",
          4141 => x"b7",
          4142 => x"96",
          4143 => x"52",
          4144 => x"78",
          4145 => x"51",
          4146 => x"08",
          4147 => x"57",
          4148 => x"98",
          4149 => x"0d",
          4150 => x"82",
          4151 => x"08",
          4152 => x"73",
          4153 => x"08",
          4154 => x"82",
          4155 => x"e0",
          4156 => x"3d",
          4157 => x"8b",
          4158 => x"24",
          4159 => x"f7",
          4160 => x"98",
          4161 => x"0d",
          4162 => x"95",
          4163 => x"98",
          4164 => x"e0",
          4165 => x"d0",
          4166 => x"98",
          4167 => x"38",
          4168 => x"2b",
          4169 => x"76",
          4170 => x"02",
          4171 => x"81",
          4172 => x"9e",
          4173 => x"c9",
          4174 => x"15",
          4175 => x"84",
          4176 => x"55",
          4177 => x"0d",
          4178 => x"3d",
          4179 => x"80",
          4180 => x"fd",
          4181 => x"e7",
          4182 => x"82",
          4183 => x"80",
          4184 => x"08",
          4185 => x"d5",
          4186 => x"83",
          4187 => x"52",
          4188 => x"08",
          4189 => x"38",
          4190 => x"ff",
          4191 => x"57",
          4192 => x"80",
          4193 => x"c2",
          4194 => x"3d",
          4195 => x"3f",
          4196 => x"98",
          4197 => x"51",
          4198 => x"57",
          4199 => x"da",
          4200 => x"3f",
          4201 => x"38",
          4202 => x"82",
          4203 => x"08",
          4204 => x"09",
          4205 => x"ee",
          4206 => x"3d",
          4207 => x"a0",
          4208 => x"11",
          4209 => x"2e",
          4210 => x"81",
          4211 => x"56",
          4212 => x"78",
          4213 => x"9c",
          4214 => x"18",
          4215 => x"ff",
          4216 => x"74",
          4217 => x"e1",
          4218 => x"34",
          4219 => x"81",
          4220 => x"3d",
          4221 => x"80",
          4222 => x"29",
          4223 => x"33",
          4224 => x"2e",
          4225 => x"33",
          4226 => x"16",
          4227 => x"55",
          4228 => x"54",
          4229 => x"34",
          4230 => x"70",
          4231 => x"09",
          4232 => x"39",
          4233 => x"59",
          4234 => x"5c",
          4235 => x"7a",
          4236 => x"df",
          4237 => x"7d",
          4238 => x"57",
          4239 => x"08",
          4240 => x"38",
          4241 => x"38",
          4242 => x"92",
          4243 => x"70",
          4244 => x"38",
          4245 => x"70",
          4246 => x"82",
          4247 => x"89",
          4248 => x"b7",
          4249 => x"bc",
          4250 => x"15",
          4251 => x"bb",
          4252 => x"26",
          4253 => x"70",
          4254 => x"18",
          4255 => x"88",
          4256 => x"52",
          4257 => x"e0",
          4258 => x"81",
          4259 => x"08",
          4260 => x"98",
          4261 => x"0c",
          4262 => x"76",
          4263 => x"94",
          4264 => x"16",
          4265 => x"51",
          4266 => x"38",
          4267 => x"3f",
          4268 => x"98",
          4269 => x"56",
          4270 => x"b5",
          4271 => x"73",
          4272 => x"b0",
          4273 => x"27",
          4274 => x"9e",
          4275 => x"0c",
          4276 => x"2e",
          4277 => x"b4",
          4278 => x"38",
          4279 => x"80",
          4280 => x"81",
          4281 => x"e0",
          4282 => x"54",
          4283 => x"73",
          4284 => x"c0",
          4285 => x"83",
          4286 => x"38",
          4287 => x"77",
          4288 => x"e0",
          4289 => x"3d",
          4290 => x"2e",
          4291 => x"fc",
          4292 => x"e0",
          4293 => x"82",
          4294 => x"76",
          4295 => x"3f",
          4296 => x"98",
          4297 => x"70",
          4298 => x"a2",
          4299 => x"70",
          4300 => x"2e",
          4301 => x"51",
          4302 => x"88",
          4303 => x"84",
          4304 => x"bc",
          4305 => x"74",
          4306 => x"85",
          4307 => x"38",
          4308 => x"e0",
          4309 => x"3d",
          4310 => x"70",
          4311 => x"98",
          4312 => x"73",
          4313 => x"0d",
          4314 => x"71",
          4315 => x"e0",
          4316 => x"80",
          4317 => x"98",
          4318 => x"3f",
          4319 => x"39",
          4320 => x"c1",
          4321 => x"82",
          4322 => x"06",
          4323 => x"e0",
          4324 => x"51",
          4325 => x"ff",
          4326 => x"84",
          4327 => x"2c",
          4328 => x"51",
          4329 => x"87",
          4330 => x"57",
          4331 => x"3d",
          4332 => x"98",
          4333 => x"38",
          4334 => x"82",
          4335 => x"08",
          4336 => x"70",
          4337 => x"85",
          4338 => x"2e",
          4339 => x"80",
          4340 => x"3d",
          4341 => x"55",
          4342 => x"52",
          4343 => x"e0",
          4344 => x"82",
          4345 => x"9c",
          4346 => x"59",
          4347 => x"38",
          4348 => x"5b",
          4349 => x"39",
          4350 => x"59",
          4351 => x"c0",
          4352 => x"92",
          4353 => x"3f",
          4354 => x"38",
          4355 => x"38",
          4356 => x"e0",
          4357 => x"81",
          4358 => x"14",
          4359 => x"39",
          4360 => x"57",
          4361 => x"18",
          4362 => x"82",
          4363 => x"08",
          4364 => x"12",
          4365 => x"82",
          4366 => x"14",
          4367 => x"98",
          4368 => x"70",
          4369 => x"51",
          4370 => x"a9",
          4371 => x"0a",
          4372 => x"84",
          4373 => x"ff",
          4374 => x"38",
          4375 => x"0c",
          4376 => x"74",
          4377 => x"0c",
          4378 => x"79",
          4379 => x"57",
          4380 => x"56",
          4381 => x"91",
          4382 => x"90",
          4383 => x"06",
          4384 => x"2e",
          4385 => x"73",
          4386 => x"73",
          4387 => x"88",
          4388 => x"8c",
          4389 => x"19",
          4390 => x"08",
          4391 => x"82",
          4392 => x"06",
          4393 => x"08",
          4394 => x"82",
          4395 => x"54",
          4396 => x"27",
          4397 => x"e0",
          4398 => x"bc",
          4399 => x"17",
          4400 => x"80",
          4401 => x"75",
          4402 => x"34",
          4403 => x"89",
          4404 => x"53",
          4405 => x"3d",
          4406 => x"08",
          4407 => x"38",
          4408 => x"3d",
          4409 => x"e0",
          4410 => x"81",
          4411 => x"70",
          4412 => x"56",
          4413 => x"98",
          4414 => x"38",
          4415 => x"06",
          4416 => x"38",
          4417 => x"3f",
          4418 => x"70",
          4419 => x"2e",
          4420 => x"98",
          4421 => x"38",
          4422 => x"76",
          4423 => x"b5",
          4424 => x"82",
          4425 => x"e0",
          4426 => x"90",
          4427 => x"e0",
          4428 => x"d0",
          4429 => x"88",
          4430 => x"38",
          4431 => x"98",
          4432 => x"82",
          4433 => x"55",
          4434 => x"80",
          4435 => x"77",
          4436 => x"98",
          4437 => x"ff",
          4438 => x"55",
          4439 => x"0d",
          4440 => x"3d",
          4441 => x"d7",
          4442 => x"82",
          4443 => x"5e",
          4444 => x"cb",
          4445 => x"82",
          4446 => x"82",
          4447 => x"2e",
          4448 => x"80",
          4449 => x"06",
          4450 => x"38",
          4451 => x"52",
          4452 => x"98",
          4453 => x"08",
          4454 => x"08",
          4455 => x"82",
          4456 => x"09",
          4457 => x"ba",
          4458 => x"98",
          4459 => x"3f",
          4460 => x"98",
          4461 => x"52",
          4462 => x"78",
          4463 => x"54",
          4464 => x"88",
          4465 => x"ff",
          4466 => x"11",
          4467 => x"53",
          4468 => x"51",
          4469 => x"0b",
          4470 => x"80",
          4471 => x"3f",
          4472 => x"77",
          4473 => x"98",
          4474 => x"38",
          4475 => x"05",
          4476 => x"64",
          4477 => x"64",
          4478 => x"54",
          4479 => x"ff",
          4480 => x"54",
          4481 => x"51",
          4482 => x"98",
          4483 => x"0d",
          4484 => x"3f",
          4485 => x"52",
          4486 => x"e0",
          4487 => x"82",
          4488 => x"52",
          4489 => x"3f",
          4490 => x"98",
          4491 => x"05",
          4492 => x"73",
          4493 => x"08",
          4494 => x"ff",
          4495 => x"92",
          4496 => x"3f",
          4497 => x"8c",
          4498 => x"e0",
          4499 => x"08",
          4500 => x"a3",
          4501 => x"81",
          4502 => x"2e",
          4503 => x"51",
          4504 => x"08",
          4505 => x"38",
          4506 => x"8d",
          4507 => x"b9",
          4508 => x"34",
          4509 => x"81",
          4510 => x"74",
          4511 => x"78",
          4512 => x"16",
          4513 => x"51",
          4514 => x"38",
          4515 => x"52",
          4516 => x"e0",
          4517 => x"aa",
          4518 => x"80",
          4519 => x"08",
          4520 => x"82",
          4521 => x"58",
          4522 => x"c1",
          4523 => x"2e",
          4524 => x"75",
          4525 => x"78",
          4526 => x"39",
          4527 => x"51",
          4528 => x"55",
          4529 => x"51",
          4530 => x"08",
          4531 => x"3d",
          4532 => x"df",
          4533 => x"05",
          4534 => x"cc",
          4535 => x"3f",
          4536 => x"98",
          4537 => x"52",
          4538 => x"3f",
          4539 => x"98",
          4540 => x"33",
          4541 => x"aa",
          4542 => x"8b",
          4543 => x"07",
          4544 => x"34",
          4545 => x"78",
          4546 => x"98",
          4547 => x"96",
          4548 => x"56",
          4549 => x"95",
          4550 => x"98",
          4551 => x"cb",
          4552 => x"d0",
          4553 => x"98",
          4554 => x"38",
          4555 => x"06",
          4556 => x"16",
          4557 => x"07",
          4558 => x"f2",
          4559 => x"34",
          4560 => x"e0",
          4561 => x"0c",
          4562 => x"6a",
          4563 => x"cc",
          4564 => x"3f",
          4565 => x"08",
          4566 => x"80",
          4567 => x"81",
          4568 => x"55",
          4569 => x"5d",
          4570 => x"52",
          4571 => x"98",
          4572 => x"d2",
          4573 => x"f8",
          4574 => x"e0",
          4575 => x"08",
          4576 => x"56",
          4577 => x"59",
          4578 => x"56",
          4579 => x"75",
          4580 => x"2e",
          4581 => x"33",
          4582 => x"38",
          4583 => x"06",
          4584 => x"76",
          4585 => x"54",
          4586 => x"80",
          4587 => x"53",
          4588 => x"98",
          4589 => x"38",
          4590 => x"56",
          4591 => x"56",
          4592 => x"75",
          4593 => x"3f",
          4594 => x"82",
          4595 => x"e6",
          4596 => x"b4",
          4597 => x"3f",
          4598 => x"08",
          4599 => x"dd",
          4600 => x"70",
          4601 => x"6d",
          4602 => x"27",
          4603 => x"51",
          4604 => x"08",
          4605 => x"82",
          4606 => x"83",
          4607 => x"95",
          4608 => x"ff",
          4609 => x"38",
          4610 => x"9b",
          4611 => x"38",
          4612 => x"89",
          4613 => x"27",
          4614 => x"81",
          4615 => x"2a",
          4616 => x"34",
          4617 => x"05",
          4618 => x"51",
          4619 => x"38",
          4620 => x"81",
          4621 => x"2e",
          4622 => x"15",
          4623 => x"09",
          4624 => x"75",
          4625 => x"52",
          4626 => x"db",
          4627 => x"e0",
          4628 => x"74",
          4629 => x"98",
          4630 => x"38",
          4631 => x"74",
          4632 => x"08",
          4633 => x"38",
          4634 => x"38",
          4635 => x"3f",
          4636 => x"98",
          4637 => x"98",
          4638 => x"3f",
          4639 => x"8b",
          4640 => x"91",
          4641 => x"34",
          4642 => x"e0",
          4643 => x"e0",
          4644 => x"3d",
          4645 => x"cb",
          4646 => x"72",
          4647 => x"82",
          4648 => x"08",
          4649 => x"77",
          4650 => x"38",
          4651 => x"90",
          4652 => x"06",
          4653 => x"54",
          4654 => x"39",
          4655 => x"11",
          4656 => x"54",
          4657 => x"ff",
          4658 => x"07",
          4659 => x"90",
          4660 => x"55",
          4661 => x"08",
          4662 => x"77",
          4663 => x"51",
          4664 => x"55",
          4665 => x"38",
          4666 => x"2e",
          4667 => x"ff",
          4668 => x"08",
          4669 => x"2e",
          4670 => x"74",
          4671 => x"81",
          4672 => x"ff",
          4673 => x"7b",
          4674 => x"81",
          4675 => x"06",
          4676 => x"52",
          4677 => x"e0",
          4678 => x"80",
          4679 => x"56",
          4680 => x"ff",
          4681 => x"55",
          4682 => x"1b",
          4683 => x"33",
          4684 => x"34",
          4685 => x"08",
          4686 => x"75",
          4687 => x"33",
          4688 => x"77",
          4689 => x"3d",
          4690 => x"02",
          4691 => x"3d",
          4692 => x"8b",
          4693 => x"24",
          4694 => x"84",
          4695 => x"51",
          4696 => x"75",
          4697 => x"98",
          4698 => x"82",
          4699 => x"81",
          4700 => x"82",
          4701 => x"81",
          4702 => x"da",
          4703 => x"51",
          4704 => x"9a",
          4705 => x"51",
          4706 => x"08",
          4707 => x"92",
          4708 => x"38",
          4709 => x"2e",
          4710 => x"87",
          4711 => x"78",
          4712 => x"19",
          4713 => x"38",
          4714 => x"2a",
          4715 => x"59",
          4716 => x"56",
          4717 => x"51",
          4718 => x"64",
          4719 => x"74",
          4720 => x"89",
          4721 => x"8b",
          4722 => x"92",
          4723 => x"ff",
          4724 => x"d4",
          4725 => x"38",
          4726 => x"33",
          4727 => x"38",
          4728 => x"3f",
          4729 => x"52",
          4730 => x"98",
          4731 => x"05",
          4732 => x"f7",
          4733 => x"8a",
          4734 => x"06",
          4735 => x"74",
          4736 => x"56",
          4737 => x"7f",
          4738 => x"27",
          4739 => x"80",
          4740 => x"70",
          4741 => x"95",
          4742 => x"2e",
          4743 => x"74",
          4744 => x"06",
          4745 => x"2e",
          4746 => x"2e",
          4747 => x"ae",
          4748 => x"82",
          4749 => x"2e",
          4750 => x"82",
          4751 => x"70",
          4752 => x"86",
          4753 => x"52",
          4754 => x"e0",
          4755 => x"70",
          4756 => x"0b",
          4757 => x"05",
          4758 => x"27",
          4759 => x"ae",
          4760 => x"82",
          4761 => x"2e",
          4762 => x"82",
          4763 => x"70",
          4764 => x"86",
          4765 => x"52",
          4766 => x"e0",
          4767 => x"e0",
          4768 => x"81",
          4769 => x"e0",
          4770 => x"83",
          4771 => x"89",
          4772 => x"1f",
          4773 => x"ff",
          4774 => x"31",
          4775 => x"83",
          4776 => x"1c",
          4777 => x"1d",
          4778 => x"31",
          4779 => x"87",
          4780 => x"7a",
          4781 => x"9a",
          4782 => x"7d",
          4783 => x"82",
          4784 => x"80",
          4785 => x"81",
          4786 => x"ad",
          4787 => x"80",
          4788 => x"e0",
          4789 => x"38",
          4790 => x"86",
          4791 => x"81",
          4792 => x"83",
          4793 => x"08",
          4794 => x"ed",
          4795 => x"27",
          4796 => x"55",
          4797 => x"38",
          4798 => x"38",
          4799 => x"86",
          4800 => x"7a",
          4801 => x"82",
          4802 => x"81",
          4803 => x"ff",
          4804 => x"7b",
          4805 => x"51",
          4806 => x"1c",
          4807 => x"96",
          4808 => x"91",
          4809 => x"55",
          4810 => x"74",
          4811 => x"51",
          4812 => x"52",
          4813 => x"f8",
          4814 => x"1b",
          4815 => x"52",
          4816 => x"7e",
          4817 => x"3f",
          4818 => x"cb",
          4819 => x"c3",
          4820 => x"52",
          4821 => x"82",
          4822 => x"3f",
          4823 => x"8c",
          4824 => x"8d",
          4825 => x"1c",
          4826 => x"93",
          4827 => x"1b",
          4828 => x"52",
          4829 => x"7c",
          4830 => x"51",
          4831 => x"a4",
          4832 => x"93",
          4833 => x"51",
          4834 => x"52",
          4835 => x"8c",
          4836 => x"52",
          4837 => x"56",
          4838 => x"7d",
          4839 => x"38",
          4840 => x"7f",
          4841 => x"53",
          4842 => x"3f",
          4843 => x"51",
          4844 => x"e4",
          4845 => x"8b",
          4846 => x"1b",
          4847 => x"83",
          4848 => x"82",
          4849 => x"bc",
          4850 => x"52",
          4851 => x"54",
          4852 => x"ff",
          4853 => x"7a",
          4854 => x"80",
          4855 => x"9a",
          4856 => x"a2",
          4857 => x"8b",
          4858 => x"51",
          4859 => x"7d",
          4860 => x"52",
          4861 => x"55",
          4862 => x"74",
          4863 => x"7f",
          4864 => x"98",
          4865 => x"82",
          4866 => x"8b",
          4867 => x"56",
          4868 => x"77",
          4869 => x"7d",
          4870 => x"57",
          4871 => x"76",
          4872 => x"ff",
          4873 => x"81",
          4874 => x"56",
          4875 => x"83",
          4876 => x"ff",
          4877 => x"82",
          4878 => x"2e",
          4879 => x"52",
          4880 => x"56",
          4881 => x"64",
          4882 => x"16",
          4883 => x"53",
          4884 => x"3f",
          4885 => x"06",
          4886 => x"53",
          4887 => x"3f",
          4888 => x"89",
          4889 => x"75",
          4890 => x"0b",
          4891 => x"76",
          4892 => x"fd",
          4893 => x"3f",
          4894 => x"98",
          4895 => x"86",
          4896 => x"16",
          4897 => x"ff",
          4898 => x"1b",
          4899 => x"77",
          4900 => x"d3",
          4901 => x"a2",
          4902 => x"ff",
          4903 => x"98",
          4904 => x"8a",
          4905 => x"98",
          4906 => x"9a",
          4907 => x"60",
          4908 => x"5a",
          4909 => x"8d",
          4910 => x"fc",
          4911 => x"7a",
          4912 => x"8c",
          4913 => x"38",
          4914 => x"81",
          4915 => x"06",
          4916 => x"76",
          4917 => x"98",
          4918 => x"0d",
          4919 => x"59",
          4920 => x"87",
          4921 => x"84",
          4922 => x"38",
          4923 => x"56",
          4924 => x"bb",
          4925 => x"05",
          4926 => x"08",
          4927 => x"70",
          4928 => x"30",
          4929 => x"0c",
          4930 => x"0d",
          4931 => x"08",
          4932 => x"89",
          4933 => x"16",
          4934 => x"82",
          4935 => x"08",
          4936 => x"88",
          4937 => x"74",
          4938 => x"04",
          4939 => x"53",
          4940 => x"3f",
          4941 => x"ea",
          4942 => x"6a",
          4943 => x"d8",
          4944 => x"3f",
          4945 => x"0d",
          4946 => x"05",
          4947 => x"72",
          4948 => x"ff",
          4949 => x"ff",
          4950 => x"2e",
          4951 => x"2e",
          4952 => x"72",
          4953 => x"83",
          4954 => x"ff",
          4955 => x"ec",
          4956 => x"81",
          4957 => x"51",
          4958 => x"0d",
          4959 => x"22",
          4960 => x"51",
          4961 => x"38",
          4962 => x"2e",
          4963 => x"ff",
          4964 => x"ec",
          4965 => x"e0",
          4966 => x"3d",
          4967 => x"26",
          4968 => x"06",
          4969 => x"72",
          4970 => x"75",
          4971 => x"70",
          4972 => x"52",
          4973 => x"82",
          4974 => x"81",
          4975 => x"53",
          4976 => x"88",
          4977 => x"82",
          4978 => x"71",
          4979 => x"54",
          4980 => x"31",
          4981 => x"a4",
          4982 => x"12",
          4983 => x"39",
          4984 => x"51",
          4985 => x"39",
          4986 => x"ff",
          4987 => x"38",
          4988 => x"71",
          4989 => x"3d",
          4990 => x"00",
          4991 => x"ff",
          4992 => x"00",
          4993 => x"00",
          4994 => x"00",
          4995 => x"00",
          4996 => x"00",
          4997 => x"00",
          4998 => x"00",
          4999 => x"00",
          5000 => x"00",
          5001 => x"00",
          5002 => x"00",
          5003 => x"00",
          5004 => x"00",
          5005 => x"00",
          5006 => x"00",
          5007 => x"00",
          5008 => x"00",
          5009 => x"00",
          5010 => x"00",
          5011 => x"00",
          5012 => x"00",
          5013 => x"00",
          5014 => x"00",
          5015 => x"00",
          5016 => x"00",
          5017 => x"00",
          5018 => x"00",
          5019 => x"00",
          5020 => x"00",
          5021 => x"00",
          5022 => x"00",
          5023 => x"00",
          5024 => x"00",
          5025 => x"00",
          5026 => x"00",
          5027 => x"00",
          5028 => x"00",
          5029 => x"00",
          5030 => x"00",
          5031 => x"00",
          5032 => x"00",
          5033 => x"00",
          5034 => x"00",
          5035 => x"00",
          5036 => x"00",
          5037 => x"00",
          5038 => x"00",
          5039 => x"00",
          5040 => x"00",
          5041 => x"00",
          5042 => x"00",
          5043 => x"00",
          5044 => x"00",
          5045 => x"00",
          5046 => x"00",
          5047 => x"00",
          5048 => x"00",
          5049 => x"00",
          5050 => x"00",
          5051 => x"00",
          5052 => x"00",
          5053 => x"00",
          5054 => x"00",
          5055 => x"00",
          5056 => x"00",
          5057 => x"00",
          5058 => x"00",
          5059 => x"00",
          5060 => x"00",
          5061 => x"00",
          5062 => x"00",
          5063 => x"00",
          5064 => x"69",
          5065 => x"69",
          5066 => x"69",
          5067 => x"6c",
          5068 => x"65",
          5069 => x"63",
          5070 => x"63",
          5071 => x"64",
          5072 => x"64",
          5073 => x"65",
          5074 => x"65",
          5075 => x"69",
          5076 => x"66",
          5077 => x"00",
          5078 => x"65",
          5079 => x"65",
          5080 => x"6e",
          5081 => x"62",
          5082 => x"62",
          5083 => x"69",
          5084 => x"64",
          5085 => x"45",
          5086 => x"6e",
          5087 => x"65",
          5088 => x"69",
          5089 => x"72",
          5090 => x"6f",
          5091 => x"6f",
          5092 => x"6f",
          5093 => x"6f",
          5094 => x"6e",
          5095 => x"69",
          5096 => x"00",
          5097 => x"73",
          5098 => x"2e",
          5099 => x"61",
          5100 => x"65",
          5101 => x"00",
          5102 => x"68",
          5103 => x"6e",
          5104 => x"00",
          5105 => x"20",
          5106 => x"72",
          5107 => x"2e",
          5108 => x"20",
          5109 => x"69",
          5110 => x"69",
          5111 => x"69",
          5112 => x"65",
          5113 => x"00",
          5114 => x"6d",
          5115 => x"20",
          5116 => x"74",
          5117 => x"64",
          5118 => x"6b",
          5119 => x"74",
          5120 => x"64",
          5121 => x"75",
          5122 => x"61",
          5123 => x"6e",
          5124 => x"00",
          5125 => x"69",
          5126 => x"64",
          5127 => x"66",
          5128 => x"6d",
          5129 => x"00",
          5130 => x"61",
          5131 => x"20",
          5132 => x"00",
          5133 => x"65",
          5134 => x"63",
          5135 => x"00",
          5136 => x"73",
          5137 => x"6e",
          5138 => x"72",
          5139 => x"25",
          5140 => x"73",
          5141 => x"25",
          5142 => x"73",
          5143 => x"00",
          5144 => x"00",
          5145 => x"00",
          5146 => x"30",
          5147 => x"20",
          5148 => x"00",
          5149 => x"00",
          5150 => x"7c",
          5151 => x"4f",
          5152 => x"20",
          5153 => x"2f",
          5154 => x"31",
          5155 => x"5a",
          5156 => x"20",
          5157 => x"73",
          5158 => x"0a",
          5159 => x"6e",
          5160 => x"20",
          5161 => x"00",
          5162 => x"20",
          5163 => x"70",
          5164 => x"6e",
          5165 => x"00",
          5166 => x"20",
          5167 => x"72",
          5168 => x"4f",
          5169 => x"69",
          5170 => x"74",
          5171 => x"20",
          5172 => x"72",
          5173 => x"41",
          5174 => x"69",
          5175 => x"74",
          5176 => x"20",
          5177 => x"72",
          5178 => x"41",
          5179 => x"69",
          5180 => x"74",
          5181 => x"6e",
          5182 => x"6d",
          5183 => x"6e",
          5184 => x"74",
          5185 => x"00",
          5186 => x"78",
          5187 => x"00",
          5188 => x"70",
          5189 => x"3a",
          5190 => x"64",
          5191 => x"74",
          5192 => x"73",
          5193 => x"30",
          5194 => x"65",
          5195 => x"61",
          5196 => x"00",
          5197 => x"6c",
          5198 => x"2e",
          5199 => x"6f",
          5200 => x"2e",
          5201 => x"72",
          5202 => x"00",
          5203 => x"28",
          5204 => x"25",
          5205 => x"38",
          5206 => x"75",
          5207 => x"72",
          5208 => x"6c",
          5209 => x"30",
          5210 => x"58",
          5211 => x"30",
          5212 => x"58",
          5213 => x"20",
          5214 => x"00",
          5215 => x"74",
          5216 => x"65",
          5217 => x"78",
          5218 => x"61",
          5219 => x"6f",
          5220 => x"38",
          5221 => x"00",
          5222 => x"72",
          5223 => x"20",
          5224 => x"64",
          5225 => x"65",
          5226 => x"67",
          5227 => x"61",
          5228 => x"00",
          5229 => x"72",
          5230 => x"67",
          5231 => x"50",
          5232 => x"64",
          5233 => x"2e",
          5234 => x"64",
          5235 => x"00",
          5236 => x"73",
          5237 => x"6f",
          5238 => x"00",
          5239 => x"79",
          5240 => x"74",
          5241 => x"6e",
          5242 => x"65",
          5243 => x"61",
          5244 => x"75",
          5245 => x"2e",
          5246 => x"69",
          5247 => x"72",
          5248 => x"2e",
          5249 => x"2f",
          5250 => x"64",
          5251 => x"64",
          5252 => x"6f",
          5253 => x"74",
          5254 => x"28",
          5255 => x"43",
          5256 => x"29",
          5257 => x"69",
          5258 => x"6c",
          5259 => x"3a",
          5260 => x"42",
          5261 => x"20",
          5262 => x"30",
          5263 => x"20",
          5264 => x"20",
          5265 => x"38",
          5266 => x"2e",
          5267 => x"4e",
          5268 => x"20",
          5269 => x"30",
          5270 => x"20",
          5271 => x"20",
          5272 => x"38",
          5273 => x"2e",
          5274 => x"41",
          5275 => x"20",
          5276 => x"30",
          5277 => x"20",
          5278 => x"52",
          5279 => x"76",
          5280 => x"30",
          5281 => x"20",
          5282 => x"31",
          5283 => x"6d",
          5284 => x"30",
          5285 => x"20",
          5286 => x"43",
          5287 => x"61",
          5288 => x"30",
          5289 => x"20",
          5290 => x"4f",
          5291 => x"00",
          5292 => x"42",
          5293 => x"20",
          5294 => x"00",
          5295 => x"53",
          5296 => x"50",
          5297 => x"73",
          5298 => x"20",
          5299 => x"65",
          5300 => x"74",
          5301 => x"65",
          5302 => x"38",
          5303 => x"20",
          5304 => x"65",
          5305 => x"61",
          5306 => x"65",
          5307 => x"38",
          5308 => x"20",
          5309 => x"20",
          5310 => x"64",
          5311 => x"20",
          5312 => x"38",
          5313 => x"69",
          5314 => x"20",
          5315 => x"64",
          5316 => x"20",
          5317 => x"20",
          5318 => x"34",
          5319 => x"20",
          5320 => x"6d",
          5321 => x"46",
          5322 => x"20",
          5323 => x"2e",
          5324 => x"0a",
          5325 => x"44",
          5326 => x"63",
          5327 => x"20",
          5328 => x"3d",
          5329 => x"64",
          5330 => x"20",
          5331 => x"6f",
          5332 => x"4d",
          5333 => x"46",
          5334 => x"2e",
          5335 => x"0a",
          5336 => x"00",
          5337 => x"6d",
          5338 => x"00",
          5339 => x"56",
          5340 => x"6e",
          5341 => x"00",
          5342 => x"00",
          5343 => x"00",
          5344 => x"00",
          5345 => x"00",
          5346 => x"00",
          5347 => x"00",
          5348 => x"00",
          5349 => x"00",
          5350 => x"00",
          5351 => x"00",
          5352 => x"00",
          5353 => x"00",
          5354 => x"00",
          5355 => x"00",
          5356 => x"00",
          5357 => x"00",
          5358 => x"00",
          5359 => x"00",
          5360 => x"00",
          5361 => x"00",
          5362 => x"00",
          5363 => x"00",
          5364 => x"00",
          5365 => x"00",
          5366 => x"00",
          5367 => x"00",
          5368 => x"00",
          5369 => x"00",
          5370 => x"00",
          5371 => x"00",
          5372 => x"00",
          5373 => x"00",
          5374 => x"5b",
          5375 => x"5b",
          5376 => x"5b",
          5377 => x"5b",
          5378 => x"5b",
          5379 => x"5b",
          5380 => x"00",
          5381 => x"00",
          5382 => x"00",
          5383 => x"00",
          5384 => x"00",
          5385 => x"69",
          5386 => x"69",
          5387 => x"00",
          5388 => x"20",
          5389 => x"61",
          5390 => x"20",
          5391 => x"68",
          5392 => x"72",
          5393 => x"74",
          5394 => x"00",
          5395 => x"74",
          5396 => x"72",
          5397 => x"73",
          5398 => x"6c",
          5399 => x"62",
          5400 => x"44",
          5401 => x"3f",
          5402 => x"2c",
          5403 => x"41",
          5404 => x"00",
          5405 => x"44",
          5406 => x"4f",
          5407 => x"20",
          5408 => x"20",
          5409 => x"4d",
          5410 => x"54",
          5411 => x"00",
          5412 => x"00",
          5413 => x"03",
          5414 => x"16",
          5415 => x"9a",
          5416 => x"45",
          5417 => x"92",
          5418 => x"99",
          5419 => x"49",
          5420 => x"a9",
          5421 => x"b1",
          5422 => x"b9",
          5423 => x"c1",
          5424 => x"c9",
          5425 => x"d1",
          5426 => x"d9",
          5427 => x"e1",
          5428 => x"e9",
          5429 => x"f1",
          5430 => x"f9",
          5431 => x"2e",
          5432 => x"22",
          5433 => x"00",
          5434 => x"10",
          5435 => x"00",
          5436 => x"04",
          5437 => x"00",
          5438 => x"e9",
          5439 => x"e5",
          5440 => x"e8",
          5441 => x"c4",
          5442 => x"c6",
          5443 => x"fb",
          5444 => x"dc",
          5445 => x"a7",
          5446 => x"f3",
          5447 => x"aa",
          5448 => x"ac",
          5449 => x"ab",
          5450 => x"93",
          5451 => x"62",
          5452 => x"51",
          5453 => x"5b",
          5454 => x"2c",
          5455 => x"5e",
          5456 => x"69",
          5457 => x"6c",
          5458 => x"65",
          5459 => x"53",
          5460 => x"0c",
          5461 => x"90",
          5462 => x"93",
          5463 => x"b5",
          5464 => x"a9",
          5465 => x"b5",
          5466 => x"65",
          5467 => x"f7",
          5468 => x"b7",
          5469 => x"a0",
          5470 => x"e0",
          5471 => x"ff",
          5472 => x"30",
          5473 => x"10",
          5474 => x"06",
          5475 => x"81",
          5476 => x"84",
          5477 => x"89",
          5478 => x"8d",
          5479 => x"91",
          5480 => x"f6",
          5481 => x"98",
          5482 => x"9d",
          5483 => x"a0",
          5484 => x"a4",
          5485 => x"a9",
          5486 => x"ac",
          5487 => x"b1",
          5488 => x"b5",
          5489 => x"b8",
          5490 => x"bc",
          5491 => x"c1",
          5492 => x"c5",
          5493 => x"c7",
          5494 => x"cd",
          5495 => x"8e",
          5496 => x"03",
          5497 => x"f8",
          5498 => x"3a",
          5499 => x"3b",
          5500 => x"40",
          5501 => x"0a",
          5502 => x"86",
          5503 => x"58",
          5504 => x"5c",
          5505 => x"93",
          5506 => x"64",
          5507 => x"97",
          5508 => x"6c",
          5509 => x"70",
          5510 => x"74",
          5511 => x"78",
          5512 => x"7c",
          5513 => x"a6",
          5514 => x"84",
          5515 => x"ae",
          5516 => x"45",
          5517 => x"90",
          5518 => x"03",
          5519 => x"ac",
          5520 => x"89",
          5521 => x"c2",
          5522 => x"c4",
          5523 => x"8c",
          5524 => x"18",
          5525 => x"f3",
          5526 => x"f7",
          5527 => x"fa",
          5528 => x"10",
          5529 => x"36",
          5530 => x"01",
          5531 => x"61",
          5532 => x"7d",
          5533 => x"96",
          5534 => x"08",
          5535 => x"08",
          5536 => x"06",
          5537 => x"52",
          5538 => x"56",
          5539 => x"70",
          5540 => x"c8",
          5541 => x"da",
          5542 => x"ea",
          5543 => x"80",
          5544 => x"a0",
          5545 => x"b8",
          5546 => x"cc",
          5547 => x"02",
          5548 => x"01",
          5549 => x"fc",
          5550 => x"70",
          5551 => x"83",
          5552 => x"2f",
          5553 => x"06",
          5554 => x"64",
          5555 => x"1a",
          5556 => x"00",
          5557 => x"00",
          5558 => x"00",
          5559 => x"00",
          5560 => x"00",
          5561 => x"00",
          5562 => x"00",
          5563 => x"00",
          5564 => x"00",
          5565 => x"00",
          5566 => x"00",
          5567 => x"00",
          5568 => x"00",
          5569 => x"00",
          5570 => x"00",
          5571 => x"00",
          5572 => x"00",
          5573 => x"00",
          5574 => x"00",
          5575 => x"00",
          5576 => x"00",
          5577 => x"00",
          5578 => x"00",
          5579 => x"00",
          5580 => x"00",
          5581 => x"00",
          5582 => x"00",
          5583 => x"00",
          5584 => x"00",
          5585 => x"00",
          5586 => x"00",
          5587 => x"00",
          5588 => x"00",
          5589 => x"00",
          5590 => x"00",
          5591 => x"00",
          5592 => x"00",
          5593 => x"00",
          5594 => x"00",
          5595 => x"00",
          5596 => x"00",
          5597 => x"00",
          5598 => x"00",
          5599 => x"00",
          5600 => x"00",
          5601 => x"00",
          5602 => x"00",
          5603 => x"00",
          5604 => x"00",
          5605 => x"00",
          5606 => x"00",
          5607 => x"00",
          5608 => x"00",
          5609 => x"00",
          5610 => x"81",
          5611 => x"7f",
          5612 => x"00",
          5613 => x"00",
          5614 => x"f5",
          5615 => x"00",
          5616 => x"01",
          5617 => x"00",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"00",
          5630 => x"00",
          5631 => x"00",
          5632 => x"00",
          5633 => x"00",
          5634 => x"03",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"08",
             6 => x"04",
             7 => x"00",
             8 => x"71",
             9 => x"81",
            10 => x"ff",
            11 => x"00",
            12 => x"71",
            13 => x"83",
            14 => x"2b",
            15 => x"0b",
            16 => x"72",
            17 => x"09",
            18 => x"07",
            19 => x"00",
            20 => x"72",
            21 => x"51",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"09",
            26 => x"0a",
            27 => x"51",
            28 => x"72",
            29 => x"51",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"0b",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"72",
            45 => x"0b",
            46 => x"00",
            47 => x"00",
            48 => x"72",
            49 => x"09",
            50 => x"06",
            51 => x"00",
            52 => x"71",
            53 => x"06",
            54 => x"0b",
            55 => x"51",
            56 => x"72",
            57 => x"81",
            58 => x"51",
            59 => x"00",
            60 => x"72",
            61 => x"81",
            62 => x"53",
            63 => x"00",
            64 => x"71",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"72",
            69 => x"04",
            70 => x"00",
            71 => x"00",
            72 => x"72",
            73 => x"07",
            74 => x"00",
            75 => x"00",
            76 => x"71",
            77 => x"81",
            78 => x"81",
            79 => x"00",
            80 => x"71",
            81 => x"ec",
            82 => x"06",
            83 => x"00",
            84 => x"88",
            85 => x"0b",
            86 => x"88",
            87 => x"0c",
            88 => x"88",
            89 => x"0b",
            90 => x"88",
            91 => x"0c",
            92 => x"72",
            93 => x"81",
            94 => x"73",
            95 => x"07",
            96 => x"72",
            97 => x"09",
            98 => x"06",
            99 => x"06",
           100 => x"05",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"04",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"71",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"04",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"02",
           117 => x"04",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"02",
           126 => x"ff",
           127 => x"ff",
           128 => x"00",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"96",
           135 => x"0b",
           136 => x"0b",
           137 => x"d6",
           138 => x"0b",
           139 => x"0b",
           140 => x"98",
           141 => x"0b",
           142 => x"0b",
           143 => x"da",
           144 => x"0b",
           145 => x"0b",
           146 => x"9e",
           147 => x"0b",
           148 => x"0b",
           149 => x"e2",
           150 => x"0b",
           151 => x"0b",
           152 => x"a6",
           153 => x"0b",
           154 => x"0b",
           155 => x"ea",
           156 => x"0b",
           157 => x"0b",
           158 => x"ae",
           159 => x"0b",
           160 => x"0b",
           161 => x"f2",
           162 => x"0b",
           163 => x"0b",
           164 => x"b6",
           165 => x"0b",
           166 => x"0b",
           167 => x"fa",
           168 => x"0b",
           169 => x"0b",
           170 => x"be",
           171 => x"0b",
           172 => x"0b",
           173 => x"82",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"0c",
           194 => x"08",
           195 => x"a4",
           196 => x"08",
           197 => x"a4",
           198 => x"08",
           199 => x"a4",
           200 => x"08",
           201 => x"a4",
           202 => x"08",
           203 => x"a4",
           204 => x"08",
           205 => x"a4",
           206 => x"a4",
           207 => x"e0",
           208 => x"e0",
           209 => x"82",
           210 => x"e0",
           211 => x"82",
           212 => x"e0",
           213 => x"82",
           214 => x"e0",
           215 => x"82",
           216 => x"82",
           217 => x"04",
           218 => x"2d",
           219 => x"90",
           220 => x"dd",
           221 => x"80",
           222 => x"fd",
           223 => x"c0",
           224 => x"80",
           225 => x"80",
           226 => x"0c",
           227 => x"08",
           228 => x"a4",
           229 => x"a4",
           230 => x"e0",
           231 => x"e0",
           232 => x"82",
           233 => x"82",
           234 => x"04",
           235 => x"2d",
           236 => x"90",
           237 => x"ce",
           238 => x"80",
           239 => x"82",
           240 => x"c0",
           241 => x"82",
           242 => x"80",
           243 => x"0c",
           244 => x"08",
           245 => x"a4",
           246 => x"a4",
           247 => x"e0",
           248 => x"e0",
           249 => x"82",
           250 => x"82",
           251 => x"04",
           252 => x"2d",
           253 => x"90",
           254 => x"cd",
           255 => x"80",
           256 => x"9b",
           257 => x"c0",
           258 => x"82",
           259 => x"80",
           260 => x"0c",
           261 => x"08",
           262 => x"a4",
           263 => x"a4",
           264 => x"e0",
           265 => x"e0",
           266 => x"82",
           267 => x"82",
           268 => x"04",
           269 => x"2d",
           270 => x"90",
           271 => x"99",
           272 => x"80",
           273 => x"a2",
           274 => x"c0",
           275 => x"81",
           276 => x"80",
           277 => x"0c",
           278 => x"08",
           279 => x"a4",
           280 => x"a4",
           281 => x"e0",
           282 => x"e0",
           283 => x"82",
           284 => x"82",
           285 => x"04",
           286 => x"2d",
           287 => x"90",
           288 => x"d9",
           289 => x"80",
           290 => x"fb",
           291 => x"c0",
           292 => x"80",
           293 => x"80",
           294 => x"0c",
           295 => x"08",
           296 => x"a4",
           297 => x"a4",
           298 => x"e0",
           299 => x"e0",
           300 => x"82",
           301 => x"82",
           302 => x"04",
           303 => x"2d",
           304 => x"90",
           305 => x"89",
           306 => x"80",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"10",
           311 => x"00",
           312 => x"09",
           313 => x"2b",
           314 => x"04",
           315 => x"05",
           316 => x"72",
           317 => x"51",
           318 => x"70",
           319 => x"71",
           320 => x"0b",
           321 => x"fa",
           322 => x"02",
           323 => x"82",
           324 => x"e0",
           325 => x"a4",
           326 => x"a4",
           327 => x"fc",
           328 => x"e0",
           329 => x"f8",
           330 => x"05",
           331 => x"54",
           332 => x"04",
           333 => x"a4",
           334 => x"08",
           335 => x"81",
           336 => x"52",
           337 => x"a4",
           338 => x"8d",
           339 => x"f4",
           340 => x"a4",
           341 => x"e0",
           342 => x"82",
           343 => x"e0",
           344 => x"a4",
           345 => x"08",
           346 => x"38",
           347 => x"05",
           348 => x"a4",
           349 => x"3f",
           350 => x"a4",
           351 => x"a4",
           352 => x"81",
           353 => x"a4",
           354 => x"82",
           355 => x"e0",
           356 => x"71",
           357 => x"05",
           358 => x"8c",
           359 => x"05",
           360 => x"fc",
           361 => x"a4",
           362 => x"34",
           363 => x"70",
           364 => x"52",
           365 => x"82",
           366 => x"e0",
           367 => x"02",
           368 => x"86",
           369 => x"34",
           370 => x"82",
           371 => x"0a",
           372 => x"0c",
           373 => x"82",
           374 => x"e0",
           375 => x"e0",
           376 => x"e0",
           377 => x"54",
           378 => x"70",
           379 => x"82",
           380 => x"e0",
           381 => x"54",
           382 => x"dc",
           383 => x"54",
           384 => x"04",
           385 => x"a4",
           386 => x"08",
           387 => x"fc",
           388 => x"05",
           389 => x"05",
           390 => x"05",
           391 => x"98",
           392 => x"05",
           393 => x"08",
           394 => x"87",
           395 => x"82",
           396 => x"0c",
           397 => x"a4",
           398 => x"08",
           399 => x"14",
           400 => x"08",
           401 => x"81",
           402 => x"51",
           403 => x"0b",
           404 => x"96",
           405 => x"05",
           406 => x"e0",
           407 => x"ff",
           408 => x"38",
           409 => x"81",
           410 => x"0c",
           411 => x"70",
           412 => x"95",
           413 => x"05",
           414 => x"38",
           415 => x"53",
           416 => x"e0",
           417 => x"b0",
           418 => x"82",
           419 => x"98",
           420 => x"72",
           421 => x"05",
           422 => x"70",
           423 => x"80",
           424 => x"e4",
           425 => x"53",
           426 => x"23",
           427 => x"e8",
           428 => x"2c",
           429 => x"11",
           430 => x"72",
           431 => x"82",
           432 => x"82",
           433 => x"15",
           434 => x"e0",
           435 => x"a4",
           436 => x"70",
           437 => x"25",
           438 => x"a4",
           439 => x"08",
           440 => x"81",
           441 => x"38",
           442 => x"70",
           443 => x"2c",
           444 => x"53",
           445 => x"23",
           446 => x"e4",
           447 => x"06",
           448 => x"38",
           449 => x"70",
           450 => x"53",
           451 => x"a4",
           452 => x"08",
           453 => x"a4",
           454 => x"a4",
           455 => x"92",
           456 => x"05",
           457 => x"11",
           458 => x"04",
           459 => x"70",
           460 => x"a4",
           461 => x"08",
           462 => x"53",
           463 => x"23",
           464 => x"e4",
           465 => x"53",
           466 => x"23",
           467 => x"e4",
           468 => x"53",
           469 => x"23",
           470 => x"e4",
           471 => x"72",
           472 => x"80",
           473 => x"34",
           474 => x"e4",
           475 => x"72",
           476 => x"fb",
           477 => x"08",
           478 => x"ec",
           479 => x"82",
           480 => x"e3",
           481 => x"34",
           482 => x"90",
           483 => x"05",
           484 => x"90",
           485 => x"82",
           486 => x"e0",
           487 => x"51",
           488 => x"05",
           489 => x"08",
           490 => x"90",
           491 => x"08",
           492 => x"a4",
           493 => x"08",
           494 => x"81",
           495 => x"2e",
           496 => x"05",
           497 => x"2c",
           498 => x"08",
           499 => x"98",
           500 => x"f4",
           501 => x"08",
           502 => x"82",
           503 => x"a4",
           504 => x"08",
           505 => x"08",
           506 => x"54",
           507 => x"23",
           508 => x"90",
           509 => x"05",
           510 => x"90",
           511 => x"08",
           512 => x"e4",
           513 => x"06",
           514 => x"ab",
           515 => x"33",
           516 => x"53",
           517 => x"52",
           518 => x"08",
           519 => x"05",
           520 => x"fc",
           521 => x"e0",
           522 => x"08",
           523 => x"ec",
           524 => x"f4",
           525 => x"72",
           526 => x"8a",
           527 => x"05",
           528 => x"51",
           529 => x"82",
           530 => x"e0",
           531 => x"82",
           532 => x"08",
           533 => x"53",
           534 => x"05",
           535 => x"08",
           536 => x"05",
           537 => x"dc",
           538 => x"dc",
           539 => x"05",
           540 => x"08",
           541 => x"08",
           542 => x"53",
           543 => x"23",
           544 => x"30",
           545 => x"82",
           546 => x"ff",
           547 => x"a4",
           548 => x"88",
           549 => x"23",
           550 => x"05",
           551 => x"72",
           552 => x"80",
           553 => x"05",
           554 => x"f4",
           555 => x"05",
           556 => x"51",
           557 => x"82",
           558 => x"e0",
           559 => x"82",
           560 => x"08",
           561 => x"53",
           562 => x"05",
           563 => x"08",
           564 => x"05",
           565 => x"d8",
           566 => x"d8",
           567 => x"05",
           568 => x"22",
           569 => x"e0",
           570 => x"a8",
           571 => x"0c",
           572 => x"82",
           573 => x"e0",
           574 => x"70",
           575 => x"82",
           576 => x"82",
           577 => x"e0",
           578 => x"a4",
           579 => x"53",
           580 => x"a4",
           581 => x"54",
           582 => x"70",
           583 => x"82",
           584 => x"39",
           585 => x"53",
           586 => x"82",
           587 => x"e0",
           588 => x"e0",
           589 => x"82",
           590 => x"05",
           591 => x"82",
           592 => x"53",
           593 => x"52",
           594 => x"08",
           595 => x"0c",
           596 => x"08",
           597 => x"82",
           598 => x"e0",
           599 => x"75",
           600 => x"08",
           601 => x"e4",
           602 => x"72",
           603 => x"08",
           604 => x"72",
           605 => x"82",
           606 => x"86",
           607 => x"72",
           608 => x"a4",
           609 => x"82",
           610 => x"e0",
           611 => x"82",
           612 => x"e0",
           613 => x"72",
           614 => x"82",
           615 => x"05",
           616 => x"05",
           617 => x"cc",
           618 => x"e0",
           619 => x"a4",
           620 => x"08",
           621 => x"e4",
           622 => x"06",
           623 => x"d0",
           624 => x"33",
           625 => x"e0",
           626 => x"51",
           627 => x"e0",
           628 => x"06",
           629 => x"e4",
           630 => x"08",
           631 => x"08",
           632 => x"54",
           633 => x"34",
           634 => x"70",
           635 => x"53",
           636 => x"a4",
           637 => x"70",
           638 => x"2c",
           639 => x"82",
           640 => x"75",
           641 => x"08",
           642 => x"a4",
           643 => x"70",
           644 => x"2c",
           645 => x"82",
           646 => x"75",
           647 => x"08",
           648 => x"e4",
           649 => x"53",
           650 => x"ec",
           651 => x"82",
           652 => x"90",
           653 => x"73",
           654 => x"88",
           655 => x"3f",
           656 => x"05",
           657 => x"51",
           658 => x"82",
           659 => x"ad",
           660 => x"82",
           661 => x"84",
           662 => x"72",
           663 => x"08",
           664 => x"a5",
           665 => x"e4",
           666 => x"06",
           667 => x"38",
           668 => x"52",
           669 => x"a4",
           670 => x"70",
           671 => x"2e",
           672 => x"05",
           673 => x"82",
           674 => x"72",
           675 => x"82",
           676 => x"82",
           677 => x"89",
           678 => x"05",
           679 => x"51",
           680 => x"82",
           681 => x"11",
           682 => x"ec",
           683 => x"2c",
           684 => x"82",
           685 => x"b0",
           686 => x"e0",
           687 => x"2a",
           688 => x"80",
           689 => x"e8",
           690 => x"82",
           691 => x"98",
           692 => x"73",
           693 => x"88",
           694 => x"3f",
           695 => x"05",
           696 => x"51",
           697 => x"a4",
           698 => x"54",
           699 => x"23",
           700 => x"53",
           701 => x"a4",
           702 => x"87",
           703 => x"08",
           704 => x"2e",
           705 => x"a4",
           706 => x"a4",
           707 => x"3f",
           708 => x"f8",
           709 => x"09",
           710 => x"a4",
           711 => x"53",
           712 => x"23",
           713 => x"83",
           714 => x"e0",
           715 => x"e0",
           716 => x"52",
           717 => x"81",
           718 => x"0c",
           719 => x"82",
           720 => x"72",
           721 => x"cb",
           722 => x"22",
           723 => x"a4",
           724 => x"ff",
           725 => x"80",
           726 => x"05",
           727 => x"05",
           728 => x"3f",
           729 => x"81",
           730 => x"0c",
           731 => x"f0",
           732 => x"38",
           733 => x"52",
           734 => x"ff",
           735 => x"0c",
           736 => x"70",
           737 => x"39",
           738 => x"70",
           739 => x"53",
           740 => x"e0",
           741 => x"54",
           742 => x"05",
           743 => x"51",
           744 => x"e0",
           745 => x"51",
           746 => x"a4",
           747 => x"a4",
           748 => x"3f",
           749 => x"05",
           750 => x"08",
           751 => x"09",
           752 => x"e0",
           753 => x"82",
           754 => x"0b",
           755 => x"8a",
           756 => x"23",
           757 => x"88",
           758 => x"f8",
           759 => x"ea",
           760 => x"08",
           761 => x"08",
           762 => x"a4",
           763 => x"0c",
           764 => x"04",
           765 => x"a4",
           766 => x"08",
           767 => x"08",
           768 => x"08",
           769 => x"08",
           770 => x"3d",
           771 => x"e0",
           772 => x"fb",
           773 => x"08",
           774 => x"85",
           775 => x"32",
           776 => x"53",
           777 => x"82",
           778 => x"92",
           779 => x"08",
           780 => x"88",
           781 => x"08",
           782 => x"a4",
           783 => x"06",
           784 => x"fb",
           785 => x"82",
           786 => x"90",
           787 => x"e0",
           788 => x"b1",
           789 => x"f8",
           790 => x"fc",
           791 => x"8a",
           792 => x"82",
           793 => x"8a",
           794 => x"f8",
           795 => x"05",
           796 => x"05",
           797 => x"05",
           798 => x"0d",
           799 => x"a4",
           800 => x"3d",
           801 => x"f8",
           802 => x"05",
           803 => x"70",
           804 => x"51",
           805 => x"ff",
           806 => x"0c",
           807 => x"88",
           808 => x"a4",
           809 => x"e0",
           810 => x"82",
           811 => x"81",
           812 => x"38",
           813 => x"82",
           814 => x"82",
           815 => x"90",
           816 => x"e0",
           817 => x"ab",
           818 => x"f8",
           819 => x"a4",
           820 => x"a4",
           821 => x"a4",
           822 => x"0c",
           823 => x"04",
           824 => x"a4",
           825 => x"08",
           826 => x"08",
           827 => x"70",
           828 => x"0d",
           829 => x"a4",
           830 => x"3d",
           831 => x"08",
           832 => x"81",
           833 => x"51",
           834 => x"0b",
           835 => x"81",
           836 => x"05",
           837 => x"70",
           838 => x"80",
           839 => x"08",
           840 => x"8c",
           841 => x"88",
           842 => x"a4",
           843 => x"82",
           844 => x"57",
           845 => x"81",
           846 => x"8c",
           847 => x"8c",
           848 => x"05",
           849 => x"05",
           850 => x"e0",
           851 => x"a4",
           852 => x"a4",
           853 => x"06",
           854 => x"72",
           855 => x"a3",
           856 => x"08",
           857 => x"0c",
           858 => x"70",
           859 => x"51",
           860 => x"a4",
           861 => x"08",
           862 => x"87",
           863 => x"82",
           864 => x"0c",
           865 => x"88",
           866 => x"32",
           867 => x"71",
           868 => x"e0",
           869 => x"39",
           870 => x"85",
           871 => x"06",
           872 => x"80",
           873 => x"05",
           874 => x"08",
           875 => x"bf",
           876 => x"82",
           877 => x"11",
           878 => x"e0",
           879 => x"33",
           880 => x"0c",
           881 => x"e0",
           882 => x"33",
           883 => x"51",
           884 => x"38",
           885 => x"70",
           886 => x"fc",
           887 => x"08",
           888 => x"a4",
           889 => x"08",
           890 => x"33",
           891 => x"14",
           892 => x"f8",
           893 => x"a4",
           894 => x"05",
           895 => x"e0",
           896 => x"a4",
           897 => x"08",
           898 => x"08",
           899 => x"0c",
           900 => x"08",
           901 => x"a4",
           902 => x"08",
           903 => x"88",
           904 => x"a4",
           905 => x"a4",
           906 => x"81",
           907 => x"f0",
           908 => x"e0",
           909 => x"82",
           910 => x"07",
           911 => x"05",
           912 => x"08",
           913 => x"33",
           914 => x"a4",
           915 => x"e0",
           916 => x"08",
           917 => x"a4",
           918 => x"06",
           919 => x"0c",
           920 => x"f8",
           921 => x"3d",
           922 => x"e0",
           923 => x"fd",
           924 => x"05",
           925 => x"0c",
           926 => x"82",
           927 => x"e0",
           928 => x"82",
           929 => x"05",
           930 => x"08",
           931 => x"08",
           932 => x"90",
           933 => x"08",
           934 => x"38",
           935 => x"82",
           936 => x"82",
           937 => x"e0",
           938 => x"a4",
           939 => x"a4",
           940 => x"08",
           941 => x"a4",
           942 => x"08",
           943 => x"a4",
           944 => x"08",
           945 => x"38",
           946 => x"ff",
           947 => x"0c",
           948 => x"ff",
           949 => x"0c",
           950 => x"82",
           951 => x"51",
           952 => x"82",
           953 => x"05",
           954 => x"82",
           955 => x"05",
           956 => x"82",
           957 => x"2e",
           958 => x"05",
           959 => x"08",
           960 => x"a4",
           961 => x"08",
           962 => x"34",
           963 => x"81",
           964 => x"0c",
           965 => x"88",
           966 => x"51",
           967 => x"04",
           968 => x"a4",
           969 => x"08",
           970 => x"fc",
           971 => x"05",
           972 => x"08",
           973 => x"a4",
           974 => x"06",
           975 => x"da",
           976 => x"08",
           977 => x"05",
           978 => x"08",
           979 => x"31",
           980 => x"3d",
           981 => x"e0",
           982 => x"fe",
           983 => x"05",
           984 => x"0c",
           985 => x"52",
           986 => x"05",
           987 => x"8c",
           988 => x"05",
           989 => x"e0",
           990 => x"82",
           991 => x"81",
           992 => x"38",
           993 => x"88",
           994 => x"51",
           995 => x"04",
           996 => x"a4",
           997 => x"08",
           998 => x"fc",
           999 => x"05",
          1000 => x"0c",
          1001 => x"80",
          1002 => x"08",
          1003 => x"a4",
          1004 => x"08",
          1005 => x"a4",
          1006 => x"08",
          1007 => x"82",
          1008 => x"70",
          1009 => x"08",
          1010 => x"05",
          1011 => x"08",
          1012 => x"a4",
          1013 => x"e0",
          1014 => x"39",
          1015 => x"70",
          1016 => x"0d",
          1017 => x"a4",
          1018 => x"3d",
          1019 => x"08",
          1020 => x"a4",
          1021 => x"82",
          1022 => x"05",
          1023 => x"82",
          1024 => x"33",
          1025 => x"51",
          1026 => x"39",
          1027 => x"52",
          1028 => x"05",
          1029 => x"88",
          1030 => x"51",
          1031 => x"a4",
          1032 => x"82",
          1033 => x"05",
          1034 => x"82",
          1035 => x"2e",
          1036 => x"a4",
          1037 => x"e8",
          1038 => x"08",
          1039 => x"ff",
          1040 => x"0c",
          1041 => x"8c",
          1042 => x"08",
          1043 => x"8c",
          1044 => x"8c",
          1045 => x"fc",
          1046 => x"08",
          1047 => x"a4",
          1048 => x"71",
          1049 => x"05",
          1050 => x"39",
          1051 => x"05",
          1052 => x"08",
          1053 => x"82",
          1054 => x"08",
          1055 => x"0d",
          1056 => x"52",
          1057 => x"51",
          1058 => x"70",
          1059 => x"82",
          1060 => x"05",
          1061 => x"3f",
          1062 => x"a4",
          1063 => x"a4",
          1064 => x"0b",
          1065 => x"bc",
          1066 => x"08",
          1067 => x"05",
          1068 => x"08",
          1069 => x"08",
          1070 => x"08",
          1071 => x"82",
          1072 => x"08",
          1073 => x"08",
          1074 => x"88",
          1075 => x"82",
          1076 => x"0c",
          1077 => x"88",
          1078 => x"05",
          1079 => x"08",
          1080 => x"08",
          1081 => x"e0",
          1082 => x"33",
          1083 => x"81",
          1084 => x"0c",
          1085 => x"80",
          1086 => x"8c",
          1087 => x"08",
          1088 => x"8c",
          1089 => x"be",
          1090 => x"08",
          1091 => x"05",
          1092 => x"08",
          1093 => x"31",
          1094 => x"0c",
          1095 => x"08",
          1096 => x"82",
          1097 => x"08",
          1098 => x"0d",
          1099 => x"82",
          1100 => x"e0",
          1101 => x"80",
          1102 => x"05",
          1103 => x"90",
          1104 => x"05",
          1105 => x"90",
          1106 => x"05",
          1107 => x"a4",
          1108 => x"e0",
          1109 => x"71",
          1110 => x"05",
          1111 => x"fc",
          1112 => x"a4",
          1113 => x"98",
          1114 => x"a4",
          1115 => x"82",
          1116 => x"e0",
          1117 => x"e0",
          1118 => x"3f",
          1119 => x"98",
          1120 => x"a4",
          1121 => x"82",
          1122 => x"0b",
          1123 => x"82",
          1124 => x"2e",
          1125 => x"05",
          1126 => x"98",
          1127 => x"05",
          1128 => x"08",
          1129 => x"e4",
          1130 => x"05",
          1131 => x"a4",
          1132 => x"3f",
          1133 => x"08",
          1134 => x"a4",
          1135 => x"82",
          1136 => x"e0",
          1137 => x"e0",
          1138 => x"a4",
          1139 => x"08",
          1140 => x"fc",
          1141 => x"e0",
          1142 => x"38",
          1143 => x"05",
          1144 => x"08",
          1145 => x"82",
          1146 => x"09",
          1147 => x"08",
          1148 => x"08",
          1149 => x"82",
          1150 => x"05",
          1151 => x"82",
          1152 => x"e0",
          1153 => x"e0",
          1154 => x"a4",
          1155 => x"08",
          1156 => x"08",
          1157 => x"a4",
          1158 => x"82",
          1159 => x"e0",
          1160 => x"81",
          1161 => x"05",
          1162 => x"05",
          1163 => x"88",
          1164 => x"82",
          1165 => x"e0",
          1166 => x"82",
          1167 => x"82",
          1168 => x"e0",
          1169 => x"a4",
          1170 => x"82",
          1171 => x"05",
          1172 => x"ec",
          1173 => x"05",
          1174 => x"f0",
          1175 => x"05",
          1176 => x"08",
          1177 => x"08",
          1178 => x"05",
          1179 => x"08",
          1180 => x"05",
          1181 => x"53",
          1182 => x"08",
          1183 => x"a4",
          1184 => x"a4",
          1185 => x"08",
          1186 => x"08",
          1187 => x"a4",
          1188 => x"0c",
          1189 => x"04",
          1190 => x"a4",
          1191 => x"08",
          1192 => x"fc",
          1193 => x"05",
          1194 => x"8c",
          1195 => x"f0",
          1196 => x"e0",
          1197 => x"a4",
          1198 => x"08",
          1199 => x"a4",
          1200 => x"a4",
          1201 => x"e0",
          1202 => x"a4",
          1203 => x"08",
          1204 => x"fc",
          1205 => x"51",
          1206 => x"a4",
          1207 => x"0b",
          1208 => x"82",
          1209 => x"e0",
          1210 => x"82",
          1211 => x"82",
          1212 => x"2a",
          1213 => x"82",
          1214 => x"e0",
          1215 => x"e0",
          1216 => x"a4",
          1217 => x"51",
          1218 => x"e0",
          1219 => x"80",
          1220 => x"0c",
          1221 => x"82",
          1222 => x"0b",
          1223 => x"31",
          1224 => x"71",
          1225 => x"0c",
          1226 => x"82",
          1227 => x"82",
          1228 => x"e0",
          1229 => x"51",
          1230 => x"e0",
          1231 => x"80",
          1232 => x"0c",
          1233 => x"82",
          1234 => x"0b",
          1235 => x"31",
          1236 => x"71",
          1237 => x"0c",
          1238 => x"82",
          1239 => x"82",
          1240 => x"0b",
          1241 => x"31",
          1242 => x"81",
          1243 => x"70",
          1244 => x"08",
          1245 => x"e0",
          1246 => x"51",
          1247 => x"e0",
          1248 => x"02",
          1249 => x"82",
          1250 => x"82",
          1251 => x"84",
          1252 => x"82",
          1253 => x"82",
          1254 => x"31",
          1255 => x"53",
          1256 => x"04",
          1257 => x"a4",
          1258 => x"08",
          1259 => x"08",
          1260 => x"e0",
          1261 => x"53",
          1262 => x"04",
          1263 => x"a4",
          1264 => x"e0",
          1265 => x"a4",
          1266 => x"38",
          1267 => x"51",
          1268 => x"70",
          1269 => x"52",
          1270 => x"05",
          1271 => x"0c",
          1272 => x"80",
          1273 => x"88",
          1274 => x"e0",
          1275 => x"05",
          1276 => x"e0",
          1277 => x"a4",
          1278 => x"08",
          1279 => x"08",
          1280 => x"e0",
          1281 => x"05",
          1282 => x"08",
          1283 => x"08",
          1284 => x"e0",
          1285 => x"e0",
          1286 => x"ba",
          1287 => x"08",
          1288 => x"08",
          1289 => x"8d",
          1290 => x"e8",
          1291 => x"a4",
          1292 => x"e0",
          1293 => x"a4",
          1294 => x"08",
          1295 => x"08",
          1296 => x"fc",
          1297 => x"05",
          1298 => x"05",
          1299 => x"88",
          1300 => x"a4",
          1301 => x"08",
          1302 => x"38",
          1303 => x"10",
          1304 => x"ff",
          1305 => x"08",
          1306 => x"a4",
          1307 => x"08",
          1308 => x"a4",
          1309 => x"a4",
          1310 => x"08",
          1311 => x"f4",
          1312 => x"a4",
          1313 => x"71",
          1314 => x"0c",
          1315 => x"81",
          1316 => x"0c",
          1317 => x"82",
          1318 => x"82",
          1319 => x"31",
          1320 => x"82",
          1321 => x"05",
          1322 => x"51",
          1323 => x"fe",
          1324 => x"05",
          1325 => x"05",
          1326 => x"05",
          1327 => x"0d",
          1328 => x"a4",
          1329 => x"3d",
          1330 => x"fc",
          1331 => x"05",
          1332 => x"08",
          1333 => x"0c",
          1334 => x"82",
          1335 => x"82",
          1336 => x"e0",
          1337 => x"a4",
          1338 => x"e0",
          1339 => x"e0",
          1340 => x"a4",
          1341 => x"08",
          1342 => x"a4",
          1343 => x"a4",
          1344 => x"08",
          1345 => x"f4",
          1346 => x"f8",
          1347 => x"05",
          1348 => x"05",
          1349 => x"82",
          1350 => x"08",
          1351 => x"a4",
          1352 => x"e0",
          1353 => x"0d",
          1354 => x"a4",
          1355 => x"3d",
          1356 => x"f0",
          1357 => x"05",
          1358 => x"a4",
          1359 => x"53",
          1360 => x"08",
          1361 => x"53",
          1362 => x"38",
          1363 => x"70",
          1364 => x"39",
          1365 => x"53",
          1366 => x"38",
          1367 => x"05",
          1368 => x"08",
          1369 => x"08",
          1370 => x"08",
          1371 => x"f8",
          1372 => x"81",
          1373 => x"08",
          1374 => x"71",
          1375 => x"82",
          1376 => x"e0",
          1377 => x"a4",
          1378 => x"08",
          1379 => x"38",
          1380 => x"80",
          1381 => x"90",
          1382 => x"34",
          1383 => x"70",
          1384 => x"51",
          1385 => x"f8",
          1386 => x"82",
          1387 => x"e0",
          1388 => x"81",
          1389 => x"72",
          1390 => x"34",
          1391 => x"f8",
          1392 => x"38",
          1393 => x"05",
          1394 => x"08",
          1395 => x"90",
          1396 => x"33",
          1397 => x"39",
          1398 => x"05",
          1399 => x"e0",
          1400 => x"82",
          1401 => x"af",
          1402 => x"08",
          1403 => x"83",
          1404 => x"a4",
          1405 => x"8a",
          1406 => x"34",
          1407 => x"05",
          1408 => x"33",
          1409 => x"82",
          1410 => x"80",
          1411 => x"a4",
          1412 => x"53",
          1413 => x"34",
          1414 => x"d0",
          1415 => x"08",
          1416 => x"f8",
          1417 => x"38",
          1418 => x"f9",
          1419 => x"08",
          1420 => x"f8",
          1421 => x"38",
          1422 => x"05",
          1423 => x"08",
          1424 => x"f4",
          1425 => x"8d",
          1426 => x"ec",
          1427 => x"a4",
          1428 => x"a4",
          1429 => x"a4",
          1430 => x"e0",
          1431 => x"a4",
          1432 => x"05",
          1433 => x"55",
          1434 => x"f8",
          1435 => x"a4",
          1436 => x"2e",
          1437 => x"05",
          1438 => x"05",
          1439 => x"08",
          1440 => x"71",
          1441 => x"08",
          1442 => x"ec",
          1443 => x"3d",
          1444 => x"e0",
          1445 => x"f7",
          1446 => x"08",
          1447 => x"8c",
          1448 => x"e0",
          1449 => x"51",
          1450 => x"a4",
          1451 => x"06",
          1452 => x"91",
          1453 => x"08",
          1454 => x"ce",
          1455 => x"33",
          1456 => x"a4",
          1457 => x"f0",
          1458 => x"05",
          1459 => x"70",
          1460 => x"a4",
          1461 => x"08",
          1462 => x"09",
          1463 => x"a4",
          1464 => x"05",
          1465 => x"33",
          1466 => x"82",
          1467 => x"e0",
          1468 => x"a4",
          1469 => x"b6",
          1470 => x"08",
          1471 => x"39",
          1472 => x"05",
          1473 => x"08",
          1474 => x"08",
          1475 => x"08",
          1476 => x"0b",
          1477 => x"82",
          1478 => x"08",
          1479 => x"53",
          1480 => x"05",
          1481 => x"08",
          1482 => x"8d",
          1483 => x"ec",
          1484 => x"a4",
          1485 => x"27",
          1486 => x"05",
          1487 => x"8d",
          1488 => x"ec",
          1489 => x"82",
          1490 => x"39",
          1491 => x"53",
          1492 => x"a4",
          1493 => x"26",
          1494 => x"e0",
          1495 => x"39",
          1496 => x"05",
          1497 => x"fc",
          1498 => x"05",
          1499 => x"38",
          1500 => x"53",
          1501 => x"e0",
          1502 => x"51",
          1503 => x"05",
          1504 => x"33",
          1505 => x"a4",
          1506 => x"08",
          1507 => x"ad",
          1508 => x"33",
          1509 => x"a4",
          1510 => x"08",
          1511 => x"8d",
          1512 => x"ec",
          1513 => x"a4",
          1514 => x"08",
          1515 => x"26",
          1516 => x"08",
          1517 => x"e0",
          1518 => x"e0",
          1519 => x"e0",
          1520 => x"82",
          1521 => x"e0",
          1522 => x"81",
          1523 => x"52",
          1524 => x"08",
          1525 => x"e0",
          1526 => x"80",
          1527 => x"fc",
          1528 => x"fc",
          1529 => x"05",
          1530 => x"08",
          1531 => x"a4",
          1532 => x"08",
          1533 => x"8b",
          1534 => x"f8",
          1535 => x"56",
          1536 => x"8c",
          1537 => x"33",
          1538 => x"73",
          1539 => x"81",
          1540 => x"90",
          1541 => x"52",
          1542 => x"08",
          1543 => x"76",
          1544 => x"e0",
          1545 => x"54",
          1546 => x"17",
          1547 => x"77",
          1548 => x"e0",
          1549 => x"a0",
          1550 => x"3d",
          1551 => x"8e",
          1552 => x"05",
          1553 => x"51",
          1554 => x"80",
          1555 => x"f2",
          1556 => x"39",
          1557 => x"82",
          1558 => x"be",
          1559 => x"d4",
          1560 => x"51",
          1561 => x"80",
          1562 => x"39",
          1563 => x"bf",
          1564 => x"51",
          1565 => x"39",
          1566 => x"c0",
          1567 => x"51",
          1568 => x"39",
          1569 => x"c1",
          1570 => x"0d",
          1571 => x"56",
          1572 => x"52",
          1573 => x"87",
          1574 => x"82",
          1575 => x"9a",
          1576 => x"53",
          1577 => x"b1",
          1578 => x"3d",
          1579 => x"05",
          1580 => x"70",
          1581 => x"59",
          1582 => x"38",
          1583 => x"ff",
          1584 => x"82",
          1585 => x"70",
          1586 => x"e0",
          1587 => x"b9",
          1588 => x"98",
          1589 => x"96",
          1590 => x"77",
          1591 => x"82",
          1592 => x"08",
          1593 => x"89",
          1594 => x"d7",
          1595 => x"9f",
          1596 => x"80",
          1597 => x"06",
          1598 => x"90",
          1599 => x"98",
          1600 => x"3f",
          1601 => x"96",
          1602 => x"02",
          1603 => x"ff",
          1604 => x"fe",
          1605 => x"38",
          1606 => x"2e",
          1607 => x"56",
          1608 => x"53",
          1609 => x"e0",
          1610 => x"77",
          1611 => x"04",
          1612 => x"8c",
          1613 => x"15",
          1614 => x"5e",
          1615 => x"e0",
          1616 => x"58",
          1617 => x"72",
          1618 => x"80",
          1619 => x"52",
          1620 => x"3f",
          1621 => x"3f",
          1622 => x"38",
          1623 => x"2e",
          1624 => x"53",
          1625 => x"52",
          1626 => x"3f",
          1627 => x"ae",
          1628 => x"39",
          1629 => x"38",
          1630 => x"ff",
          1631 => x"d8",
          1632 => x"55",
          1633 => x"27",
          1634 => x"e4",
          1635 => x"82",
          1636 => x"81",
          1637 => x"a0",
          1638 => x"82",
          1639 => x"80",
          1640 => x"74",
          1641 => x"72",
          1642 => x"53",
          1643 => x"75",
          1644 => x"53",
          1645 => x"fe",
          1646 => x"52",
          1647 => x"08",
          1648 => x"15",
          1649 => x"51",
          1650 => x"5c",
          1651 => x"e0",
          1652 => x"51",
          1653 => x"ac",
          1654 => x"e0",
          1655 => x"70",
          1656 => x"70",
          1657 => x"06",
          1658 => x"80",
          1659 => x"fd",
          1660 => x"26",
          1661 => x"e0",
          1662 => x"3d",
          1663 => x"51",
          1664 => x"82",
          1665 => x"82",
          1666 => x"82",
          1667 => x"82",
          1668 => x"51",
          1669 => x"84",
          1670 => x"04",
          1671 => x"08",
          1672 => x"bf",
          1673 => x"3f",
          1674 => x"2a",
          1675 => x"2e",
          1676 => x"82",
          1677 => x"51",
          1678 => x"81",
          1679 => x"38",
          1680 => x"dc",
          1681 => x"f7",
          1682 => x"51",
          1683 => x"51",
          1684 => x"99",
          1685 => x"72",
          1686 => x"71",
          1687 => x"c7",
          1688 => x"3f",
          1689 => x"2a",
          1690 => x"2e",
          1691 => x"82",
          1692 => x"51",
          1693 => x"81",
          1694 => x"38",
          1695 => x"a8",
          1696 => x"ff",
          1697 => x"51",
          1698 => x"51",
          1699 => x"99",
          1700 => x"72",
          1701 => x"71",
          1702 => x"cf",
          1703 => x"3f",
          1704 => x"3f",
          1705 => x"77",
          1706 => x"55",
          1707 => x"ec",
          1708 => x"54",
          1709 => x"8c",
          1710 => x"b6",
          1711 => x"82",
          1712 => x"71",
          1713 => x"82",
          1714 => x"9c",
          1715 => x"06",
          1716 => x"52",
          1717 => x"e0",
          1718 => x"e0",
          1719 => x"39",
          1720 => x"3f",
          1721 => x"34",
          1722 => x"73",
          1723 => x"82",
          1724 => x"aa",
          1725 => x"0c",
          1726 => x"80",
          1727 => x"a4",
          1728 => x"c8",
          1729 => x"ff",
          1730 => x"06",
          1731 => x"82",
          1732 => x"3f",
          1733 => x"51",
          1734 => x"08",
          1735 => x"51",
          1736 => x"82",
          1737 => x"97",
          1738 => x"79",
          1739 => x"84",
          1740 => x"98",
          1741 => x"59",
          1742 => x"78",
          1743 => x"2e",
          1744 => x"38",
          1745 => x"bc",
          1746 => x"78",
          1747 => x"80",
          1748 => x"2e",
          1749 => x"80",
          1750 => x"f9",
          1751 => x"88",
          1752 => x"a7",
          1753 => x"2e",
          1754 => x"8b",
          1755 => x"38",
          1756 => x"8a",
          1757 => x"ff",
          1758 => x"ec",
          1759 => x"2e",
          1760 => x"11",
          1761 => x"3f",
          1762 => x"af",
          1763 => x"ff",
          1764 => x"e0",
          1765 => x"08",
          1766 => x"db",
          1767 => x"27",
          1768 => x"70",
          1769 => x"f5",
          1770 => x"80",
          1771 => x"c6",
          1772 => x"fd",
          1773 => x"53",
          1774 => x"82",
          1775 => x"38",
          1776 => x"84",
          1777 => x"98",
          1778 => x"c4",
          1779 => x"5a",
          1780 => x"59",
          1781 => x"34",
          1782 => x"3d",
          1783 => x"51",
          1784 => x"80",
          1785 => x"fc",
          1786 => x"ce",
          1787 => x"fc",
          1788 => x"53",
          1789 => x"82",
          1790 => x"38",
          1791 => x"3f",
          1792 => x"62",
          1793 => x"78",
          1794 => x"54",
          1795 => x"94",
          1796 => x"63",
          1797 => x"51",
          1798 => x"3d",
          1799 => x"51",
          1800 => x"80",
          1801 => x"78",
          1802 => x"08",
          1803 => x"33",
          1804 => x"de",
          1805 => x"fe",
          1806 => x"82",
          1807 => x"de",
          1808 => x"38",
          1809 => x"82",
          1810 => x"88",
          1811 => x"39",
          1812 => x"45",
          1813 => x"84",
          1814 => x"98",
          1815 => x"33",
          1816 => x"de",
          1817 => x"de",
          1818 => x"38",
          1819 => x"82",
          1820 => x"88",
          1821 => x"39",
          1822 => x"2e",
          1823 => x"99",
          1824 => x"80",
          1825 => x"44",
          1826 => x"05",
          1827 => x"ff",
          1828 => x"e0",
          1829 => x"63",
          1830 => x"81",
          1831 => x"72",
          1832 => x"51",
          1833 => x"7a",
          1834 => x"c5",
          1835 => x"55",
          1836 => x"51",
          1837 => x"87",
          1838 => x"53",
          1839 => x"82",
          1840 => x"38",
          1841 => x"84",
          1842 => x"98",
          1843 => x"02",
          1844 => x"81",
          1845 => x"53",
          1846 => x"82",
          1847 => x"39",
          1848 => x"c8",
          1849 => x"f8",
          1850 => x"ff",
          1851 => x"59",
          1852 => x"79",
          1853 => x"11",
          1854 => x"3f",
          1855 => x"38",
          1856 => x"79",
          1857 => x"39",
          1858 => x"3f",
          1859 => x"11",
          1860 => x"3f",
          1861 => x"97",
          1862 => x"ff",
          1863 => x"e0",
          1864 => x"59",
          1865 => x"82",
          1866 => x"fe",
          1867 => x"df",
          1868 => x"38",
          1869 => x"52",
          1870 => x"3f",
          1871 => x"52",
          1872 => x"46",
          1873 => x"b7",
          1874 => x"82",
          1875 => x"f0",
          1876 => x"ad",
          1877 => x"93",
          1878 => x"22",
          1879 => x"42",
          1880 => x"ff",
          1881 => x"3d",
          1882 => x"51",
          1883 => x"80",
          1884 => x"f0",
          1885 => x"e5",
          1886 => x"a0",
          1887 => x"84",
          1888 => x"53",
          1889 => x"82",
          1890 => x"39",
          1891 => x"e4",
          1892 => x"f8",
          1893 => x"ff",
          1894 => x"59",
          1895 => x"79",
          1896 => x"11",
          1897 => x"3f",
          1898 => x"38",
          1899 => x"05",
          1900 => x"51",
          1901 => x"b5",
          1902 => x"05",
          1903 => x"08",
          1904 => x"82",
          1905 => x"64",
          1906 => x"11",
          1907 => x"3f",
          1908 => x"9f",
          1909 => x"ff",
          1910 => x"82",
          1911 => x"38",
          1912 => x"ac",
          1913 => x"39",
          1914 => x"3f",
          1915 => x"82",
          1916 => x"80",
          1917 => x"f4",
          1918 => x"80",
          1919 => x"79",
          1920 => x"08",
          1921 => x"82",
          1922 => x"b5",
          1923 => x"3f",
          1924 => x"5a",
          1925 => x"82",
          1926 => x"82",
          1927 => x"38",
          1928 => x"7a",
          1929 => x"8c",
          1930 => x"ad",
          1931 => x"56",
          1932 => x"53",
          1933 => x"b0",
          1934 => x"39",
          1935 => x"51",
          1936 => x"82",
          1937 => x"90",
          1938 => x"ff",
          1939 => x"80",
          1940 => x"ff",
          1941 => x"82",
          1942 => x"7c",
          1943 => x"0a",
          1944 => x"ff",
          1945 => x"e0",
          1946 => x"70",
          1947 => x"5b",
          1948 => x"83",
          1949 => x"78",
          1950 => x"81",
          1951 => x"38",
          1952 => x"59",
          1953 => x"81",
          1954 => x"ff",
          1955 => x"3f",
          1956 => x"ff",
          1957 => x"3d",
          1958 => x"87",
          1959 => x"87",
          1960 => x"3f",
          1961 => x"08",
          1962 => x"51",
          1963 => x"08",
          1964 => x"70",
          1965 => x"72",
          1966 => x"08",
          1967 => x"84",
          1968 => x"72",
          1969 => x"8c",
          1970 => x"0c",
          1971 => x"94",
          1972 => x"84",
          1973 => x"34",
          1974 => x"3d",
          1975 => x"82",
          1976 => x"93",
          1977 => x"b4",
          1978 => x"b4",
          1979 => x"d2",
          1980 => x"8c",
          1981 => x"70",
          1982 => x"72",
          1983 => x"51",
          1984 => x"38",
          1985 => x"51",
          1986 => x"38",
          1987 => x"73",
          1988 => x"84",
          1989 => x"52",
          1990 => x"54",
          1991 => x"38",
          1992 => x"33",
          1993 => x"81",
          1994 => x"ea",
          1995 => x"a0",
          1996 => x"54",
          1997 => x"25",
          1998 => x"2e",
          1999 => x"54",
          2000 => x"82",
          2001 => x"fc",
          2002 => x"2e",
          2003 => x"72",
          2004 => x"08",
          2005 => x"53",
          2006 => x"0d",
          2007 => x"33",
          2008 => x"8b",
          2009 => x"ff",
          2010 => x"81",
          2011 => x"52",
          2012 => x"13",
          2013 => x"80",
          2014 => x"52",
          2015 => x"13",
          2016 => x"26",
          2017 => x"87",
          2018 => x"38",
          2019 => x"72",
          2020 => x"13",
          2021 => x"13",
          2022 => x"13",
          2023 => x"13",
          2024 => x"13",
          2025 => x"87",
          2026 => x"98",
          2027 => x"9c",
          2028 => x"0c",
          2029 => x"7f",
          2030 => x"7d",
          2031 => x"7d",
          2032 => x"5a",
          2033 => x"b4",
          2034 => x"c0",
          2035 => x"34",
          2036 => x"85",
          2037 => x"5a",
          2038 => x"a4",
          2039 => x"c0",
          2040 => x"23",
          2041 => x"06",
          2042 => x"86",
          2043 => x"84",
          2044 => x"82",
          2045 => x"06",
          2046 => x"9b",
          2047 => x"0d",
          2048 => x"72",
          2049 => x"72",
          2050 => x"80",
          2051 => x"80",
          2052 => x"39",
          2053 => x"98",
          2054 => x"ff",
          2055 => x"54",
          2056 => x"38",
          2057 => x"70",
          2058 => x"70",
          2059 => x"0c",
          2060 => x"80",
          2061 => x"81",
          2062 => x"08",
          2063 => x"ff",
          2064 => x"e3",
          2065 => x"3d",
          2066 => x"05",
          2067 => x"ff",
          2068 => x"84",
          2069 => x"c0",
          2070 => x"2a",
          2071 => x"80",
          2072 => x"81",
          2073 => x"81",
          2074 => x"80",
          2075 => x"81",
          2076 => x"73",
          2077 => x"80",
          2078 => x"c0",
          2079 => x"82",
          2080 => x"ff",
          2081 => x"30",
          2082 => x"82",
          2083 => x"f9",
          2084 => x"77",
          2085 => x"7a",
          2086 => x"b0",
          2087 => x"87",
          2088 => x"86",
          2089 => x"08",
          2090 => x"56",
          2091 => x"91",
          2092 => x"d7",
          2093 => x"51",
          2094 => x"93",
          2095 => x"ff",
          2096 => x"87",
          2097 => x"86",
          2098 => x"74",
          2099 => x"89",
          2100 => x"54",
          2101 => x"53",
          2102 => x"38",
          2103 => x"de",
          2104 => x"57",
          2105 => x"75",
          2106 => x"94",
          2107 => x"81",
          2108 => x"8c",
          2109 => x"51",
          2110 => x"70",
          2111 => x"8d",
          2112 => x"51",
          2113 => x"ff",
          2114 => x"70",
          2115 => x"90",
          2116 => x"33",
          2117 => x"70",
          2118 => x"0c",
          2119 => x"82",
          2120 => x"54",
          2121 => x"80",
          2122 => x"51",
          2123 => x"06",
          2124 => x"38",
          2125 => x"94",
          2126 => x"87",
          2127 => x"81",
          2128 => x"84",
          2129 => x"e0",
          2130 => x"98",
          2131 => x"b0",
          2132 => x"87",
          2133 => x"86",
          2134 => x"08",
          2135 => x"51",
          2136 => x"38",
          2137 => x"94",
          2138 => x"87",
          2139 => x"98",
          2140 => x"71",
          2141 => x"04",
          2142 => x"08",
          2143 => x"70",
          2144 => x"9e",
          2145 => x"c0",
          2146 => x"87",
          2147 => x"0c",
          2148 => x"c0",
          2149 => x"de",
          2150 => x"82",
          2151 => x"08",
          2152 => x"b0",
          2153 => x"9e",
          2154 => x"c0",
          2155 => x"87",
          2156 => x"0c",
          2157 => x"e0",
          2158 => x"de",
          2159 => x"51",
          2160 => x"9e",
          2161 => x"c0",
          2162 => x"87",
          2163 => x"0c",
          2164 => x"0b",
          2165 => x"80",
          2166 => x"2e",
          2167 => x"f9",
          2168 => x"08",
          2169 => x"52",
          2170 => x"71",
          2171 => x"c0",
          2172 => x"06",
          2173 => x"38",
          2174 => x"80",
          2175 => x"88",
          2176 => x"80",
          2177 => x"de",
          2178 => x"90",
          2179 => x"52",
          2180 => x"52",
          2181 => x"87",
          2182 => x"80",
          2183 => x"83",
          2184 => x"34",
          2185 => x"70",
          2186 => x"70",
          2187 => x"82",
          2188 => x"9e",
          2189 => x"51",
          2190 => x"81",
          2191 => x"0b",
          2192 => x"80",
          2193 => x"2e",
          2194 => x"81",
          2195 => x"08",
          2196 => x"52",
          2197 => x"71",
          2198 => x"c0",
          2199 => x"51",
          2200 => x"81",
          2201 => x"c0",
          2202 => x"70",
          2203 => x"df",
          2204 => x"90",
          2205 => x"52",
          2206 => x"71",
          2207 => x"90",
          2208 => x"2a",
          2209 => x"34",
          2210 => x"70",
          2211 => x"2e",
          2212 => x"87",
          2213 => x"87",
          2214 => x"34",
          2215 => x"82",
          2216 => x"82",
          2217 => x"89",
          2218 => x"bb",
          2219 => x"be",
          2220 => x"80",
          2221 => x"82",
          2222 => x"c8",
          2223 => x"de",
          2224 => x"38",
          2225 => x"08",
          2226 => x"ff",
          2227 => x"54",
          2228 => x"b4",
          2229 => x"52",
          2230 => x"3f",
          2231 => x"2e",
          2232 => x"de",
          2233 => x"b0",
          2234 => x"fe",
          2235 => x"82",
          2236 => x"11",
          2237 => x"88",
          2238 => x"73",
          2239 => x"33",
          2240 => x"8b",
          2241 => x"80",
          2242 => x"52",
          2243 => x"3f",
          2244 => x"2e",
          2245 => x"82",
          2246 => x"82",
          2247 => x"89",
          2248 => x"d6",
          2249 => x"80",
          2250 => x"ff",
          2251 => x"54",
          2252 => x"e8",
          2253 => x"81",
          2254 => x"82",
          2255 => x"82",
          2256 => x"89",
          2257 => x"8e",
          2258 => x"86",
          2259 => x"cb",
          2260 => x"de",
          2261 => x"ff",
          2262 => x"52",
          2263 => x"3f",
          2264 => x"3f",
          2265 => x"90",
          2266 => x"ec",
          2267 => x"51",
          2268 => x"08",
          2269 => x"54",
          2270 => x"cc",
          2271 => x"de",
          2272 => x"38",
          2273 => x"c0",
          2274 => x"82",
          2275 => x"76",
          2276 => x"08",
          2277 => x"e3",
          2278 => x"80",
          2279 => x"56",
          2280 => x"b7",
          2281 => x"84",
          2282 => x"82",
          2283 => x"51",
          2284 => x"a4",
          2285 => x"3d",
          2286 => x"52",
          2287 => x"29",
          2288 => x"04",
          2289 => x"cd",
          2290 => x"51",
          2291 => x"39",
          2292 => x"cd",
          2293 => x"3d",
          2294 => x"80",
          2295 => x"82",
          2296 => x"0c",
          2297 => x"70",
          2298 => x"2c",
          2299 => x"53",
          2300 => x"cd",
          2301 => x"25",
          2302 => x"12",
          2303 => x"33",
          2304 => x"81",
          2305 => x"e0",
          2306 => x"3d",
          2307 => x"33",
          2308 => x"2e",
          2309 => x"88",
          2310 => x"fc",
          2311 => x"3f",
          2312 => x"ff",
          2313 => x"53",
          2314 => x"53",
          2315 => x"3f",
          2316 => x"f6",
          2317 => x"05",
          2318 => x"82",
          2319 => x"df",
          2320 => x"5a",
          2321 => x"74",
          2322 => x"33",
          2323 => x"81",
          2324 => x"fe",
          2325 => x"82",
          2326 => x"df",
          2327 => x"74",
          2328 => x"52",
          2329 => x"df",
          2330 => x"df",
          2331 => x"93",
          2332 => x"df",
          2333 => x"82",
          2334 => x"ac",
          2335 => x"a4",
          2336 => x"53",
          2337 => x"3f",
          2338 => x"81",
          2339 => x"51",
          2340 => x"04",
          2341 => x"93",
          2342 => x"89",
          2343 => x"73",
          2344 => x"73",
          2345 => x"df",
          2346 => x"71",
          2347 => x"f0",
          2348 => x"99",
          2349 => x"0c",
          2350 => x"81",
          2351 => x"51",
          2352 => x"08",
          2353 => x"53",
          2354 => x"56",
          2355 => x"08",
          2356 => x"a9",
          2357 => x"80",
          2358 => x"38",
          2359 => x"17",
          2360 => x"76",
          2361 => x"57",
          2362 => x"09",
          2363 => x"0d",
          2364 => x"ad",
          2365 => x"58",
          2366 => x"80",
          2367 => x"81",
          2368 => x"08",
          2369 => x"70",
          2370 => x"e0",
          2371 => x"51",
          2372 => x"08",
          2373 => x"e0",
          2374 => x"98",
          2375 => x"80",
          2376 => x"72",
          2377 => x"77",
          2378 => x"82",
          2379 => x"51",
          2380 => x"08",
          2381 => x"51",
          2382 => x"09",
          2383 => x"51",
          2384 => x"a7",
          2385 => x"e0",
          2386 => x"82",
          2387 => x"f6",
          2388 => x"72",
          2389 => x"2e",
          2390 => x"78",
          2391 => x"81",
          2392 => x"58",
          2393 => x"86",
          2394 => x"54",
          2395 => x"70",
          2396 => x"82",
          2397 => x"08",
          2398 => x"98",
          2399 => x"55",
          2400 => x"2e",
          2401 => x"ac",
          2402 => x"11",
          2403 => x"82",
          2404 => x"ff",
          2405 => x"b1",
          2406 => x"06",
          2407 => x"39",
          2408 => x"54",
          2409 => x"54",
          2410 => x"0d",
          2411 => x"b2",
          2412 => x"5a",
          2413 => x"e8",
          2414 => x"73",
          2415 => x"33",
          2416 => x"76",
          2417 => x"76",
          2418 => x"ad",
          2419 => x"e0",
          2420 => x"e0",
          2421 => x"93",
          2422 => x"51",
          2423 => x"08",
          2424 => x"51",
          2425 => x"82",
          2426 => x"08",
          2427 => x"52",
          2428 => x"98",
          2429 => x"2e",
          2430 => x"e0",
          2431 => x"82",
          2432 => x"e0",
          2433 => x"98",
          2434 => x"80",
          2435 => x"06",
          2436 => x"1b",
          2437 => x"7b",
          2438 => x"2e",
          2439 => x"39",
          2440 => x"38",
          2441 => x"38",
          2442 => x"51",
          2443 => x"98",
          2444 => x"ff",
          2445 => x"82",
          2446 => x"98",
          2447 => x"2b",
          2448 => x"70",
          2449 => x"08",
          2450 => x"59",
          2451 => x"73",
          2452 => x"27",
          2453 => x"81",
          2454 => x"55",
          2455 => x"53",
          2456 => x"82",
          2457 => x"73",
          2458 => x"d0",
          2459 => x"80",
          2460 => x"98",
          2461 => x"55",
          2462 => x"74",
          2463 => x"e0",
          2464 => x"cc",
          2465 => x"2e",
          2466 => x"82",
          2467 => x"98",
          2468 => x"2b",
          2469 => x"82",
          2470 => x"51",
          2471 => x"77",
          2472 => x"82",
          2473 => x"0b",
          2474 => x"f7",
          2475 => x"d4",
          2476 => x"af",
          2477 => x"73",
          2478 => x"29",
          2479 => x"04",
          2480 => x"2e",
          2481 => x"55",
          2482 => x"2b",
          2483 => x"24",
          2484 => x"81",
          2485 => x"81",
          2486 => x"f7",
          2487 => x"82",
          2488 => x"74",
          2489 => x"ae",
          2490 => x"33",
          2491 => x"14",
          2492 => x"f7",
          2493 => x"81",
          2494 => x"f7",
          2495 => x"77",
          2496 => x"52",
          2497 => x"97",
          2498 => x"81",
          2499 => x"f7",
          2500 => x"24",
          2501 => x"98",
          2502 => x"33",
          2503 => x"fc",
          2504 => x"88",
          2505 => x"80",
          2506 => x"98",
          2507 => x"55",
          2508 => x"39",
          2509 => x"34",
          2510 => x"c1",
          2511 => x"39",
          2512 => x"06",
          2513 => x"38",
          2514 => x"73",
          2515 => x"73",
          2516 => x"08",
          2517 => x"82",
          2518 => x"98",
          2519 => x"56",
          2520 => x"1a",
          2521 => x"fb",
          2522 => x"96",
          2523 => x"81",
          2524 => x"f7",
          2525 => x"24",
          2526 => x"a0",
          2527 => x"dc",
          2528 => x"82",
          2529 => x"74",
          2530 => x"fc",
          2531 => x"3f",
          2532 => x"0a",
          2533 => x"33",
          2534 => x"38",
          2535 => x"7a",
          2536 => x"fc",
          2537 => x"3f",
          2538 => x"c7",
          2539 => x"06",
          2540 => x"33",
          2541 => x"53",
          2542 => x"84",
          2543 => x"f7",
          2544 => x"34",
          2545 => x"0d",
          2546 => x"80",
          2547 => x"08",
          2548 => x"82",
          2549 => x"82",
          2550 => x"54",
          2551 => x"f7",
          2552 => x"f9",
          2553 => x"f7",
          2554 => x"2c",
          2555 => x"74",
          2556 => x"81",
          2557 => x"08",
          2558 => x"3f",
          2559 => x"0a",
          2560 => x"33",
          2561 => x"38",
          2562 => x"ff",
          2563 => x"70",
          2564 => x"d8",
          2565 => x"24",
          2566 => x"52",
          2567 => x"81",
          2568 => x"70",
          2569 => x"51",
          2570 => x"fb",
          2571 => x"ff",
          2572 => x"54",
          2573 => x"fb",
          2574 => x"82",
          2575 => x"52",
          2576 => x"dc",
          2577 => x"d8",
          2578 => x"d6",
          2579 => x"53",
          2580 => x"ee",
          2581 => x"80",
          2582 => x"39",
          2583 => x"55",
          2584 => x"ff",
          2585 => x"82",
          2586 => x"81",
          2587 => x"79",
          2588 => x"81",
          2589 => x"90",
          2590 => x"80",
          2591 => x"c0",
          2592 => x"d8",
          2593 => x"06",
          2594 => x"ff",
          2595 => x"fa",
          2596 => x"f6",
          2597 => x"3f",
          2598 => x"06",
          2599 => x"74",
          2600 => x"99",
          2601 => x"f7",
          2602 => x"ff",
          2603 => x"51",
          2604 => x"7a",
          2605 => x"08",
          2606 => x"74",
          2607 => x"98",
          2608 => x"98",
          2609 => x"74",
          2610 => x"81",
          2611 => x"89",
          2612 => x"7a",
          2613 => x"d8",
          2614 => x"f5",
          2615 => x"81",
          2616 => x"56",
          2617 => x"82",
          2618 => x"73",
          2619 => x"33",
          2620 => x"eb",
          2621 => x"80",
          2622 => x"08",
          2623 => x"82",
          2624 => x"82",
          2625 => x"3d",
          2626 => x"88",
          2627 => x"23",
          2628 => x"fa",
          2629 => x"e0",
          2630 => x"34",
          2631 => x"e0",
          2632 => x"76",
          2633 => x"54",
          2634 => x"34",
          2635 => x"22",
          2636 => x"83",
          2637 => x"51",
          2638 => x"89",
          2639 => x"88",
          2640 => x"11",
          2641 => x"76",
          2642 => x"ff",
          2643 => x"72",
          2644 => x"82",
          2645 => x"51",
          2646 => x"3d",
          2647 => x"05",
          2648 => x"71",
          2649 => x"2b",
          2650 => x"70",
          2651 => x"07",
          2652 => x"81",
          2653 => x"53",
          2654 => x"53",
          2655 => x"18",
          2656 => x"88",
          2657 => x"74",
          2658 => x"70",
          2659 => x"88",
          2660 => x"f8",
          2661 => x"73",
          2662 => x"54",
          2663 => x"81",
          2664 => x"82",
          2665 => x"34",
          2666 => x"04",
          2667 => x"02",
          2668 => x"2b",
          2669 => x"33",
          2670 => x"58",
          2671 => x"84",
          2672 => x"2b",
          2673 => x"52",
          2674 => x"34",
          2675 => x"11",
          2676 => x"71",
          2677 => x"72",
          2678 => x"71",
          2679 => x"56",
          2680 => x"87",
          2681 => x"70",
          2682 => x"07",
          2683 => x"2a",
          2684 => x"34",
          2685 => x"04",
          2686 => x"82",
          2687 => x"11",
          2688 => x"2b",
          2689 => x"81",
          2690 => x"2b",
          2691 => x"56",
          2692 => x"f6",
          2693 => x"e0",
          2694 => x"12",
          2695 => x"07",
          2696 => x"71",
          2697 => x"ff",
          2698 => x"5a",
          2699 => x"54",
          2700 => x"13",
          2701 => x"70",
          2702 => x"71",
          2703 => x"72",
          2704 => x"88",
          2705 => x"70",
          2706 => x"72",
          2707 => x"3d",
          2708 => x"88",
          2709 => x"70",
          2710 => x"83",
          2711 => x"2b",
          2712 => x"73",
          2713 => x"88",
          2714 => x"22",
          2715 => x"53",
          2716 => x"14",
          2717 => x"70",
          2718 => x"71",
          2719 => x"72",
          2720 => x"71",
          2721 => x"55",
          2722 => x"83",
          2723 => x"82",
          2724 => x"2b",
          2725 => x"87",
          2726 => x"82",
          2727 => x"83",
          2728 => x"fd",
          2729 => x"83",
          2730 => x"12",
          2731 => x"07",
          2732 => x"71",
          2733 => x"42",
          2734 => x"54",
          2735 => x"80",
          2736 => x"84",
          2737 => x"71",
          2738 => x"11",
          2739 => x"55",
          2740 => x"06",
          2741 => x"88",
          2742 => x"13",
          2743 => x"2a",
          2744 => x"16",
          2745 => x"88",
          2746 => x"34",
          2747 => x"88",
          2748 => x"85",
          2749 => x"70",
          2750 => x"07",
          2751 => x"2a",
          2752 => x"34",
          2753 => x"04",
          2754 => x"88",
          2755 => x"80",
          2756 => x"3f",
          2757 => x"80",
          2758 => x"e0",
          2759 => x"e0",
          2760 => x"33",
          2761 => x"56",
          2762 => x"78",
          2763 => x"17",
          2764 => x"2b",
          2765 => x"31",
          2766 => x"27",
          2767 => x"79",
          2768 => x"38",
          2769 => x"85",
          2770 => x"54",
          2771 => x"2e",
          2772 => x"76",
          2773 => x"70",
          2774 => x"07",
          2775 => x"5a",
          2776 => x"38",
          2777 => x"81",
          2778 => x"81",
          2779 => x"06",
          2780 => x"81",
          2781 => x"52",
          2782 => x"88",
          2783 => x"12",
          2784 => x"07",
          2785 => x"17",
          2786 => x"2a",
          2787 => x"34",
          2788 => x"15",
          2789 => x"2b",
          2790 => x"87",
          2791 => x"88",
          2792 => x"54",
          2793 => x"34",
          2794 => x"11",
          2795 => x"71",
          2796 => x"74",
          2797 => x"87",
          2798 => x"16",
          2799 => x"33",
          2800 => x"53",
          2801 => x"16",
          2802 => x"88",
          2803 => x"e0",
          2804 => x"3d",
          2805 => x"84",
          2806 => x"80",
          2807 => x"3f",
          2808 => x"e0",
          2809 => x"3d",
          2810 => x"42",
          2811 => x"09",
          2812 => x"7b",
          2813 => x"82",
          2814 => x"7e",
          2815 => x"7e",
          2816 => x"8f",
          2817 => x"ff",
          2818 => x"31",
          2819 => x"70",
          2820 => x"12",
          2821 => x"31",
          2822 => x"29",
          2823 => x"33",
          2824 => x"70",
          2825 => x"41",
          2826 => x"5b",
          2827 => x"81",
          2828 => x"ff",
          2829 => x"83",
          2830 => x"88",
          2831 => x"71",
          2832 => x"47",
          2833 => x"8b",
          2834 => x"ff",
          2835 => x"fe",
          2836 => x"09",
          2837 => x"c0",
          2838 => x"81",
          2839 => x"24",
          2840 => x"81",
          2841 => x"24",
          2842 => x"33",
          2843 => x"53",
          2844 => x"78",
          2845 => x"08",
          2846 => x"53",
          2847 => x"11",
          2848 => x"ce",
          2849 => x"05",
          2850 => x"81",
          2851 => x"24",
          2852 => x"3f",
          2853 => x"33",
          2854 => x"53",
          2855 => x"78",
          2856 => x"08",
          2857 => x"53",
          2858 => x"11",
          2859 => x"f6",
          2860 => x"05",
          2861 => x"83",
          2862 => x"7f",
          2863 => x"98",
          2864 => x"2e",
          2865 => x"e0",
          2866 => x"73",
          2867 => x"78",
          2868 => x"78",
          2869 => x"2b",
          2870 => x"51",
          2871 => x"e0",
          2872 => x"3d",
          2873 => x"fb",
          2874 => x"82",
          2875 => x"73",
          2876 => x"51",
          2877 => x"98",
          2878 => x"0d",
          2879 => x"70",
          2880 => x"11",
          2881 => x"83",
          2882 => x"9b",
          2883 => x"33",
          2884 => x"80",
          2885 => x"92",
          2886 => x"80",
          2887 => x"72",
          2888 => x"81",
          2889 => x"8c",
          2890 => x"06",
          2891 => x"87",
          2892 => x"38",
          2893 => x"71",
          2894 => x"51",
          2895 => x"e0",
          2896 => x"33",
          2897 => x"3d",
          2898 => x"64",
          2899 => x"40",
          2900 => x"cd",
          2901 => x"7a",
          2902 => x"72",
          2903 => x"11",
          2904 => x"92",
          2905 => x"58",
          2906 => x"76",
          2907 => x"70",
          2908 => x"54",
          2909 => x"52",
          2910 => x"81",
          2911 => x"53",
          2912 => x"78",
          2913 => x"2e",
          2914 => x"52",
          2915 => x"08",
          2916 => x"84",
          2917 => x"87",
          2918 => x"70",
          2919 => x"ff",
          2920 => x"81",
          2921 => x"57",
          2922 => x"80",
          2923 => x"78",
          2924 => x"80",
          2925 => x"81",
          2926 => x"0c",
          2927 => x"60",
          2928 => x"33",
          2929 => x"74",
          2930 => x"98",
          2931 => x"78",
          2932 => x"77",
          2933 => x"11",
          2934 => x"92",
          2935 => x"85",
          2936 => x"7d",
          2937 => x"08",
          2938 => x"53",
          2939 => x"70",
          2940 => x"18",
          2941 => x"51",
          2942 => x"c0",
          2943 => x"87",
          2944 => x"2e",
          2945 => x"38",
          2946 => x"15",
          2947 => x"52",
          2948 => x"39",
          2949 => x"80",
          2950 => x"90",
          2951 => x"71",
          2952 => x"38",
          2953 => x"80",
          2954 => x"72",
          2955 => x"04",
          2956 => x"a3",
          2957 => x"33",
          2958 => x"3f",
          2959 => x"83",
          2960 => x"87",
          2961 => x"76",
          2962 => x"93",
          2963 => x"8c",
          2964 => x"38",
          2965 => x"c6",
          2966 => x"81",
          2967 => x"71",
          2968 => x"8c",
          2969 => x"98",
          2970 => x"73",
          2971 => x"72",
          2972 => x"f7",
          2973 => x"88",
          2974 => x"80",
          2975 => x"56",
          2976 => x"88",
          2977 => x"81",
          2978 => x"07",
          2979 => x"3d",
          2980 => x"11",
          2981 => x"71",
          2982 => x"72",
          2983 => x"82",
          2984 => x"54",
          2985 => x"0d",
          2986 => x"52",
          2987 => x"34",
          2988 => x"83",
          2989 => x"75",
          2990 => x"54",
          2991 => x"70",
          2992 => x"51",
          2993 => x"70",
          2994 => x"3d",
          2995 => x"77",
          2996 => x"38",
          2997 => x"70",
          2998 => x"eb",
          2999 => x"0d",
          3000 => x"72",
          3001 => x"51",
          3002 => x"fc",
          3003 => x"53",
          3004 => x"70",
          3005 => x"ff",
          3006 => x"2e",
          3007 => x"71",
          3008 => x"04",
          3009 => x"89",
          3010 => x"11",
          3011 => x"70",
          3012 => x"0d",
          3013 => x"04",
          3014 => x"70",
          3015 => x"55",
          3016 => x"98",
          3017 => x"38",
          3018 => x"a2",
          3019 => x"ff",
          3020 => x"73",
          3021 => x"98",
          3022 => x"0d",
          3023 => x"56",
          3024 => x"81",
          3025 => x"70",
          3026 => x"e4",
          3027 => x"09",
          3028 => x"08",
          3029 => x"a8",
          3030 => x"56",
          3031 => x"16",
          3032 => x"06",
          3033 => x"78",
          3034 => x"3f",
          3035 => x"98",
          3036 => x"0d",
          3037 => x"b4",
          3038 => x"fe",
          3039 => x"82",
          3040 => x"74",
          3041 => x"51",
          3042 => x"80",
          3043 => x"74",
          3044 => x"0c",
          3045 => x"7a",
          3046 => x"e0",
          3047 => x"81",
          3048 => x"2e",
          3049 => x"17",
          3050 => x"06",
          3051 => x"e0",
          3052 => x"56",
          3053 => x"84",
          3054 => x"8b",
          3055 => x"eb",
          3056 => x"84",
          3057 => x"17",
          3058 => x"d3",
          3059 => x"17",
          3060 => x"81",
          3061 => x"53",
          3062 => x"c4",
          3063 => x"80",
          3064 => x"3f",
          3065 => x"38",
          3066 => x"8a",
          3067 => x"fe",
          3068 => x"56",
          3069 => x"38",
          3070 => x"16",
          3071 => x"98",
          3072 => x"0d",
          3073 => x"81",
          3074 => x"15",
          3075 => x"33",
          3076 => x"38",
          3077 => x"2e",
          3078 => x"2e",
          3079 => x"81",
          3080 => x"08",
          3081 => x"3f",
          3082 => x"74",
          3083 => x"81",
          3084 => x"05",
          3085 => x"f5",
          3086 => x"38",
          3087 => x"33",
          3088 => x"06",
          3089 => x"53",
          3090 => x"06",
          3091 => x"a8",
          3092 => x"bd",
          3093 => x"38",
          3094 => x"b8",
          3095 => x"98",
          3096 => x"39",
          3097 => x"52",
          3098 => x"98",
          3099 => x"fc",
          3100 => x"ba",
          3101 => x"06",
          3102 => x"e0",
          3103 => x"3d",
          3104 => x"82",
          3105 => x"76",
          3106 => x"75",
          3107 => x"38",
          3108 => x"2e",
          3109 => x"2e",
          3110 => x"81",
          3111 => x"08",
          3112 => x"3f",
          3113 => x"98",
          3114 => x"06",
          3115 => x"06",
          3116 => x"2e",
          3117 => x"06",
          3118 => x"53",
          3119 => x"34",
          3120 => x"52",
          3121 => x"98",
          3122 => x"94",
          3123 => x"05",
          3124 => x"38",
          3125 => x"06",
          3126 => x"74",
          3127 => x"a8",
          3128 => x"9d",
          3129 => x"e0",
          3130 => x"ff",
          3131 => x"06",
          3132 => x"3f",
          3133 => x"08",
          3134 => x"82",
          3135 => x"08",
          3136 => x"82",
          3137 => x"05",
          3138 => x"3f",
          3139 => x"74",
          3140 => x"81",
          3141 => x"98",
          3142 => x"0d",
          3143 => x"56",
          3144 => x"9c",
          3145 => x"2e",
          3146 => x"51",
          3147 => x"54",
          3148 => x"93",
          3149 => x"54",
          3150 => x"54",
          3151 => x"fb",
          3152 => x"82",
          3153 => x"38",
          3154 => x"38",
          3155 => x"38",
          3156 => x"d6",
          3157 => x"9c",
          3158 => x"57",
          3159 => x"81",
          3160 => x"81",
          3161 => x"55",
          3162 => x"54",
          3163 => x"0d",
          3164 => x"08",
          3165 => x"17",
          3166 => x"9c",
          3167 => x"58",
          3168 => x"fd",
          3169 => x"08",
          3170 => x"08",
          3171 => x"82",
          3172 => x"98",
          3173 => x"94",
          3174 => x"2e",
          3175 => x"81",
          3176 => x"9c",
          3177 => x"56",
          3178 => x"80",
          3179 => x"09",
          3180 => x"08",
          3181 => x"30",
          3182 => x"07",
          3183 => x"55",
          3184 => x"98",
          3185 => x"08",
          3186 => x"9c",
          3187 => x"85",
          3188 => x"81",
          3189 => x"89",
          3190 => x"ac",
          3191 => x"3f",
          3192 => x"38",
          3193 => x"2e",
          3194 => x"98",
          3195 => x"70",
          3196 => x"7c",
          3197 => x"f8",
          3198 => x"ff",
          3199 => x"ff",
          3200 => x"3f",
          3201 => x"08",
          3202 => x"80",
          3203 => x"94",
          3204 => x"53",
          3205 => x"82",
          3206 => x"75",
          3207 => x"05",
          3208 => x"26",
          3209 => x"84",
          3210 => x"18",
          3211 => x"2e",
          3212 => x"39",
          3213 => x"81",
          3214 => x"0c",
          3215 => x"7a",
          3216 => x"e0",
          3217 => x"98",
          3218 => x"51",
          3219 => x"82",
          3220 => x"84",
          3221 => x"52",
          3222 => x"39",
          3223 => x"75",
          3224 => x"19",
          3225 => x"ed",
          3226 => x"2e",
          3227 => x"70",
          3228 => x"53",
          3229 => x"0c",
          3230 => x"7a",
          3231 => x"f0",
          3232 => x"9f",
          3233 => x"90",
          3234 => x"aa",
          3235 => x"88",
          3236 => x"38",
          3237 => x"17",
          3238 => x"fe",
          3239 => x"80",
          3240 => x"2b",
          3241 => x"73",
          3242 => x"e0",
          3243 => x"ff",
          3244 => x"98",
          3245 => x"82",
          3246 => x"58",
          3247 => x"39",
          3248 => x"82",
          3249 => x"94",
          3250 => x"58",
          3251 => x"81",
          3252 => x"98",
          3253 => x"b8",
          3254 => x"82",
          3255 => x"f8",
          3256 => x"08",
          3257 => x"0a",
          3258 => x"15",
          3259 => x"72",
          3260 => x"ff",
          3261 => x"13",
          3262 => x"74",
          3263 => x"22",
          3264 => x"38",
          3265 => x"05",
          3266 => x"8a",
          3267 => x"3f",
          3268 => x"81",
          3269 => x"ff",
          3270 => x"ff",
          3271 => x"82",
          3272 => x"7b",
          3273 => x"55",
          3274 => x"73",
          3275 => x"08",
          3276 => x"80",
          3277 => x"e0",
          3278 => x"55",
          3279 => x"38",
          3280 => x"fb",
          3281 => x"38",
          3282 => x"51",
          3283 => x"98",
          3284 => x"16",
          3285 => x"74",
          3286 => x"04",
          3287 => x"5b",
          3288 => x"ac",
          3289 => x"e0",
          3290 => x"98",
          3291 => x"51",
          3292 => x"54",
          3293 => x"82",
          3294 => x"33",
          3295 => x"09",
          3296 => x"e0",
          3297 => x"55",
          3298 => x"8e",
          3299 => x"09",
          3300 => x"e0",
          3301 => x"fd",
          3302 => x"82",
          3303 => x"38",
          3304 => x"38",
          3305 => x"8b",
          3306 => x"9a",
          3307 => x"e0",
          3308 => x"70",
          3309 => x"09",
          3310 => x"eb",
          3311 => x"2b",
          3312 => x"0c",
          3313 => x"77",
          3314 => x"9a",
          3315 => x"76",
          3316 => x"09",
          3317 => x"52",
          3318 => x"3d",
          3319 => x"80",
          3320 => x"81",
          3321 => x"56",
          3322 => x"ff",
          3323 => x"38",
          3324 => x"0d",
          3325 => x"59",
          3326 => x"70",
          3327 => x"83",
          3328 => x"51",
          3329 => x"5b",
          3330 => x"9c",
          3331 => x"86",
          3332 => x"15",
          3333 => x"58",
          3334 => x"98",
          3335 => x"81",
          3336 => x"98",
          3337 => x"06",
          3338 => x"53",
          3339 => x"77",
          3340 => x"09",
          3341 => x"7f",
          3342 => x"ef",
          3343 => x"81",
          3344 => x"06",
          3345 => x"8d",
          3346 => x"90",
          3347 => x"5d",
          3348 => x"9c",
          3349 => x"2e",
          3350 => x"1e",
          3351 => x"3f",
          3352 => x"06",
          3353 => x"70",
          3354 => x"51",
          3355 => x"a8",
          3356 => x"3f",
          3357 => x"06",
          3358 => x"81",
          3359 => x"1a",
          3360 => x"14",
          3361 => x"2e",
          3362 => x"57",
          3363 => x"70",
          3364 => x"55",
          3365 => x"fe",
          3366 => x"80",
          3367 => x"06",
          3368 => x"72",
          3369 => x"51",
          3370 => x"81",
          3371 => x"38",
          3372 => x"80",
          3373 => x"e0",
          3374 => x"89",
          3375 => x"86",
          3376 => x"82",
          3377 => x"f2",
          3378 => x"80",
          3379 => x"e0",
          3380 => x"83",
          3381 => x"ff",
          3382 => x"52",
          3383 => x"98",
          3384 => x"85",
          3385 => x"57",
          3386 => x"39",
          3387 => x"ff",
          3388 => x"75",
          3389 => x"83",
          3390 => x"8f",
          3391 => x"74",
          3392 => x"38",
          3393 => x"81",
          3394 => x"38",
          3395 => x"54",
          3396 => x"33",
          3397 => x"08",
          3398 => x"7c",
          3399 => x"8d",
          3400 => x"81",
          3401 => x"9a",
          3402 => x"e0",
          3403 => x"74",
          3404 => x"06",
          3405 => x"75",
          3406 => x"77",
          3407 => x"98",
          3408 => x"80",
          3409 => x"80",
          3410 => x"3f",
          3411 => x"70",
          3412 => x"80",
          3413 => x"08",
          3414 => x"75",
          3415 => x"2e",
          3416 => x"5b",
          3417 => x"33",
          3418 => x"55",
          3419 => x"80",
          3420 => x"22",
          3421 => x"70",
          3422 => x"81",
          3423 => x"93",
          3424 => x"e0",
          3425 => x"7e",
          3426 => x"06",
          3427 => x"19",
          3428 => x"3f",
          3429 => x"38",
          3430 => x"0c",
          3431 => x"82",
          3432 => x"08",
          3433 => x"e0",
          3434 => x"3d",
          3435 => x"81",
          3436 => x"73",
          3437 => x"70",
          3438 => x"8d",
          3439 => x"22",
          3440 => x"a0",
          3441 => x"5f",
          3442 => x"05",
          3443 => x"82",
          3444 => x"34",
          3445 => x"58",
          3446 => x"e2",
          3447 => x"7a",
          3448 => x"06",
          3449 => x"74",
          3450 => x"55",
          3451 => x"07",
          3452 => x"81",
          3453 => x"2e",
          3454 => x"56",
          3455 => x"38",
          3456 => x"05",
          3457 => x"bf",
          3458 => x"87",
          3459 => x"ff",
          3460 => x"74",
          3461 => x"54",
          3462 => x"b5",
          3463 => x"ad",
          3464 => x"e3",
          3465 => x"2e",
          3466 => x"2e",
          3467 => x"55",
          3468 => x"70",
          3469 => x"77",
          3470 => x"16",
          3471 => x"8a",
          3472 => x"58",
          3473 => x"27",
          3474 => x"82",
          3475 => x"5b",
          3476 => x"87",
          3477 => x"38",
          3478 => x"98",
          3479 => x"df",
          3480 => x"1b",
          3481 => x"81",
          3482 => x"81",
          3483 => x"52",
          3484 => x"82",
          3485 => x"79",
          3486 => x"08",
          3487 => x"38",
          3488 => x"d4",
          3489 => x"71",
          3490 => x"3f",
          3491 => x"98",
          3492 => x"f5",
          3493 => x"ff",
          3494 => x"51",
          3495 => x"57",
          3496 => x"8c",
          3497 => x"ff",
          3498 => x"34",
          3499 => x"98",
          3500 => x"08",
          3501 => x"77",
          3502 => x"73",
          3503 => x"10",
          3504 => x"54",
          3505 => x"76",
          3506 => x"38",
          3507 => x"8c",
          3508 => x"ff",
          3509 => x"22",
          3510 => x"c0",
          3511 => x"83",
          3512 => x"f7",
          3513 => x"e0",
          3514 => x"59",
          3515 => x"52",
          3516 => x"98",
          3517 => x"38",
          3518 => x"9c",
          3519 => x"53",
          3520 => x"df",
          3521 => x"33",
          3522 => x"34",
          3523 => x"74",
          3524 => x"04",
          3525 => x"12",
          3526 => x"55",
          3527 => x"74",
          3528 => x"08",
          3529 => x"38",
          3530 => x"8d",
          3531 => x"e0",
          3532 => x"53",
          3533 => x"34",
          3534 => x"82",
          3535 => x"bf",
          3536 => x"e0",
          3537 => x"84",
          3538 => x"54",
          3539 => x"0d",
          3540 => x"08",
          3541 => x"34",
          3542 => x"38",
          3543 => x"38",
          3544 => x"70",
          3545 => x"77",
          3546 => x"70",
          3547 => x"97",
          3548 => x"ff",
          3549 => x"26",
          3550 => x"76",
          3551 => x"58",
          3552 => x"2b",
          3553 => x"82",
          3554 => x"55",
          3555 => x"76",
          3556 => x"72",
          3557 => x"55",
          3558 => x"78",
          3559 => x"52",
          3560 => x"80",
          3561 => x"55",
          3562 => x"08",
          3563 => x"54",
          3564 => x"80",
          3565 => x"53",
          3566 => x"82",
          3567 => x"5a",
          3568 => x"81",
          3569 => x"b7",
          3570 => x"84",
          3571 => x"70",
          3572 => x"54",
          3573 => x"80",
          3574 => x"05",
          3575 => x"70",
          3576 => x"8a",
          3577 => x"88",
          3578 => x"96",
          3579 => x"76",
          3580 => x"81",
          3581 => x"1a",
          3582 => x"80",
          3583 => x"56",
          3584 => x"72",
          3585 => x"8c",
          3586 => x"87",
          3587 => x"72",
          3588 => x"72",
          3589 => x"83",
          3590 => x"70",
          3591 => x"15",
          3592 => x"59",
          3593 => x"05",
          3594 => x"1c",
          3595 => x"85",
          3596 => x"08",
          3597 => x"9c",
          3598 => x"aa",
          3599 => x"96",
          3600 => x"98",
          3601 => x"d8",
          3602 => x"19",
          3603 => x"0d",
          3604 => x"70",
          3605 => x"83",
          3606 => x"92",
          3607 => x"98",
          3608 => x"81",
          3609 => x"56",
          3610 => x"83",
          3611 => x"70",
          3612 => x"51",
          3613 => x"0c",
          3614 => x"26",
          3615 => x"34",
          3616 => x"82",
          3617 => x"63",
          3618 => x"54",
          3619 => x"da",
          3620 => x"2e",
          3621 => x"82",
          3622 => x"10",
          3623 => x"55",
          3624 => x"82",
          3625 => x"70",
          3626 => x"71",
          3627 => x"73",
          3628 => x"38",
          3629 => x"52",
          3630 => x"82",
          3631 => x"81",
          3632 => x"1a",
          3633 => x"ff",
          3634 => x"70",
          3635 => x"09",
          3636 => x"80",
          3637 => x"79",
          3638 => x"74",
          3639 => x"78",
          3640 => x"79",
          3641 => x"80",
          3642 => x"06",
          3643 => x"73",
          3644 => x"38",
          3645 => x"81",
          3646 => x"80",
          3647 => x"58",
          3648 => x"a0",
          3649 => x"34",
          3650 => x"38",
          3651 => x"34",
          3652 => x"38",
          3653 => x"22",
          3654 => x"30",
          3655 => x"56",
          3656 => x"87",
          3657 => x"78",
          3658 => x"23",
          3659 => x"39",
          3660 => x"80",
          3661 => x"56",
          3662 => x"06",
          3663 => x"70",
          3664 => x"f2",
          3665 => x"ff",
          3666 => x"06",
          3667 => x"80",
          3668 => x"70",
          3669 => x"38",
          3670 => x"19",
          3671 => x"15",
          3672 => x"09",
          3673 => x"52",
          3674 => x"70",
          3675 => x"70",
          3676 => x"80",
          3677 => x"96",
          3678 => x"80",
          3679 => x"8c",
          3680 => x"83",
          3681 => x"5b",
          3682 => x"7c",
          3683 => x"80",
          3684 => x"55",
          3685 => x"2e",
          3686 => x"38",
          3687 => x"81",
          3688 => x"7c",
          3689 => x"ff",
          3690 => x"38",
          3691 => x"75",
          3692 => x"98",
          3693 => x"2a",
          3694 => x"80",
          3695 => x"82",
          3696 => x"ff",
          3697 => x"73",
          3698 => x"7f",
          3699 => x"a0",
          3700 => x"75",
          3701 => x"75",
          3702 => x"d1",
          3703 => x"98",
          3704 => x"77",
          3705 => x"bf",
          3706 => x"7b",
          3707 => x"73",
          3708 => x"e0",
          3709 => x"55",
          3710 => x"74",
          3711 => x"a0",
          3712 => x"09",
          3713 => x"1f",
          3714 => x"88",
          3715 => x"5c",
          3716 => x"8d",
          3717 => x"2e",
          3718 => x"07",
          3719 => x"51",
          3720 => x"54",
          3721 => x"07",
          3722 => x"51",
          3723 => x"88",
          3724 => x"51",
          3725 => x"ab",
          3726 => x"08",
          3727 => x"08",
          3728 => x"38",
          3729 => x"82",
          3730 => x"96",
          3731 => x"2e",
          3732 => x"1f",
          3733 => x"81",
          3734 => x"b7",
          3735 => x"51",
          3736 => x"70",
          3737 => x"55",
          3738 => x"08",
          3739 => x"52",
          3740 => x"98",
          3741 => x"75",
          3742 => x"04",
          3743 => x"08",
          3744 => x"59",
          3745 => x"70",
          3746 => x"52",
          3747 => x"ee",
          3748 => x"81",
          3749 => x"81",
          3750 => x"26",
          3751 => x"06",
          3752 => x"80",
          3753 => x"59",
          3754 => x"70",
          3755 => x"05",
          3756 => x"53",
          3757 => x"70",
          3758 => x"12",
          3759 => x"12",
          3760 => x"30",
          3761 => x"2e",
          3762 => x"be",
          3763 => x"30",
          3764 => x"2a",
          3765 => x"2e",
          3766 => x"55",
          3767 => x"39",
          3768 => x"7c",
          3769 => x"f7",
          3770 => x"0c",
          3771 => x"78",
          3772 => x"0b",
          3773 => x"d1",
          3774 => x"08",
          3775 => x"ce",
          3776 => x"ff",
          3777 => x"d4",
          3778 => x"38",
          3779 => x"74",
          3780 => x"38",
          3781 => x"30",
          3782 => x"54",
          3783 => x"09",
          3784 => x"d1",
          3785 => x"87",
          3786 => x"e0",
          3787 => x"53",
          3788 => x"51",
          3789 => x"55",
          3790 => x"38",
          3791 => x"88",
          3792 => x"02",
          3793 => x"55",
          3794 => x"3f",
          3795 => x"80",
          3796 => x"c7",
          3797 => x"82",
          3798 => x"8c",
          3799 => x"73",
          3800 => x"33",
          3801 => x"81",
          3802 => x"e0",
          3803 => x"06",
          3804 => x"2e",
          3805 => x"81",
          3806 => x"f7",
          3807 => x"77",
          3808 => x"81",
          3809 => x"51",
          3810 => x"81",
          3811 => x"83",
          3812 => x"2e",
          3813 => x"06",
          3814 => x"38",
          3815 => x"9c",
          3816 => x"06",
          3817 => x"81",
          3818 => x"19",
          3819 => x"38",
          3820 => x"83",
          3821 => x"80",
          3822 => x"cb",
          3823 => x"76",
          3824 => x"16",
          3825 => x"d7",
          3826 => x"33",
          3827 => x"31",
          3828 => x"05",
          3829 => x"08",
          3830 => x"38",
          3831 => x"82",
          3832 => x"80",
          3833 => x"58",
          3834 => x"38",
          3835 => x"77",
          3836 => x"16",
          3837 => x"81",
          3838 => x"8d",
          3839 => x"80",
          3840 => x"e0",
          3841 => x"72",
          3842 => x"d7",
          3843 => x"3f",
          3844 => x"06",
          3845 => x"51",
          3846 => x"58",
          3847 => x"33",
          3848 => x"ff",
          3849 => x"55",
          3850 => x"38",
          3851 => x"80",
          3852 => x"8a",
          3853 => x"ff",
          3854 => x"86",
          3855 => x"c9",
          3856 => x"98",
          3857 => x"15",
          3858 => x"76",
          3859 => x"c8",
          3860 => x"ff",
          3861 => x"d8",
          3862 => x"98",
          3863 => x"cb",
          3864 => x"ff",
          3865 => x"83",
          3866 => x"71",
          3867 => x"26",
          3868 => x"74",
          3869 => x"82",
          3870 => x"08",
          3871 => x"98",
          3872 => x"83",
          3873 => x"26",
          3874 => x"26",
          3875 => x"56",
          3876 => x"15",
          3877 => x"0c",
          3878 => x"1d",
          3879 => x"2e",
          3880 => x"14",
          3881 => x"08",
          3882 => x"72",
          3883 => x"80",
          3884 => x"e0",
          3885 => x"2b",
          3886 => x"2e",
          3887 => x"0c",
          3888 => x"38",
          3889 => x"81",
          3890 => x"89",
          3891 => x"08",
          3892 => x"15",
          3893 => x"80",
          3894 => x"09",
          3895 => x"14",
          3896 => x"08",
          3897 => x"2e",
          3898 => x"1b",
          3899 => x"e0",
          3900 => x"98",
          3901 => x"51",
          3902 => x"83",
          3903 => x"d5",
          3904 => x"b8",
          3905 => x"98",
          3906 => x"09",
          3907 => x"51",
          3908 => x"86",
          3909 => x"06",
          3910 => x"ea",
          3911 => x"0c",
          3912 => x"82",
          3913 => x"74",
          3914 => x"53",
          3915 => x"15",
          3916 => x"0c",
          3917 => x"75",
          3918 => x"04",
          3919 => x"73",
          3920 => x"72",
          3921 => x"71",
          3922 => x"84",
          3923 => x"09",
          3924 => x"51",
          3925 => x"08",
          3926 => x"74",
          3927 => x"78",
          3928 => x"98",
          3929 => x"0d",
          3930 => x"3d",
          3931 => x"8b",
          3932 => x"24",
          3933 => x"29",
          3934 => x"55",
          3935 => x"34",
          3936 => x"80",
          3937 => x"75",
          3938 => x"3d",
          3939 => x"3f",
          3940 => x"e0",
          3941 => x"3d",
          3942 => x"05",
          3943 => x"2e",
          3944 => x"54",
          3945 => x"84",
          3946 => x"e0",
          3947 => x"84",
          3948 => x"3d",
          3949 => x"e0",
          3950 => x"92",
          3951 => x"98",
          3952 => x"38",
          3953 => x"80",
          3954 => x"95",
          3955 => x"aa",
          3956 => x"e0",
          3957 => x"05",
          3958 => x"38",
          3959 => x"54",
          3960 => x"83",
          3961 => x"83",
          3962 => x"06",
          3963 => x"38",
          3964 => x"82",
          3965 => x"0a",
          3966 => x"3f",
          3967 => x"80",
          3968 => x"3f",
          3969 => x"db",
          3970 => x"34",
          3971 => x"b4",
          3972 => x"52",
          3973 => x"3f",
          3974 => x"98",
          3975 => x"82",
          3976 => x"84",
          3977 => x"73",
          3978 => x"ad",
          3979 => x"51",
          3980 => x"81",
          3981 => x"87",
          3982 => x"51",
          3983 => x"7b",
          3984 => x"82",
          3985 => x"83",
          3986 => x"80",
          3987 => x"58",
          3988 => x"63",
          3989 => x"57",
          3990 => x"82",
          3991 => x"9c",
          3992 => x"e0",
          3993 => x"1b",
          3994 => x"22",
          3995 => x"80",
          3996 => x"1a",
          3997 => x"85",
          3998 => x"80",
          3999 => x"08",
          4000 => x"98",
          4001 => x"70",
          4002 => x"39",
          4003 => x"82",
          4004 => x"08",
          4005 => x"e0",
          4006 => x"83",
          4007 => x"74",
          4008 => x"54",
          4009 => x"75",
          4010 => x"98",
          4011 => x"ff",
          4012 => x"76",
          4013 => x"e0",
          4014 => x"39",
          4015 => x"05",
          4016 => x"0c",
          4017 => x"98",
          4018 => x"63",
          4019 => x"7e",
          4020 => x"51",
          4021 => x"55",
          4022 => x"19",
          4023 => x"74",
          4024 => x"81",
          4025 => x"82",
          4026 => x"1a",
          4027 => x"0b",
          4028 => x"39",
          4029 => x"55",
          4030 => x"7b",
          4031 => x"08",
          4032 => x"81",
          4033 => x"05",
          4034 => x"a8",
          4035 => x"55",
          4036 => x"51",
          4037 => x"55",
          4038 => x"ff",
          4039 => x"0c",
          4040 => x"93",
          4041 => x"ff",
          4042 => x"7c",
          4043 => x"80",
          4044 => x"22",
          4045 => x"38",
          4046 => x"53",
          4047 => x"b8",
          4048 => x"d6",
          4049 => x"74",
          4050 => x"77",
          4051 => x"84",
          4052 => x"08",
          4053 => x"ff",
          4054 => x"ba",
          4055 => x"08",
          4056 => x"57",
          4057 => x"56",
          4058 => x"8d",
          4059 => x"38",
          4060 => x"06",
          4061 => x"bd",
          4062 => x"17",
          4063 => x"18",
          4064 => x"39",
          4065 => x"90",
          4066 => x"63",
          4067 => x"7e",
          4068 => x"51",
          4069 => x"55",
          4070 => x"18",
          4071 => x"74",
          4072 => x"70",
          4073 => x"56",
          4074 => x"38",
          4075 => x"82",
          4076 => x"19",
          4077 => x"18",
          4078 => x"27",
          4079 => x"2e",
          4080 => x"83",
          4081 => x"38",
          4082 => x"89",
          4083 => x"75",
          4084 => x"9c",
          4085 => x"08",
          4086 => x"e0",
          4087 => x"80",
          4088 => x"ff",
          4089 => x"38",
          4090 => x"85",
          4091 => x"b4",
          4092 => x"81",
          4093 => x"85",
          4094 => x"38",
          4095 => x"bf",
          4096 => x"2e",
          4097 => x"1b",
          4098 => x"2e",
          4099 => x"11",
          4100 => x"85",
          4101 => x"76",
          4102 => x"ff",
          4103 => x"fe",
          4104 => x"31",
          4105 => x"84",
          4106 => x"89",
          4107 => x"ff",
          4108 => x"83",
          4109 => x"de",
          4110 => x"26",
          4111 => x"3f",
          4112 => x"7e",
          4113 => x"19",
          4114 => x"84",
          4115 => x"27",
          4116 => x"52",
          4117 => x"e0",
          4118 => x"7c",
          4119 => x"1f",
          4120 => x"7e",
          4121 => x"76",
          4122 => x"1e",
          4123 => x"0c",
          4124 => x"74",
          4125 => x"8c",
          4126 => x"33",
          4127 => x"34",
          4128 => x"90",
          4129 => x"8b",
          4130 => x"f2",
          4131 => x"82",
          4132 => x"16",
          4133 => x"51",
          4134 => x"38",
          4135 => x"bb",
          4136 => x"82",
          4137 => x"16",
          4138 => x"55",
          4139 => x"53",
          4140 => x"3f",
          4141 => x"ff",
          4142 => x"52",
          4143 => x"76",
          4144 => x"3f",
          4145 => x"78",
          4146 => x"98",
          4147 => x"55",
          4148 => x"e0",
          4149 => x"3d",
          4150 => x"3f",
          4151 => x"98",
          4152 => x"52",
          4153 => x"98",
          4154 => x"38",
          4155 => x"82",
          4156 => x"ff",
          4157 => x"3f",
          4158 => x"08",
          4159 => x"82",
          4160 => x"e0",
          4161 => x"3d",
          4162 => x"52",
          4163 => x"e0",
          4164 => x"80",
          4165 => x"3d",
          4166 => x"e0",
          4167 => x"bc",
          4168 => x"98",
          4169 => x"38",
          4170 => x"39",
          4171 => x"70",
          4172 => x"2e",
          4173 => x"54",
          4174 => x"98",
          4175 => x"08",
          4176 => x"85",
          4177 => x"3d",
          4178 => x"e1",
          4179 => x"5b",
          4180 => x"3d",
          4181 => x"51",
          4182 => x"57",
          4183 => x"7b",
          4184 => x"11",
          4185 => x"80",
          4186 => x"82",
          4187 => x"70",
          4188 => x"98",
          4189 => x"ef",
          4190 => x"51",
          4191 => x"08",
          4192 => x"38",
          4193 => x"c8",
          4194 => x"d6",
          4195 => x"d4",
          4196 => x"e0",
          4197 => x"74",
          4198 => x"08",
          4199 => x"80",
          4200 => x"8b",
          4201 => x"a6",
          4202 => x"3f",
          4203 => x"98",
          4204 => x"2e",
          4205 => x"81",
          4206 => x"df",
          4207 => x"d6",
          4208 => x"82",
          4209 => x"80",
          4210 => x"55",
          4211 => x"56",
          4212 => x"73",
          4213 => x"2e",
          4214 => x"ff",
          4215 => x"18",
          4216 => x"33",
          4217 => x"80",
          4218 => x"74",
          4219 => x"09",
          4220 => x"e1",
          4221 => x"34",
          4222 => x"84",
          4223 => x"70",
          4224 => x"76",
          4225 => x"70",
          4226 => x"82",
          4227 => x"80",
          4228 => x"19",
          4229 => x"5c",
          4230 => x"7a",
          4231 => x"2e",
          4232 => x"97",
          4233 => x"19",
          4234 => x"05",
          4235 => x"80",
          4236 => x"80",
          4237 => x"7b",
          4238 => x"53",
          4239 => x"98",
          4240 => x"fe",
          4241 => x"f6",
          4242 => x"27",
          4243 => x"2a",
          4244 => x"83",
          4245 => x"80",
          4246 => x"2e",
          4247 => x"70",
          4248 => x"2e",
          4249 => x"fe",
          4250 => x"ff",
          4251 => x"fe",
          4252 => x"73",
          4253 => x"06",
          4254 => x"98",
          4255 => x"39",
          4256 => x"73",
          4257 => x"82",
          4258 => x"08",
          4259 => x"98",
          4260 => x"e0",
          4261 => x"16",
          4262 => x"76",
          4263 => x"31",
          4264 => x"90",
          4265 => x"06",
          4266 => x"9b",
          4267 => x"81",
          4268 => x"e0",
          4269 => x"08",
          4270 => x"ff",
          4271 => x"54",
          4272 => x"27",
          4273 => x"08",
          4274 => x"ff",
          4275 => x"16",
          4276 => x"80",
          4277 => x"ff",
          4278 => x"94",
          4279 => x"53",
          4280 => x"34",
          4281 => x"82",
          4282 => x"08",
          4283 => x"38",
          4284 => x"80",
          4285 => x"73",
          4286 => x"8c",
          4287 => x"38",
          4288 => x"82",
          4289 => x"f9",
          4290 => x"80",
          4291 => x"3d",
          4292 => x"51",
          4293 => x"55",
          4294 => x"77",
          4295 => x"dd",
          4296 => x"e0",
          4297 => x"33",
          4298 => x"24",
          4299 => x"2a",
          4300 => x"80",
          4301 => x"77",
          4302 => x"08",
          4303 => x"22",
          4304 => x"ff",
          4305 => x"55",
          4306 => x"38",
          4307 => x"84",
          4308 => x"82",
          4309 => x"fc",
          4310 => x"53",
          4311 => x"e0",
          4312 => x"08",
          4313 => x"3d",
          4314 => x"54",
          4315 => x"82",
          4316 => x"08",
          4317 => x"e0",
          4318 => x"fc",
          4319 => x"cb",
          4320 => x"51",
          4321 => x"53",
          4322 => x"81",
          4323 => x"82",
          4324 => x"73",
          4325 => x"51",
          4326 => x"08",
          4327 => x"9f",
          4328 => x"51",
          4329 => x"0c",
          4330 => x"66",
          4331 => x"97",
          4332 => x"e0",
          4333 => x"b2",
          4334 => x"3f",
          4335 => x"98",
          4336 => x"33",
          4337 => x"25",
          4338 => x"80",
          4339 => x"ce",
          4340 => x"95",
          4341 => x"65",
          4342 => x"05",
          4343 => x"82",
          4344 => x"08",
          4345 => x"08",
          4346 => x"08",
          4347 => x"91",
          4348 => x"81",
          4349 => x"c9",
          4350 => x"55",
          4351 => x"80",
          4352 => x"52",
          4353 => x"f5",
          4354 => x"cf",
          4355 => x"cc",
          4356 => x"82",
          4357 => x"05",
          4358 => x"9c",
          4359 => x"f9",
          4360 => x"08",
          4361 => x"81",
          4362 => x"3f",
          4363 => x"98",
          4364 => x"77",
          4365 => x"74",
          4366 => x"b8",
          4367 => x"e0",
          4368 => x"30",
          4369 => x"5b",
          4370 => x"ff",
          4371 => x"f0",
          4372 => x"1b",
          4373 => x"83",
          4374 => x"92",
          4375 => x"12",
          4376 => x"54",
          4377 => x"98",
          4378 => x"0d",
          4379 => x"52",
          4380 => x"08",
          4381 => x"38",
          4382 => x"38",
          4383 => x"81",
          4384 => x"80",
          4385 => x"54",
          4386 => x"38",
          4387 => x"53",
          4388 => x"b2",
          4389 => x"88",
          4390 => x"17",
          4391 => x"3f",
          4392 => x"81",
          4393 => x"98",
          4394 => x"38",
          4395 => x"77",
          4396 => x"08",
          4397 => x"82",
          4398 => x"b1",
          4399 => x"94",
          4400 => x"33",
          4401 => x"34",
          4402 => x"18",
          4403 => x"0c",
          4404 => x"82",
          4405 => x"a3",
          4406 => x"98",
          4407 => x"f9",
          4408 => x"96",
          4409 => x"82",
          4410 => x"08",
          4411 => x"33",
          4412 => x"55",
          4413 => x"75",
          4414 => x"c1",
          4415 => x"81",
          4416 => x"b1",
          4417 => x"c3",
          4418 => x"2a",
          4419 => x"80",
          4420 => x"e0",
          4421 => x"89",
          4422 => x"5c",
          4423 => x"ff",
          4424 => x"55",
          4425 => x"82",
          4426 => x"bb",
          4427 => x"82",
          4428 => x"80",
          4429 => x"2e",
          4430 => x"c1",
          4431 => x"e0",
          4432 => x"70",
          4433 => x"51",
          4434 => x"73",
          4435 => x"52",
          4436 => x"e0",
          4437 => x"51",
          4438 => x"08",
          4439 => x"3d",
          4440 => x"9a",
          4441 => x"51",
          4442 => x"54",
          4443 => x"78",
          4444 => x"58",
          4445 => x"54",
          4446 => x"54",
          4447 => x"84",
          4448 => x"02",
          4449 => x"81",
          4450 => x"fd",
          4451 => x"70",
          4452 => x"e0",
          4453 => x"98",
          4454 => x"98",
          4455 => x"38",
          4456 => x"2e",
          4457 => x"81",
          4458 => x"e0",
          4459 => x"9c",
          4460 => x"e0",
          4461 => x"a0",
          4462 => x"3f",
          4463 => x"78",
          4464 => x"82",
          4465 => x"51",
          4466 => x"b8",
          4467 => x"a0",
          4468 => x"05",
          4469 => x"ae",
          4470 => x"78",
          4471 => x"cc",
          4472 => x"34",
          4473 => x"e0",
          4474 => x"b3",
          4475 => x"96",
          4476 => x"53",
          4477 => x"3f",
          4478 => x"78",
          4479 => x"51",
          4480 => x"08",
          4481 => x"76",
          4482 => x"e0",
          4483 => x"3d",
          4484 => x"d0",
          4485 => x"05",
          4486 => x"82",
          4487 => x"08",
          4488 => x"08",
          4489 => x"cd",
          4490 => x"e0",
          4491 => x"9f",
          4492 => x"55",
          4493 => x"3d",
          4494 => x"51",
          4495 => x"52",
          4496 => x"92",
          4497 => x"c8",
          4498 => x"82",
          4499 => x"3d",
          4500 => x"65",
          4501 => x"55",
          4502 => x"84",
          4503 => x"73",
          4504 => x"98",
          4505 => x"ca",
          4506 => x"ff",
          4507 => x"a1",
          4508 => x"17",
          4509 => x"70",
          4510 => x"38",
          4511 => x"34",
          4512 => x"8b",
          4513 => x"06",
          4514 => x"e7",
          4515 => x"75",
          4516 => x"82",
          4517 => x"a5",
          4518 => x"08",
          4519 => x"98",
          4520 => x"3f",
          4521 => x"11",
          4522 => x"80",
          4523 => x"ae",
          4524 => x"53",
          4525 => x"3f",
          4526 => x"87",
          4527 => x"77",
          4528 => x"08",
          4529 => x"78",
          4530 => x"98",
          4531 => x"aa",
          4532 => x"80",
          4533 => x"e3",
          4534 => x"3d",
          4535 => x"c3",
          4536 => x"e0",
          4537 => x"66",
          4538 => x"c5",
          4539 => x"e0",
          4540 => x"05",
          4541 => x"73",
          4542 => x"09",
          4543 => x"06",
          4544 => x"15",
          4545 => x"34",
          4546 => x"e0",
          4547 => x"0c",
          4548 => x"65",
          4549 => x"52",
          4550 => x"e0",
          4551 => x"80",
          4552 => x"3d",
          4553 => x"e0",
          4554 => x"b4",
          4555 => x"a0",
          4556 => x"84",
          4557 => x"2b",
          4558 => x"9d",
          4559 => x"15",
          4560 => x"82",
          4561 => x"98",
          4562 => x"0d",
          4563 => x"3d",
          4564 => x"db",
          4565 => x"98",
          4566 => x"07",
          4567 => x"2e",
          4568 => x"55",
          4569 => x"7b",
          4570 => x"70",
          4571 => x"e0",
          4572 => x"80",
          4573 => x"b1",
          4574 => x"82",
          4575 => x"98",
          4576 => x"59",
          4577 => x"56",
          4578 => x"16",
          4579 => x"56",
          4580 => x"80",
          4581 => x"70",
          4582 => x"e8",
          4583 => x"81",
          4584 => x"57",
          4585 => x"51",
          4586 => x"73",
          4587 => x"08",
          4588 => x"e0",
          4589 => x"a7",
          4590 => x"c3",
          4591 => x"e4",
          4592 => x"56",
          4593 => x"92",
          4594 => x"76",
          4595 => x"04",
          4596 => x"ff",
          4597 => x"d3",
          4598 => x"98",
          4599 => x"82",
          4600 => x"3d",
          4601 => x"73",
          4602 => x"74",
          4603 => x"3d",
          4604 => x"98",
          4605 => x"38",
          4606 => x"3f",
          4607 => x"51",
          4608 => x"83",
          4609 => x"a3",
          4610 => x"ff",
          4611 => x"93",
          4612 => x"75",
          4613 => x"76",
          4614 => x"39",
          4615 => x"88",
          4616 => x"59",
          4617 => x"81",
          4618 => x"33",
          4619 => x"fe",
          4620 => x"73",
          4621 => x"80",
          4622 => x"75",
          4623 => x"2e",
          4624 => x"56",
          4625 => x"80",
          4626 => x"a8",
          4627 => x"82",
          4628 => x"52",
          4629 => x"e0",
          4630 => x"8d",
          4631 => x"e5",
          4632 => x"98",
          4633 => x"cc",
          4634 => x"c4",
          4635 => x"d8",
          4636 => x"e0",
          4637 => x"e0",
          4638 => x"c5",
          4639 => x"34",
          4640 => x"99",
          4641 => x"15",
          4642 => x"82",
          4643 => x"82",
          4644 => x"f2",
          4645 => x"80",
          4646 => x"55",
          4647 => x"3f",
          4648 => x"98",
          4649 => x"58",
          4650 => x"97",
          4651 => x"38",
          4652 => x"81",
          4653 => x"87",
          4654 => x"90",
          4655 => x"8a",
          4656 => x"7f",
          4657 => x"3f",
          4658 => x"72",
          4659 => x"05",
          4660 => x"55",
          4661 => x"16",
          4662 => x"76",
          4663 => x"79",
          4664 => x"7f",
          4665 => x"83",
          4666 => x"81",
          4667 => x"08",
          4668 => x"98",
          4669 => x"7b",
          4670 => x"39",
          4671 => x"09",
          4672 => x"80",
          4673 => x"78",
          4674 => x"38",
          4675 => x"81",
          4676 => x"74",
          4677 => x"82",
          4678 => x"08",
          4679 => x"16",
          4680 => x"39",
          4681 => x"0c",
          4682 => x"88",
          4683 => x"1a",
          4684 => x"1b",
          4685 => x"16",
          4686 => x"38",
          4687 => x"15",
          4688 => x"34",
          4689 => x"90",
          4690 => x"6e",
          4691 => x"9e",
          4692 => x"3f",
          4693 => x"08",
          4694 => x"08",
          4695 => x"08",
          4696 => x"80",
          4697 => x"e0",
          4698 => x"33",
          4699 => x"55",
          4700 => x"3f",
          4701 => x"70",
          4702 => x"8c",
          4703 => x"06",
          4704 => x"38",
          4705 => x"7f",
          4706 => x"98",
          4707 => x"2e",
          4708 => x"8b",
          4709 => x"80",
          4710 => x"2e",
          4711 => x"38",
          4712 => x"ff",
          4713 => x"86",
          4714 => x"89",
          4715 => x"77",
          4716 => x"81",
          4717 => x"07",
          4718 => x"38",
          4719 => x"54",
          4720 => x"8e",
          4721 => x"08",
          4722 => x"ff",
          4723 => x"83",
          4724 => x"82",
          4725 => x"a3",
          4726 => x"11",
          4727 => x"93",
          4728 => x"da",
          4729 => x"18",
          4730 => x"e0",
          4731 => x"f8",
          4732 => x"90",
          4733 => x"08",
          4734 => x"77",
          4735 => x"55",
          4736 => x"8e",
          4737 => x"74",
          4738 => x"68",
          4739 => x"81",
          4740 => x"2a",
          4741 => x"2e",
          4742 => x"82",
          4743 => x"55",
          4744 => x"81",
          4745 => x"80",
          4746 => x"83",
          4747 => x"78",
          4748 => x"0b",
          4749 => x"80",
          4750 => x"38",
          4751 => x"17",
          4752 => x"2e",
          4753 => x"79",
          4754 => x"82",
          4755 => x"05",
          4756 => x"80",
          4757 => x"8a",
          4758 => x"75",
          4759 => x"78",
          4760 => x"0b",
          4761 => x"80",
          4762 => x"38",
          4763 => x"17",
          4764 => x"2e",
          4765 => x"79",
          4766 => x"82",
          4767 => x"82",
          4768 => x"38",
          4769 => x"82",
          4770 => x"2a",
          4771 => x"17",
          4772 => x"7b",
          4773 => x"12",
          4774 => x"74",
          4775 => x"7d",
          4776 => x"76",
          4777 => x"76",
          4778 => x"60",
          4779 => x"26",
          4780 => x"31",
          4781 => x"fe",
          4782 => x"58",
          4783 => x"38",
          4784 => x"26",
          4785 => x"79",
          4786 => x"87",
          4787 => x"06",
          4788 => x"82",
          4789 => x"8f",
          4790 => x"26",
          4791 => x"63",
          4792 => x"38",
          4793 => x"98",
          4794 => x"86",
          4795 => x"79",
          4796 => x"80",
          4797 => x"83",
          4798 => x"8b",
          4799 => x"74",
          4800 => x"52",
          4801 => x"53",
          4802 => x"8f",
          4803 => x"51",
          4804 => x"34",
          4805 => x"1b",
          4806 => x"90",
          4807 => x"70",
          4808 => x"55",
          4809 => x"67",
          4810 => x"38",
          4811 => x"1b",
          4812 => x"74",
          4813 => x"3f",
          4814 => x"98",
          4815 => x"ff",
          4816 => x"3f",
          4817 => x"db",
          4818 => x"80",
          4819 => x"80",
          4820 => x"7c",
          4821 => x"3f",
          4822 => x"b3",
          4823 => x"8d",
          4824 => x"ff",
          4825 => x"c0",
          4826 => x"34",
          4827 => x"c7",
          4828 => x"0a",
          4829 => x"3f",
          4830 => x"1b",
          4831 => x"0b",
          4832 => x"34",
          4833 => x"1b",
          4834 => x"d5",
          4835 => x"ff",
          4836 => x"7a",
          4837 => x"81",
          4838 => x"38",
          4839 => x"ec",
          4840 => x"52",
          4841 => x"80",
          4842 => x"e5",
          4843 => x"7a",
          4844 => x"85",
          4845 => x"ff",
          4846 => x"e8",
          4847 => x"52",
          4848 => x"3f",
          4849 => x"8b",
          4850 => x"7a",
          4851 => x"75",
          4852 => x"51",
          4853 => x"52",
          4854 => x"56",
          4855 => x"06",
          4856 => x"8b",
          4857 => x"ff",
          4858 => x"1b",
          4859 => x"55",
          4860 => x"74",
          4861 => x"7c",
          4862 => x"38",
          4863 => x"52",
          4864 => x"e0",
          4865 => x"53",
          4866 => x"ff",
          4867 => x"31",
          4868 => x"58",
          4869 => x"55",
          4870 => x"61",
          4871 => x"57",
          4872 => x"51",
          4873 => x"08",
          4874 => x"31",
          4875 => x"7d",
          4876 => x"83",
          4877 => x"7d",
          4878 => x"80",
          4879 => x"7a",
          4880 => x"81",
          4881 => x"38",
          4882 => x"b2",
          4883 => x"08",
          4884 => x"d4",
          4885 => x"81",
          4886 => x"80",
          4887 => x"fd",
          4888 => x"ff",
          4889 => x"77",
          4890 => x"81",
          4891 => x"34",
          4892 => x"80",
          4893 => x"ea",
          4894 => x"e0",
          4895 => x"75",
          4896 => x"87",
          4897 => x"51",
          4898 => x"ca",
          4899 => x"54",
          4900 => x"84",
          4901 => x"08",
          4902 => x"51",
          4903 => x"e0",
          4904 => x"56",
          4905 => x"e0",
          4906 => x"0c",
          4907 => x"7d",
          4908 => x"05",
          4909 => x"38",
          4910 => x"53",
          4911 => x"3f",
          4912 => x"38",
          4913 => x"db",
          4914 => x"34",
          4915 => x"81",
          4916 => x"55",
          4917 => x"e0",
          4918 => x"3d",
          4919 => x"33",
          4920 => x"06",
          4921 => x"3f",
          4922 => x"be",
          4923 => x"05",
          4924 => x"56",
          4925 => x"fc",
          4926 => x"76",
          4927 => x"32",
          4928 => x"70",
          4929 => x"18",
          4930 => x"3d",
          4931 => x"11",
          4932 => x"38",
          4933 => x"8c",
          4934 => x"3f",
          4935 => x"16",
          4936 => x"38",
          4937 => x"55",
          4938 => x"0d",
          4939 => x"cc",
          4940 => x"d5",
          4941 => x"04",
          4942 => x"33",
          4943 => x"54",
          4944 => x"ae",
          4945 => x"3d",
          4946 => x"84",
          4947 => x"52",
          4948 => x"83",
          4949 => x"83",
          4950 => x"b5",
          4951 => x"80",
          4952 => x"51",
          4953 => x"70",
          4954 => x"80",
          4955 => x"d3",
          4956 => x"39",
          4957 => x"53",
          4958 => x"3d",
          4959 => x"05",
          4960 => x"53",
          4961 => x"85",
          4962 => x"b5",
          4963 => x"81",
          4964 => x"d1",
          4965 => x"82",
          4966 => x"fb",
          4967 => x"ff",
          4968 => x"ff",
          4969 => x"ff",
          4970 => x"56",
          4971 => x"30",
          4972 => x"51",
          4973 => x"70",
          4974 => x"71",
          4975 => x"55",
          4976 => x"73",
          4977 => x"29",
          4978 => x"04",
          4979 => x"22",
          4980 => x"75",
          4981 => x"51",
          4982 => x"e0",
          4983 => x"95",
          4984 => x"12",
          4985 => x"85",
          4986 => x"ff",
          4987 => x"f8",
          4988 => x"39",
          4989 => x"87",
          4990 => x"ff",
          4991 => x"ff",
          4992 => x"00",
          4993 => x"00",
          4994 => x"00",
          4995 => x"00",
          4996 => x"00",
          4997 => x"00",
          4998 => x"00",
          4999 => x"00",
          5000 => x"00",
          5001 => x"00",
          5002 => x"00",
          5003 => x"00",
          5004 => x"00",
          5005 => x"00",
          5006 => x"00",
          5007 => x"00",
          5008 => x"00",
          5009 => x"00",
          5010 => x"00",
          5011 => x"00",
          5012 => x"00",
          5013 => x"00",
          5014 => x"00",
          5015 => x"00",
          5016 => x"00",
          5017 => x"00",
          5018 => x"00",
          5019 => x"00",
          5020 => x"00",
          5021 => x"00",
          5022 => x"00",
          5023 => x"00",
          5024 => x"00",
          5025 => x"00",
          5026 => x"00",
          5027 => x"00",
          5028 => x"00",
          5029 => x"00",
          5030 => x"00",
          5031 => x"00",
          5032 => x"00",
          5033 => x"00",
          5034 => x"00",
          5035 => x"00",
          5036 => x"00",
          5037 => x"00",
          5038 => x"00",
          5039 => x"00",
          5040 => x"00",
          5041 => x"00",
          5042 => x"00",
          5043 => x"00",
          5044 => x"00",
          5045 => x"00",
          5046 => x"00",
          5047 => x"00",
          5048 => x"00",
          5049 => x"00",
          5050 => x"00",
          5051 => x"00",
          5052 => x"00",
          5053 => x"00",
          5054 => x"00",
          5055 => x"00",
          5056 => x"00",
          5057 => x"00",
          5058 => x"00",
          5059 => x"00",
          5060 => x"00",
          5061 => x"00",
          5062 => x"00",
          5063 => x"00",
          5064 => x"64",
          5065 => x"64",
          5066 => x"66",
          5067 => x"66",
          5068 => x"66",
          5069 => x"6d",
          5070 => x"6d",
          5071 => x"6d",
          5072 => x"6d",
          5073 => x"6d",
          5074 => x"6d",
          5075 => x"68",
          5076 => x"68",
          5077 => x"00",
          5078 => x"72",
          5079 => x"72",
          5080 => x"69",
          5081 => x"74",
          5082 => x"6d",
          5083 => x"6b",
          5084 => x"65",
          5085 => x"20",
          5086 => x"49",
          5087 => x"20",
          5088 => x"44",
          5089 => x"20",
          5090 => x"4e",
          5091 => x"66",
          5092 => x"4e",
          5093 => x"66",
          5094 => x"49",
          5095 => x"66",
          5096 => x"2e",
          5097 => x"73",
          5098 => x"64",
          5099 => x"20",
          5100 => x"20",
          5101 => x"00",
          5102 => x"20",
          5103 => x"69",
          5104 => x"00",
          5105 => x"73",
          5106 => x"70",
          5107 => x"64",
          5108 => x"65",
          5109 => x"20",
          5110 => x"6c",
          5111 => x"44",
          5112 => x"20",
          5113 => x"2e",
          5114 => x"6f",
          5115 => x"65",
          5116 => x"73",
          5117 => x"6e",
          5118 => x"73",
          5119 => x"61",
          5120 => x"65",
          5121 => x"6f",
          5122 => x"72",
          5123 => x"61",
          5124 => x"2e",
          5125 => x"20",
          5126 => x"65",
          5127 => x"66",
          5128 => x"20",
          5129 => x"00",
          5130 => x"6d",
          5131 => x"6e",
          5132 => x"00",
          5133 => x"6d",
          5134 => x"6e",
          5135 => x"2e",
          5136 => x"65",
          5137 => x"55",
          5138 => x"65",
          5139 => x"0a",
          5140 => x"65",
          5141 => x"20",
          5142 => x"65",
          5143 => x"00",
          5144 => x"00",
          5145 => x"58",
          5146 => x"25",
          5147 => x"20",
          5148 => x"00",
          5149 => x"00",
          5150 => x"20",
          5151 => x"7a",
          5152 => x"73",
          5153 => x"32",
          5154 => x"76",
          5155 => x"20",
          5156 => x"76",
          5157 => x"25",
          5158 => x"0a",
          5159 => x"49",
          5160 => x"74",
          5161 => x"72",
          5162 => x"72",
          5163 => x"75",
          5164 => x"69",
          5165 => x"74",
          5166 => x"4c",
          5167 => x"65",
          5168 => x"49",
          5169 => x"20",
          5170 => x"70",
          5171 => x"30",
          5172 => x"65",
          5173 => x"55",
          5174 => x"20",
          5175 => x"70",
          5176 => x"31",
          5177 => x"65",
          5178 => x"55",
          5179 => x"20",
          5180 => x"70",
          5181 => x"69",
          5182 => x"69",
          5183 => x"45",
          5184 => x"20",
          5185 => x"2e",
          5186 => x"65",
          5187 => x"00",
          5188 => x"7a",
          5189 => x"30",
          5190 => x"65",
          5191 => x"69",
          5192 => x"20",
          5193 => x"20",
          5194 => x"73",
          5195 => x"6d",
          5196 => x"2e",
          5197 => x"43",
          5198 => x"2e",
          5199 => x"43",
          5200 => x"2e",
          5201 => x"61",
          5202 => x"00",
          5203 => x"78",
          5204 => x"3e",
          5205 => x"30",
          5206 => x"44",
          5207 => x"6f",
          5208 => x"70",
          5209 => x"25",
          5210 => x"32",
          5211 => x"25",
          5212 => x"34",
          5213 => x"58",
          5214 => x"00",
          5215 => x"75",
          5216 => x"64",
          5217 => x"6c",
          5218 => x"43",
          5219 => x"63",
          5220 => x"30",
          5221 => x"0a",
          5222 => x"20",
          5223 => x"64",
          5224 => x"25",
          5225 => x"52",
          5226 => x"6e",
          5227 => x"63",
          5228 => x"2e",
          5229 => x"20",
          5230 => x"6e",
          5231 => x"5a",
          5232 => x"25",
          5233 => x"73",
          5234 => x"25",
          5235 => x"73",
          5236 => x"25",
          5237 => x"63",
          5238 => x"00",
          5239 => x"72",
          5240 => x"73",
          5241 => x"6e",
          5242 => x"63",
          5243 => x"6d",
          5244 => x"52",
          5245 => x"2e",
          5246 => x"6c",
          5247 => x"65",
          5248 => x"2e",
          5249 => x"64",
          5250 => x"25",
          5251 => x"25",
          5252 => x"43",
          5253 => x"61",
          5254 => x"20",
          5255 => x"6f",
          5256 => x"67",
          5257 => x"76",
          5258 => x"70",
          5259 => x"64",
          5260 => x"57",
          5261 => x"20",
          5262 => x"25",
          5263 => x"20",
          5264 => x"4d",
          5265 => x"30",
          5266 => x"29",
          5267 => x"49",
          5268 => x"4d",
          5269 => x"25",
          5270 => x"20",
          5271 => x"20",
          5272 => x"30",
          5273 => x"29",
          5274 => x"52",
          5275 => x"20",
          5276 => x"25",
          5277 => x"20",
          5278 => x"41",
          5279 => x"65",
          5280 => x"25",
          5281 => x"20",
          5282 => x"52",
          5283 => x"69",
          5284 => x"25",
          5285 => x"20",
          5286 => x"20",
          5287 => x"68",
          5288 => x"25",
          5289 => x"20",
          5290 => x"42",
          5291 => x"00",
          5292 => x"57",
          5293 => x"20",
          5294 => x"4c",
          5295 => x"50",
          5296 => x"53",
          5297 => x"65",
          5298 => x"20",
          5299 => x"52",
          5300 => x"63",
          5301 => x"72",
          5302 => x"30",
          5303 => x"20",
          5304 => x"4d",
          5305 => x"74",
          5306 => x"72",
          5307 => x"30",
          5308 => x"20",
          5309 => x"6b",
          5310 => x"41",
          5311 => x"20",
          5312 => x"30",
          5313 => x"4d",
          5314 => x"20",
          5315 => x"49",
          5316 => x"20",
          5317 => x"20",
          5318 => x"30",
          5319 => x"20",
          5320 => x"65",
          5321 => x"20",
          5322 => x"20",
          5323 => x"64",
          5324 => x"7a",
          5325 => x"53",
          5326 => x"6f",
          5327 => x"20",
          5328 => x"20",
          5329 => x"34",
          5330 => x"20",
          5331 => x"62",
          5332 => x"41",
          5333 => x"20",
          5334 => x"64",
          5335 => x"7a",
          5336 => x"6c",
          5337 => x"75",
          5338 => x"00",
          5339 => x"45",
          5340 => x"55",
          5341 => x"00",
          5342 => x"00",
          5343 => x"01",
          5344 => x"00",
          5345 => x"00",
          5346 => x"01",
          5347 => x"00",
          5348 => x"00",
          5349 => x"01",
          5350 => x"00",
          5351 => x"00",
          5352 => x"01",
          5353 => x"00",
          5354 => x"00",
          5355 => x"01",
          5356 => x"00",
          5357 => x"00",
          5358 => x"04",
          5359 => x"00",
          5360 => x"00",
          5361 => x"04",
          5362 => x"00",
          5363 => x"00",
          5364 => x"04",
          5365 => x"00",
          5366 => x"00",
          5367 => x"04",
          5368 => x"00",
          5369 => x"00",
          5370 => x"03",
          5371 => x"00",
          5372 => x"00",
          5373 => x"03",
          5374 => x"1b",
          5375 => x"1b",
          5376 => x"1b",
          5377 => x"1b",
          5378 => x"1b",
          5379 => x"1b",
          5380 => x"0e",
          5381 => x"0b",
          5382 => x"06",
          5383 => x"04",
          5384 => x"02",
          5385 => x"68",
          5386 => x"68",
          5387 => x"21",
          5388 => x"75",
          5389 => x"46",
          5390 => x"6f",
          5391 => x"74",
          5392 => x"6f",
          5393 => x"20",
          5394 => x"00",
          5395 => x"6f",
          5396 => x"63",
          5397 => x"69",
          5398 => x"69",
          5399 => x"61",
          5400 => x"53",
          5401 => x"3e",
          5402 => x"2b",
          5403 => x"46",
          5404 => x"32",
          5405 => x"53",
          5406 => x"4e",
          5407 => x"20",
          5408 => x"20",
          5409 => x"41",
          5410 => x"41",
          5411 => x"00",
          5412 => x"00",
          5413 => x"01",
          5414 => x"14",
          5415 => x"80",
          5416 => x"45",
          5417 => x"90",
          5418 => x"59",
          5419 => x"41",
          5420 => x"a8",
          5421 => x"b0",
          5422 => x"b8",
          5423 => x"c0",
          5424 => x"c8",
          5425 => x"d0",
          5426 => x"d8",
          5427 => x"e0",
          5428 => x"e8",
          5429 => x"f0",
          5430 => x"f8",
          5431 => x"2b",
          5432 => x"5c",
          5433 => x"7f",
          5434 => x"00",
          5435 => x"00",
          5436 => x"00",
          5437 => x"00",
          5438 => x"00",
          5439 => x"00",
          5440 => x"00",
          5441 => x"00",
          5442 => x"00",
          5443 => x"00",
          5444 => x"00",
          5445 => x"20",
          5446 => x"00",
          5447 => x"00",
          5448 => x"00",
          5449 => x"00",
          5450 => x"25",
          5451 => x"25",
          5452 => x"25",
          5453 => x"25",
          5454 => x"25",
          5455 => x"25",
          5456 => x"25",
          5457 => x"25",
          5458 => x"25",
          5459 => x"25",
          5460 => x"25",
          5461 => x"25",
          5462 => x"03",
          5463 => x"00",
          5464 => x"03",
          5465 => x"03",
          5466 => x"22",
          5467 => x"00",
          5468 => x"00",
          5469 => x"25",
          5470 => x"00",
          5471 => x"00",
          5472 => x"01",
          5473 => x"01",
          5474 => x"01",
          5475 => x"01",
          5476 => x"01",
          5477 => x"01",
          5478 => x"01",
          5479 => x"01",
          5480 => x"01",
          5481 => x"01",
          5482 => x"01",
          5483 => x"01",
          5484 => x"01",
          5485 => x"01",
          5486 => x"01",
          5487 => x"01",
          5488 => x"01",
          5489 => x"01",
          5490 => x"01",
          5491 => x"01",
          5492 => x"01",
          5493 => x"01",
          5494 => x"01",
          5495 => x"01",
          5496 => x"00",
          5497 => x"01",
          5498 => x"02",
          5499 => x"02",
          5500 => x"02",
          5501 => x"01",
          5502 => x"01",
          5503 => x"02",
          5504 => x"02",
          5505 => x"01",
          5506 => x"02",
          5507 => x"01",
          5508 => x"02",
          5509 => x"02",
          5510 => x"02",
          5511 => x"02",
          5512 => x"02",
          5513 => x"01",
          5514 => x"02",
          5515 => x"01",
          5516 => x"02",
          5517 => x"02",
          5518 => x"00",
          5519 => x"03",
          5520 => x"03",
          5521 => x"03",
          5522 => x"03",
          5523 => x"03",
          5524 => x"01",
          5525 => x"03",
          5526 => x"03",
          5527 => x"03",
          5528 => x"07",
          5529 => x"01",
          5530 => x"00",
          5531 => x"05",
          5532 => x"1d",
          5533 => x"01",
          5534 => x"06",
          5535 => x"06",
          5536 => x"06",
          5537 => x"1f",
          5538 => x"1f",
          5539 => x"1f",
          5540 => x"1f",
          5541 => x"1f",
          5542 => x"1f",
          5543 => x"1f",
          5544 => x"1f",
          5545 => x"1f",
          5546 => x"1f",
          5547 => x"06",
          5548 => x"00",
          5549 => x"1f",
          5550 => x"21",
          5551 => x"21",
          5552 => x"04",
          5553 => x"01",
          5554 => x"01",
          5555 => x"03",
          5556 => x"00",
          5557 => x"00",
          5558 => x"00",
          5559 => x"00",
          5560 => x"00",
          5561 => x"00",
          5562 => x"00",
          5563 => x"00",
          5564 => x"00",
          5565 => x"00",
          5566 => x"00",
          5567 => x"00",
          5568 => x"00",
          5569 => x"00",
          5570 => x"00",
          5571 => x"00",
          5572 => x"00",
          5573 => x"00",
          5574 => x"00",
          5575 => x"00",
          5576 => x"00",
          5577 => x"00",
          5578 => x"00",
          5579 => x"00",
          5580 => x"00",
          5581 => x"00",
          5582 => x"00",
          5583 => x"00",
          5584 => x"00",
          5585 => x"00",
          5586 => x"00",
          5587 => x"00",
          5588 => x"00",
          5589 => x"00",
          5590 => x"00",
          5591 => x"00",
          5592 => x"00",
          5593 => x"00",
          5594 => x"00",
          5595 => x"00",
          5596 => x"00",
          5597 => x"00",
          5598 => x"00",
          5599 => x"00",
          5600 => x"00",
          5601 => x"00",
          5602 => x"00",
          5603 => x"00",
          5604 => x"00",
          5605 => x"00",
          5606 => x"00",
          5607 => x"00",
          5608 => x"00",
          5609 => x"00",
          5610 => x"00",
          5611 => x"01",
          5612 => x"00",
          5613 => x"00",
          5614 => x"05",
          5615 => x"00",
          5616 => x"01",
          5617 => x"01",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"00",
          5630 => x"01",
          5631 => x"01",
          5632 => x"02",
          5633 => x"00",
          5634 => x"00",
        others => X"00"
    );

    shared variable RAM4 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"80",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"09",
             9 => x"83",
            10 => x"00",
            11 => x"00",
            12 => x"73",
            13 => x"83",
            14 => x"ff",
            15 => x"00",
            16 => x"73",
            17 => x"06",
            18 => x"00",
            19 => x"00",
            20 => x"53",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"72",
            26 => x"06",
            27 => x"00",
            28 => x"53",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"04",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"0b",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"2a",
            49 => x"05",
            50 => x"00",
            51 => x"00",
            52 => x"83",
            53 => x"2b",
            54 => x"51",
            55 => x"00",
            56 => x"70",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"70",
            61 => x"06",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"51",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"06",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"09",
            77 => x"2a",
            78 => x"00",
            79 => x"00",
            80 => x"b7",
            81 => x"08",
            82 => x"00",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"88",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"88",
            91 => x"00",
            92 => x"0a",
            93 => x"06",
            94 => x"06",
            95 => x"00",
            96 => x"0a",
            97 => x"71",
            98 => x"05",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"52",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"51",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"8c",
           134 => x"04",
           135 => x"0b",
           136 => x"8c",
           137 => x"04",
           138 => x"0b",
           139 => x"8d",
           140 => x"04",
           141 => x"0b",
           142 => x"8d",
           143 => x"04",
           144 => x"0b",
           145 => x"8e",
           146 => x"04",
           147 => x"0b",
           148 => x"8e",
           149 => x"04",
           150 => x"0b",
           151 => x"8f",
           152 => x"04",
           153 => x"0b",
           154 => x"8f",
           155 => x"04",
           156 => x"0b",
           157 => x"90",
           158 => x"04",
           159 => x"0b",
           160 => x"90",
           161 => x"04",
           162 => x"0b",
           163 => x"91",
           164 => x"04",
           165 => x"0b",
           166 => x"91",
           167 => x"04",
           168 => x"0b",
           169 => x"92",
           170 => x"04",
           171 => x"0b",
           172 => x"93",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"a4",
           193 => x"a4",
           194 => x"e0",
           195 => x"a4",
           196 => x"e0",
           197 => x"a4",
           198 => x"e0",
           199 => x"a4",
           200 => x"e0",
           201 => x"a4",
           202 => x"e0",
           203 => x"a4",
           204 => x"e0",
           205 => x"e0",
           206 => x"82",
           207 => x"82",
           208 => x"04",
           209 => x"82",
           210 => x"04",
           211 => x"82",
           212 => x"04",
           213 => x"82",
           214 => x"04",
           215 => x"2d",
           216 => x"90",
           217 => x"f6",
           218 => x"80",
           219 => x"80",
           220 => x"c0",
           221 => x"80",
           222 => x"80",
           223 => x"0c",
           224 => x"08",
           225 => x"a4",
           226 => x"a4",
           227 => x"e0",
           228 => x"e0",
           229 => x"82",
           230 => x"82",
           231 => x"04",
           232 => x"2d",
           233 => x"90",
           234 => x"e5",
           235 => x"80",
           236 => x"91",
           237 => x"c0",
           238 => x"82",
           239 => x"80",
           240 => x"0c",
           241 => x"08",
           242 => x"a4",
           243 => x"a4",
           244 => x"e0",
           245 => x"e0",
           246 => x"82",
           247 => x"82",
           248 => x"04",
           249 => x"2d",
           250 => x"90",
           251 => x"97",
           252 => x"80",
           253 => x"8e",
           254 => x"c0",
           255 => x"82",
           256 => x"80",
           257 => x"0c",
           258 => x"08",
           259 => x"a4",
           260 => x"a4",
           261 => x"e0",
           262 => x"e0",
           263 => x"82",
           264 => x"82",
           265 => x"04",
           266 => x"2d",
           267 => x"90",
           268 => x"8e",
           269 => x"80",
           270 => x"9f",
           271 => x"c0",
           272 => x"82",
           273 => x"80",
           274 => x"0c",
           275 => x"08",
           276 => x"a4",
           277 => x"a4",
           278 => x"e0",
           279 => x"e0",
           280 => x"82",
           281 => x"82",
           282 => x"04",
           283 => x"2d",
           284 => x"90",
           285 => x"f5",
           286 => x"80",
           287 => x"b8",
           288 => x"c0",
           289 => x"80",
           290 => x"80",
           291 => x"0c",
           292 => x"08",
           293 => x"a4",
           294 => x"a4",
           295 => x"e0",
           296 => x"e0",
           297 => x"82",
           298 => x"82",
           299 => x"04",
           300 => x"2d",
           301 => x"90",
           302 => x"bf",
           303 => x"80",
           304 => x"ac",
           305 => x"c0",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"00",
           311 => x"06",
           312 => x"10",
           313 => x"51",
           314 => x"ff",
           315 => x"52",
           316 => x"38",
           317 => x"98",
           318 => x"80",
           319 => x"0b",
           320 => x"80",
           321 => x"08",
           322 => x"0d",
           323 => x"82",
           324 => x"e0",
           325 => x"e0",
           326 => x"fb",
           327 => x"82",
           328 => x"08",
           329 => x"f8",
           330 => x"51",
           331 => x"0c",
           332 => x"e0",
           333 => x"a4",
           334 => x"70",
           335 => x"51",
           336 => x"e0",
           337 => x"38",
           338 => x"08",
           339 => x"e0",
           340 => x"82",
           341 => x"0b",
           342 => x"82",
           343 => x"e0",
           344 => x"a4",
           345 => x"f6",
           346 => x"8c",
           347 => x"e0",
           348 => x"90",
           349 => x"e0",
           350 => x"e0",
           351 => x"09",
           352 => x"e0",
           353 => x"39",
           354 => x"82",
           355 => x"53",
           356 => x"8c",
           357 => x"08",
           358 => x"fc",
           359 => x"08",
           360 => x"e0",
           361 => x"72",
           362 => x"08",
           363 => x"0c",
           364 => x"08",
           365 => x"82",
           366 => x"08",
           367 => x"0d",
           368 => x"05",
           369 => x"08",
           370 => x"fe",
           371 => x"05",
           372 => x"70",
           373 => x"82",
           374 => x"82",
           375 => x"82",
           376 => x"51",
           377 => x"08",
           378 => x"0c",
           379 => x"82",
           380 => x"51",
           381 => x"08",
           382 => x"0c",
           383 => x"0c",
           384 => x"e0",
           385 => x"a4",
           386 => x"08",
           387 => x"fc",
           388 => x"8c",
           389 => x"88",
           390 => x"e0",
           391 => x"f8",
           392 => x"05",
           393 => x"54",
           394 => x"04",
           395 => x"a4",
           396 => x"e0",
           397 => x"a4",
           398 => x"8c",
           399 => x"05",
           400 => x"70",
           401 => x"51",
           402 => x"ff",
           403 => x"0c",
           404 => x"8c",
           405 => x"82",
           406 => x"81",
           407 => x"fa",
           408 => x"08",
           409 => x"05",
           410 => x"22",
           411 => x"2e",
           412 => x"f8",
           413 => x"fc",
           414 => x"33",
           415 => x"82",
           416 => x"72",
           417 => x"38",
           418 => x"70",
           419 => x"53",
           420 => x"e4",
           421 => x"32",
           422 => x"72",
           423 => x"08",
           424 => x"51",
           425 => x"05",
           426 => x"08",
           427 => x"98",
           428 => x"73",
           429 => x"53",
           430 => x"34",
           431 => x"54",
           432 => x"70",
           433 => x"82",
           434 => x"e0",
           435 => x"2b",
           436 => x"80",
           437 => x"e0",
           438 => x"a4",
           439 => x"70",
           440 => x"db",
           441 => x"33",
           442 => x"90",
           443 => x"51",
           444 => x"05",
           445 => x"08",
           446 => x"81",
           447 => x"9d",
           448 => x"33",
           449 => x"51",
           450 => x"e0",
           451 => x"a4",
           452 => x"e0",
           453 => x"e0",
           454 => x"26",
           455 => x"c4",
           456 => x"dc",
           457 => x"72",
           458 => x"22",
           459 => x"e0",
           460 => x"a4",
           461 => x"51",
           462 => x"05",
           463 => x"08",
           464 => x"51",
           465 => x"05",
           466 => x"08",
           467 => x"51",
           468 => x"05",
           469 => x"08",
           470 => x"53",
           471 => x"23",
           472 => x"05",
           473 => x"08",
           474 => x"53",
           475 => x"23",
           476 => x"a4",
           477 => x"08",
           478 => x"72",
           479 => x"80",
           480 => x"05",
           481 => x"08",
           482 => x"90",
           483 => x"08",
           484 => x"72",
           485 => x"82",
           486 => x"11",
           487 => x"ec",
           488 => x"a4",
           489 => x"08",
           490 => x"a4",
           491 => x"e0",
           492 => x"a4",
           493 => x"70",
           494 => x"80",
           495 => x"e8",
           496 => x"98",
           497 => x"05",
           498 => x"e0",
           499 => x"08",
           500 => x"a4",
           501 => x"3f",
           502 => x"e0",
           503 => x"a4",
           504 => x"a4",
           505 => x"54",
           506 => x"05",
           507 => x"08",
           508 => x"90",
           509 => x"08",
           510 => x"a4",
           511 => x"08",
           512 => x"81",
           513 => x"2e",
           514 => x"05",
           515 => x"2c",
           516 => x"08",
           517 => x"98",
           518 => x"f4",
           519 => x"08",
           520 => x"82",
           521 => x"a4",
           522 => x"08",
           523 => x"08",
           524 => x"54",
           525 => x"23",
           526 => x"e4",
           527 => x"06",
           528 => x"38",
           529 => x"82",
           530 => x"05",
           531 => x"70",
           532 => x"0c",
           533 => x"90",
           534 => x"05",
           535 => x"90",
           536 => x"08",
           537 => x"08",
           538 => x"fc",
           539 => x"05",
           540 => x"a4",
           541 => x"51",
           542 => x"05",
           543 => x"08",
           544 => x"0c",
           545 => x"70",
           546 => x"e0",
           547 => x"39",
           548 => x"05",
           549 => x"e4",
           550 => x"53",
           551 => x"23",
           552 => x"f8",
           553 => x"08",
           554 => x"e4",
           555 => x"06",
           556 => x"38",
           557 => x"82",
           558 => x"05",
           559 => x"70",
           560 => x"0c",
           561 => x"90",
           562 => x"05",
           563 => x"90",
           564 => x"08",
           565 => x"08",
           566 => x"fc",
           567 => x"05",
           568 => x"82",
           569 => x"e0",
           570 => x"05",
           571 => x"08",
           572 => x"82",
           573 => x"55",
           574 => x"3f",
           575 => x"34",
           576 => x"82",
           577 => x"e0",
           578 => x"51",
           579 => x"e0",
           580 => x"33",
           581 => x"33",
           582 => x"72",
           583 => x"97",
           584 => x"08",
           585 => x"72",
           586 => x"82",
           587 => x"82",
           588 => x"34",
           589 => x"81",
           590 => x"0c",
           591 => x"70",
           592 => x"08",
           593 => x"98",
           594 => x"05",
           595 => x"05",
           596 => x"39",
           597 => x"82",
           598 => x"70",
           599 => x"a4",
           600 => x"08",
           601 => x"53",
           602 => x"a4",
           603 => x"53",
           604 => x"23",
           605 => x"70",
           606 => x"53",
           607 => x"e0",
           608 => x"2b",
           609 => x"82",
           610 => x"2c",
           611 => x"82",
           612 => x"53",
           613 => x"38",
           614 => x"fe",
           615 => x"c8",
           616 => x"08",
           617 => x"82",
           618 => x"e0",
           619 => x"a4",
           620 => x"08",
           621 => x"81",
           622 => x"80",
           623 => x"05",
           624 => x"82",
           625 => x"51",
           626 => x"82",
           627 => x"f7",
           628 => x"08",
           629 => x"a4",
           630 => x"a4",
           631 => x"54",
           632 => x"05",
           633 => x"22",
           634 => x"51",
           635 => x"e0",
           636 => x"2b",
           637 => x"88",
           638 => x"54",
           639 => x"70",
           640 => x"a4",
           641 => x"e0",
           642 => x"2b",
           643 => x"88",
           644 => x"54",
           645 => x"70",
           646 => x"a4",
           647 => x"08",
           648 => x"51",
           649 => x"08",
           650 => x"72",
           651 => x"73",
           652 => x"80",
           653 => x"08",
           654 => x"ee",
           655 => x"e4",
           656 => x"06",
           657 => x"38",
           658 => x"52",
           659 => x"39",
           660 => x"70",
           661 => x"53",
           662 => x"a4",
           663 => x"8a",
           664 => x"08",
           665 => x"81",
           666 => x"8e",
           667 => x"08",
           668 => x"e0",
           669 => x"2a",
           670 => x"80",
           671 => x"88",
           672 => x"3f",
           673 => x"53",
           674 => x"38",
           675 => x"52",
           676 => x"51",
           677 => x"e4",
           678 => x"06",
           679 => x"38",
           680 => x"ff",
           681 => x"08",
           682 => x"90",
           683 => x"38",
           684 => x"52",
           685 => x"82",
           686 => x"83",
           687 => x"72",
           688 => x"08",
           689 => x"72",
           690 => x"73",
           691 => x"80",
           692 => x"08",
           693 => x"b6",
           694 => x"e4",
           695 => x"06",
           696 => x"e0",
           697 => x"54",
           698 => x"05",
           699 => x"51",
           700 => x"e0",
           701 => x"51",
           702 => x"a4",
           703 => x"e3",
           704 => x"e0",
           705 => x"e0",
           706 => x"ce",
           707 => x"08",
           708 => x"2e",
           709 => x"e0",
           710 => x"51",
           711 => x"05",
           712 => x"72",
           713 => x"82",
           714 => x"82",
           715 => x"33",
           716 => x"08",
           717 => x"05",
           718 => x"39",
           719 => x"53",
           720 => x"80",
           721 => x"05",
           722 => x"e0",
           723 => x"ff",
           724 => x"2e",
           725 => x"88",
           726 => x"fc",
           727 => x"a6",
           728 => x"08",
           729 => x"05",
           730 => x"08",
           731 => x"a9",
           732 => x"08",
           733 => x"08",
           734 => x"05",
           735 => x"08",
           736 => x"cc",
           737 => x"22",
           738 => x"51",
           739 => x"82",
           740 => x"11",
           741 => x"ec",
           742 => x"2c",
           743 => x"82",
           744 => x"a0",
           745 => x"e0",
           746 => x"e0",
           747 => x"86",
           748 => x"e4",
           749 => x"a4",
           750 => x"2e",
           751 => x"82",
           752 => x"0b",
           753 => x"80",
           754 => x"34",
           755 => x"05",
           756 => x"08",
           757 => x"08",
           758 => x"e9",
           759 => x"05",
           760 => x"a4",
           761 => x"e0",
           762 => x"98",
           763 => x"0c",
           764 => x"e0",
           765 => x"f8",
           766 => x"05",
           767 => x"05",
           768 => x"98",
           769 => x"85",
           770 => x"82",
           771 => x"0c",
           772 => x"a4",
           773 => x"08",
           774 => x"81",
           775 => x"51",
           776 => x"0b",
           777 => x"81",
           778 => x"05",
           779 => x"08",
           780 => x"a4",
           781 => x"e0",
           782 => x"ff",
           783 => x"82",
           784 => x"53",
           785 => x"52",
           786 => x"82",
           787 => x"ff",
           788 => x"08",
           789 => x"fb",
           790 => x"53",
           791 => x"2d",
           792 => x"2e",
           793 => x"08",
           794 => x"f8",
           795 => x"f4",
           796 => x"f4",
           797 => x"3d",
           798 => x"e0",
           799 => x"fb",
           800 => x"08",
           801 => x"8c",
           802 => x"2a",
           803 => x"51",
           804 => x"38",
           805 => x"05",
           806 => x"08",
           807 => x"e0",
           808 => x"82",
           809 => x"72",
           810 => x"72",
           811 => x"b6",
           812 => x"08",
           813 => x"53",
           814 => x"52",
           815 => x"82",
           816 => x"ff",
           817 => x"08",
           818 => x"e0",
           819 => x"e0",
           820 => x"e0",
           821 => x"98",
           822 => x"0c",
           823 => x"e0",
           824 => x"fc",
           825 => x"05",
           826 => x"08",
           827 => x"3d",
           828 => x"e0",
           829 => x"fb",
           830 => x"05",
           831 => x"70",
           832 => x"51",
           833 => x"ff",
           834 => x"0c",
           835 => x"8c",
           836 => x"2a",
           837 => x"72",
           838 => x"a4",
           839 => x"08",
           840 => x"08",
           841 => x"e0",
           842 => x"70",
           843 => x"52",
           844 => x"08",
           845 => x"08",
           846 => x"05",
           847 => x"88",
           848 => x"fc",
           849 => x"82",
           850 => x"e0",
           851 => x"e0",
           852 => x"ff",
           853 => x"54",
           854 => x"72",
           855 => x"05",
           856 => x"12",
           857 => x"08",
           858 => x"0c",
           859 => x"e0",
           860 => x"a4",
           861 => x"0c",
           862 => x"04",
           863 => x"a4",
           864 => x"08",
           865 => x"81",
           866 => x"52",
           867 => x"82",
           868 => x"94",
           869 => x"08",
           870 => x"81",
           871 => x"2e",
           872 => x"88",
           873 => x"05",
           874 => x"ff",
           875 => x"34",
           876 => x"8c",
           877 => x"82",
           878 => x"11",
           879 => x"05",
           880 => x"82",
           881 => x"11",
           882 => x"51",
           883 => x"d7",
           884 => x"08",
           885 => x"08",
           886 => x"a4",
           887 => x"e0",
           888 => x"a4",
           889 => x"12",
           890 => x"85",
           891 => x"08",
           892 => x"e0",
           893 => x"81",
           894 => x"82",
           895 => x"e0",
           896 => x"11",
           897 => x"98",
           898 => x"05",
           899 => x"05",
           900 => x"e0",
           901 => x"a4",
           902 => x"08",
           903 => x"e0",
           904 => x"e0",
           905 => x"09",
           906 => x"08",
           907 => x"82",
           908 => x"39",
           909 => x"a0",
           910 => x"ec",
           911 => x"05",
           912 => x"05",
           913 => x"e0",
           914 => x"82",
           915 => x"11",
           916 => x"e0",
           917 => x"ff",
           918 => x"05",
           919 => x"08",
           920 => x"89",
           921 => x"82",
           922 => x"0c",
           923 => x"88",
           924 => x"05",
           925 => x"08",
           926 => x"82",
           927 => x"2e",
           928 => x"f8",
           929 => x"05",
           930 => x"a4",
           931 => x"08",
           932 => x"a4",
           933 => x"90",
           934 => x"08",
           935 => x"05",
           936 => x"82",
           937 => x"e0",
           938 => x"e0",
           939 => x"a4",
           940 => x"e0",
           941 => x"a4",
           942 => x"e0",
           943 => x"a4",
           944 => x"9c",
           945 => x"08",
           946 => x"05",
           947 => x"08",
           948 => x"05",
           949 => x"08",
           950 => x"53",
           951 => x"39",
           952 => x"81",
           953 => x"0c",
           954 => x"ff",
           955 => x"0c",
           956 => x"80",
           957 => x"f8",
           958 => x"a4",
           959 => x"e0",
           960 => x"a4",
           961 => x"71",
           962 => x"08",
           963 => x"05",
           964 => x"08",
           965 => x"0c",
           966 => x"0c",
           967 => x"e0",
           968 => x"a4",
           969 => x"08",
           970 => x"fc",
           971 => x"a4",
           972 => x"e0",
           973 => x"ff",
           974 => x"38",
           975 => x"05",
           976 => x"fc",
           977 => x"05",
           978 => x"08",
           979 => x"84",
           980 => x"82",
           981 => x"0c",
           982 => x"88",
           983 => x"05",
           984 => x"08",
           985 => x"8c",
           986 => x"08",
           987 => x"fc",
           988 => x"82",
           989 => x"05",
           990 => x"70",
           991 => x"84",
           992 => x"08",
           993 => x"0c",
           994 => x"0c",
           995 => x"e0",
           996 => x"a4",
           997 => x"08",
           998 => x"8c",
           999 => x"05",
          1000 => x"08",
          1001 => x"a4",
          1002 => x"e0",
          1003 => x"a4",
          1004 => x"e0",
          1005 => x"a4",
          1006 => x"38",
          1007 => x"51",
          1008 => x"05",
          1009 => x"f8",
          1010 => x"05",
          1011 => x"e0",
          1012 => x"82",
          1013 => x"ad",
          1014 => x"08",
          1015 => x"3d",
          1016 => x"e0",
          1017 => x"fd",
          1018 => x"05",
          1019 => x"e0",
          1020 => x"33",
          1021 => x"81",
          1022 => x"0c",
          1023 => x"70",
          1024 => x"54",
          1025 => x"ce",
          1026 => x"08",
          1027 => x"88",
          1028 => x"08",
          1029 => x"51",
          1030 => x"e0",
          1031 => x"39",
          1032 => x"ff",
          1033 => x"0c",
          1034 => x"80",
          1035 => x"e0",
          1036 => x"80",
          1037 => x"05",
          1038 => x"38",
          1039 => x"05",
          1040 => x"08",
          1041 => x"a4",
          1042 => x"08",
          1043 => x"70",
          1044 => x"08",
          1045 => x"a4",
          1046 => x"e0",
          1047 => x"72",
          1048 => x"fc",
          1049 => x"8a",
          1050 => x"fc",
          1051 => x"05",
          1052 => x"0d",
          1053 => x"a4",
          1054 => x"3d",
          1055 => x"08",
          1056 => x"08",
          1057 => x"08",
          1058 => x"0c",
          1059 => x"81",
          1060 => x"f7",
          1061 => x"e0",
          1062 => x"e0",
          1063 => x"80",
          1064 => x"0c",
          1065 => x"05",
          1066 => x"08",
          1067 => x"a4",
          1068 => x"a4",
          1069 => x"a4",
          1070 => x"3f",
          1071 => x"a4",
          1072 => x"a4",
          1073 => x"0c",
          1074 => x"04",
          1075 => x"a4",
          1076 => x"08",
          1077 => x"f8",
          1078 => x"05",
          1079 => x"a4",
          1080 => x"82",
          1081 => x"71",
          1082 => x"08",
          1083 => x"05",
          1084 => x"70",
          1085 => x"08",
          1086 => x"a4",
          1087 => x"08",
          1088 => x"ff",
          1089 => x"05",
          1090 => x"f8",
          1091 => x"05",
          1092 => x"08",
          1093 => x"05",
          1094 => x"05",
          1095 => x"0d",
          1096 => x"a4",
          1097 => x"3d",
          1098 => x"08",
          1099 => x"82",
          1100 => x"2e",
          1101 => x"90",
          1102 => x"08",
          1103 => x"90",
          1104 => x"08",
          1105 => x"90",
          1106 => x"e0",
          1107 => x"82",
          1108 => x"52",
          1109 => x"fc",
          1110 => x"08",
          1111 => x"e0",
          1112 => x"e0",
          1113 => x"e0",
          1114 => x"02",
          1115 => x"82",
          1116 => x"82",
          1117 => x"93",
          1118 => x"e0",
          1119 => x"e0",
          1120 => x"02",
          1121 => x"a0",
          1122 => x"0c",
          1123 => x"80",
          1124 => x"8c",
          1125 => x"e0",
          1126 => x"e4",
          1127 => x"a4",
          1128 => x"08",
          1129 => x"88",
          1130 => x"e0",
          1131 => x"c9",
          1132 => x"a4",
          1133 => x"e0",
          1134 => x"39",
          1135 => x"82",
          1136 => x"82",
          1137 => x"e0",
          1138 => x"a4",
          1139 => x"08",
          1140 => x"82",
          1141 => x"8d",
          1142 => x"e8",
          1143 => x"a4",
          1144 => x"71",
          1145 => x"2e",
          1146 => x"a4",
          1147 => x"a4",
          1148 => x"39",
          1149 => x"81",
          1150 => x"0c",
          1151 => x"82",
          1152 => x"82",
          1153 => x"e0",
          1154 => x"a4",
          1155 => x"a4",
          1156 => x"e0",
          1157 => x"0b",
          1158 => x"82",
          1159 => x"2e",
          1160 => x"f4",
          1161 => x"fc",
          1162 => x"08",
          1163 => x"07",
          1164 => x"82",
          1165 => x"70",
          1166 => x"07",
          1167 => x"82",
          1168 => x"e0",
          1169 => x"11",
          1170 => x"ff",
          1171 => x"08",
          1172 => x"ec",
          1173 => x"08",
          1174 => x"8c",
          1175 => x"05",
          1176 => x"05",
          1177 => x"f4",
          1178 => x"05",
          1179 => x"f8",
          1180 => x"51",
          1181 => x"a4",
          1182 => x"e0",
          1183 => x"e0",
          1184 => x"a4",
          1185 => x"a4",
          1186 => x"e0",
          1187 => x"98",
          1188 => x"0c",
          1189 => x"e0",
          1190 => x"a4",
          1191 => x"08",
          1192 => x"fc",
          1193 => x"70",
          1194 => x"08",
          1195 => x"82",
          1196 => x"e0",
          1197 => x"a4",
          1198 => x"e0",
          1199 => x"e0",
          1200 => x"82",
          1201 => x"e0",
          1202 => x"a4",
          1203 => x"08",
          1204 => x"51",
          1205 => x"e0",
          1206 => x"80",
          1207 => x"0c",
          1208 => x"82",
          1209 => x"0b",
          1210 => x"31",
          1211 => x"71",
          1212 => x"0c",
          1213 => x"82",
          1214 => x"82",
          1215 => x"e0",
          1216 => x"06",
          1217 => x"82",
          1218 => x"39",
          1219 => x"05",
          1220 => x"08",
          1221 => x"84",
          1222 => x"08",
          1223 => x"08",
          1224 => x"05",
          1225 => x"08",
          1226 => x"05",
          1227 => x"82",
          1228 => x"06",
          1229 => x"82",
          1230 => x"39",
          1231 => x"05",
          1232 => x"08",
          1233 => x"82",
          1234 => x"08",
          1235 => x"08",
          1236 => x"05",
          1237 => x"08",
          1238 => x"05",
          1239 => x"82",
          1240 => x"08",
          1241 => x"08",
          1242 => x"06",
          1243 => x"a4",
          1244 => x"82",
          1245 => x"51",
          1246 => x"82",
          1247 => x"08",
          1248 => x"0d",
          1249 => x"52",
          1250 => x"51",
          1251 => x"70",
          1252 => x"29",
          1253 => x"71",
          1254 => x"51",
          1255 => x"0c",
          1256 => x"e0",
          1257 => x"a4",
          1258 => x"a4",
          1259 => x"82",
          1260 => x"0c",
          1261 => x"0c",
          1262 => x"e0",
          1263 => x"82",
          1264 => x"e0",
          1265 => x"9b",
          1266 => x"08",
          1267 => x"08",
          1268 => x"0c",
          1269 => x"fc",
          1270 => x"05",
          1271 => x"08",
          1272 => x"08",
          1273 => x"82",
          1274 => x"e4",
          1275 => x"08",
          1276 => x"e0",
          1277 => x"a4",
          1278 => x"a4",
          1279 => x"08",
          1280 => x"f8",
          1281 => x"05",
          1282 => x"a4",
          1283 => x"82",
          1284 => x"82",
          1285 => x"82",
          1286 => x"05",
          1287 => x"a4",
          1288 => x"06",
          1289 => x"08",
          1290 => x"e0",
          1291 => x"82",
          1292 => x"e0",
          1293 => x"a4",
          1294 => x"a4",
          1295 => x"08",
          1296 => x"f8",
          1297 => x"88",
          1298 => x"08",
          1299 => x"e0",
          1300 => x"a4",
          1301 => x"ab",
          1302 => x"08",
          1303 => x"08",
          1304 => x"05",
          1305 => x"e0",
          1306 => x"a4",
          1307 => x"e0",
          1308 => x"e0",
          1309 => x"a4",
          1310 => x"08",
          1311 => x"e0",
          1312 => x"71",
          1313 => x"05",
          1314 => x"08",
          1315 => x"05",
          1316 => x"08",
          1317 => x"06",
          1318 => x"71",
          1319 => x"0c",
          1320 => x"ff",
          1321 => x"0c",
          1322 => x"53",
          1323 => x"f4",
          1324 => x"e8",
          1325 => x"e8",
          1326 => x"3d",
          1327 => x"e0",
          1328 => x"fb",
          1329 => x"08",
          1330 => x"88",
          1331 => x"05",
          1332 => x"05",
          1333 => x"08",
          1334 => x"2c",
          1335 => x"82",
          1336 => x"e0",
          1337 => x"82",
          1338 => x"82",
          1339 => x"e0",
          1340 => x"a4",
          1341 => x"e0",
          1342 => x"e0",
          1343 => x"a4",
          1344 => x"08",
          1345 => x"08",
          1346 => x"8c",
          1347 => x"88",
          1348 => x"3f",
          1349 => x"a4",
          1350 => x"e0",
          1351 => x"82",
          1352 => x"3d",
          1353 => x"e0",
          1354 => x"f7",
          1355 => x"08",
          1356 => x"8c",
          1357 => x"e0",
          1358 => x"51",
          1359 => x"a4",
          1360 => x"06",
          1361 => x"91",
          1362 => x"08",
          1363 => x"ce",
          1364 => x"33",
          1365 => x"a4",
          1366 => x"f0",
          1367 => x"05",
          1368 => x"70",
          1369 => x"a4",
          1370 => x"08",
          1371 => x"09",
          1372 => x"a4",
          1373 => x"05",
          1374 => x"33",
          1375 => x"82",
          1376 => x"e0",
          1377 => x"a4",
          1378 => x"b6",
          1379 => x"08",
          1380 => x"39",
          1381 => x"05",
          1382 => x"08",
          1383 => x"08",
          1384 => x"08",
          1385 => x"0b",
          1386 => x"82",
          1387 => x"08",
          1388 => x"53",
          1389 => x"05",
          1390 => x"08",
          1391 => x"8d",
          1392 => x"ec",
          1393 => x"a4",
          1394 => x"27",
          1395 => x"05",
          1396 => x"8d",
          1397 => x"ec",
          1398 => x"82",
          1399 => x"39",
          1400 => x"53",
          1401 => x"a4",
          1402 => x"26",
          1403 => x"e0",
          1404 => x"39",
          1405 => x"05",
          1406 => x"fc",
          1407 => x"05",
          1408 => x"38",
          1409 => x"53",
          1410 => x"e0",
          1411 => x"51",
          1412 => x"05",
          1413 => x"33",
          1414 => x"a4",
          1415 => x"08",
          1416 => x"ad",
          1417 => x"33",
          1418 => x"a4",
          1419 => x"08",
          1420 => x"8d",
          1421 => x"ec",
          1422 => x"a4",
          1423 => x"08",
          1424 => x"26",
          1425 => x"08",
          1426 => x"e0",
          1427 => x"e0",
          1428 => x"e0",
          1429 => x"82",
          1430 => x"e0",
          1431 => x"81",
          1432 => x"52",
          1433 => x"08",
          1434 => x"e0",
          1435 => x"80",
          1436 => x"fc",
          1437 => x"fc",
          1438 => x"05",
          1439 => x"08",
          1440 => x"a4",
          1441 => x"08",
          1442 => x"8b",
          1443 => x"82",
          1444 => x"0c",
          1445 => x"a4",
          1446 => x"08",
          1447 => x"82",
          1448 => x"08",
          1449 => x"e0",
          1450 => x"ff",
          1451 => x"06",
          1452 => x"05",
          1453 => x"53",
          1454 => x"05",
          1455 => x"06",
          1456 => x"08",
          1457 => x"88",
          1458 => x"0c",
          1459 => x"e0",
          1460 => x"a4",
          1461 => x"2e",
          1462 => x"e0",
          1463 => x"81",
          1464 => x"72",
          1465 => x"34",
          1466 => x"82",
          1467 => x"e0",
          1468 => x"2e",
          1469 => x"05",
          1470 => x"cd",
          1471 => x"f4",
          1472 => x"05",
          1473 => x"70",
          1474 => x"a4",
          1475 => x"82",
          1476 => x"34",
          1477 => x"70",
          1478 => x"51",
          1479 => x"f8",
          1480 => x"a4",
          1481 => x"26",
          1482 => x"08",
          1483 => x"e0",
          1484 => x"73",
          1485 => x"f8",
          1486 => x"38",
          1487 => x"08",
          1488 => x"0b",
          1489 => x"b2",
          1490 => x"33",
          1491 => x"e0",
          1492 => x"b9",
          1493 => x"82",
          1494 => x"a5",
          1495 => x"f4",
          1496 => x"08",
          1497 => x"f8",
          1498 => x"cf",
          1499 => x"33",
          1500 => x"82",
          1501 => x"11",
          1502 => x"f8",
          1503 => x"05",
          1504 => x"e0",
          1505 => x"a4",
          1506 => x"27",
          1507 => x"05",
          1508 => x"e0",
          1509 => x"a4",
          1510 => x"26",
          1511 => x"08",
          1512 => x"e0",
          1513 => x"a4",
          1514 => x"74",
          1515 => x"a4",
          1516 => x"82",
          1517 => x"82",
          1518 => x"82",
          1519 => x"12",
          1520 => x"82",
          1521 => x"08",
          1522 => x"51",
          1523 => x"a4",
          1524 => x"82",
          1525 => x"72",
          1526 => x"08",
          1527 => x"08",
          1528 => x"8c",
          1529 => x"05",
          1530 => x"e0",
          1531 => x"a4",
          1532 => x"0c",
          1533 => x"04",
          1534 => x"56",
          1535 => x"38",
          1536 => x"16",
          1537 => x"54",
          1538 => x"38",
          1539 => x"76",
          1540 => x"08",
          1541 => x"98",
          1542 => x"53",
          1543 => x"82",
          1544 => x"33",
          1545 => x"81",
          1546 => x"98",
          1547 => x"82",
          1548 => x"81",
          1549 => x"ff",
          1550 => x"81",
          1551 => x"fc",
          1552 => x"e4",
          1553 => x"51",
          1554 => x"80",
          1555 => x"eb",
          1556 => x"39",
          1557 => x"82",
          1558 => x"be",
          1559 => x"ec",
          1560 => x"51",
          1561 => x"bb",
          1562 => x"82",
          1563 => x"f4",
          1564 => x"a3",
          1565 => x"82",
          1566 => x"cc",
          1567 => x"8b",
          1568 => x"82",
          1569 => x"3d",
          1570 => x"56",
          1571 => x"74",
          1572 => x"39",
          1573 => x"3f",
          1574 => x"e3",
          1575 => x"79",
          1576 => x"ff",
          1577 => x"ec",
          1578 => x"e3",
          1579 => x"30",
          1580 => x"59",
          1581 => x"83",
          1582 => x"81",
          1583 => x"81",
          1584 => x"3d",
          1585 => x"82",
          1586 => x"08",
          1587 => x"c0",
          1588 => x"59",
          1589 => x"53",
          1590 => x"3f",
          1591 => x"98",
          1592 => x"2e",
          1593 => x"59",
          1594 => x"81",
          1595 => x"07",
          1596 => x"72",
          1597 => x"2e",
          1598 => x"c0",
          1599 => x"92",
          1600 => x"0c",
          1601 => x"7c",
          1602 => x"59",
          1603 => x"51",
          1604 => x"a8",
          1605 => x"81",
          1606 => x"f8",
          1607 => x"98",
          1608 => x"82",
          1609 => x"04",
          1610 => x"0d",
          1611 => x"02",
          1612 => x"73",
          1613 => x"5e",
          1614 => x"82",
          1615 => x"88",
          1616 => x"58",
          1617 => x"39",
          1618 => x"7a",
          1619 => x"ec",
          1620 => x"e4",
          1621 => x"80",
          1622 => x"a0",
          1623 => x"19",
          1624 => x"22",
          1625 => x"bc",
          1626 => x"ff",
          1627 => x"c3",
          1628 => x"8e",
          1629 => x"51",
          1630 => x"c1",
          1631 => x"15",
          1632 => x"7a",
          1633 => x"c1",
          1634 => x"39",
          1635 => x"3f",
          1636 => x"52",
          1637 => x"39",
          1638 => x"3f",
          1639 => x"38",
          1640 => x"56",
          1641 => x"80",
          1642 => x"53",
          1643 => x"51",
          1644 => x"80",
          1645 => x"08",
          1646 => x"fc",
          1647 => x"81",
          1648 => x"f4",
          1649 => x"1c",
          1650 => x"82",
          1651 => x"2c",
          1652 => x"06",
          1653 => x"82",
          1654 => x"2c",
          1655 => x"32",
          1656 => x"07",
          1657 => x"57",
          1658 => x"2e",
          1659 => x"79",
          1660 => x"82",
          1661 => x"fc",
          1662 => x"8a",
          1663 => x"52",
          1664 => x"3f",
          1665 => x"3f",
          1666 => x"53",
          1667 => x"98",
          1668 => x"2e",
          1669 => x"0d",
          1670 => x"80",
          1671 => x"99",
          1672 => x"d4",
          1673 => x"81",
          1674 => x"80",
          1675 => x"3f",
          1676 => x"80",
          1677 => x"70",
          1678 => x"92",
          1679 => x"c2",
          1680 => x"98",
          1681 => x"06",
          1682 => x"81",
          1683 => x"51",
          1684 => x"3f",
          1685 => x"52",
          1686 => x"98",
          1687 => x"dc",
          1688 => x"85",
          1689 => x"80",
          1690 => x"3f",
          1691 => x"80",
          1692 => x"70",
          1693 => x"92",
          1694 => x"c3",
          1695 => x"97",
          1696 => x"06",
          1697 => x"81",
          1698 => x"51",
          1699 => x"3f",
          1700 => x"52",
          1701 => x"97",
          1702 => x"e4",
          1703 => x"f8",
          1704 => x"0d",
          1705 => x"70",
          1706 => x"d9",
          1707 => x"33",
          1708 => x"c4",
          1709 => x"8b",
          1710 => x"70",
          1711 => x"82",
          1712 => x"0b",
          1713 => x"db",
          1714 => x"81",
          1715 => x"74",
          1716 => x"82",
          1717 => x"82",
          1718 => x"91",
          1719 => x"e7",
          1720 => x"9c",
          1721 => x"54",
          1722 => x"38",
          1723 => x"51",
          1724 => x"98",
          1725 => x"0d",
          1726 => x"f7",
          1727 => x"80",
          1728 => x"81",
          1729 => x"81",
          1730 => x"53",
          1731 => x"f9",
          1732 => x"c4",
          1733 => x"98",
          1734 => x"ac",
          1735 => x"5e",
          1736 => x"3f",
          1737 => x"52",
          1738 => x"ff",
          1739 => x"e0",
          1740 => x"51",
          1741 => x"38",
          1742 => x"bd",
          1743 => x"90",
          1744 => x"78",
          1745 => x"39",
          1746 => x"78",
          1747 => x"bf",
          1748 => x"78",
          1749 => x"80",
          1750 => x"2e",
          1751 => x"89",
          1752 => x"83",
          1753 => x"24",
          1754 => x"f1",
          1755 => x"2e",
          1756 => x"3d",
          1757 => x"51",
          1758 => x"80",
          1759 => x"fc",
          1760 => x"97",
          1761 => x"fe",
          1762 => x"53",
          1763 => x"82",
          1764 => x"98",
          1765 => x"a5",
          1766 => x"7b",
          1767 => x"7a",
          1768 => x"26",
          1769 => x"ff",
          1770 => x"eb",
          1771 => x"2e",
          1772 => x"11",
          1773 => x"3f",
          1774 => x"c8",
          1775 => x"ff",
          1776 => x"e0",
          1777 => x"82",
          1778 => x"64",
          1779 => x"62",
          1780 => x"79",
          1781 => x"b5",
          1782 => x"05",
          1783 => x"08",
          1784 => x"fe",
          1785 => x"ea",
          1786 => x"2e",
          1787 => x"11",
          1788 => x"3f",
          1789 => x"d0",
          1790 => x"94",
          1791 => x"38",
          1792 => x"5b",
          1793 => x"7a",
          1794 => x"c5",
          1795 => x"1a",
          1796 => x"8a",
          1797 => x"b5",
          1798 => x"05",
          1799 => x"08",
          1800 => x"59",
          1801 => x"b4",
          1802 => x"fd",
          1803 => x"82",
          1804 => x"de",
          1805 => x"38",
          1806 => x"82",
          1807 => x"88",
          1808 => x"39",
          1809 => x"2e",
          1810 => x"89",
          1811 => x"05",
          1812 => x"ff",
          1813 => x"e0",
          1814 => x"fc",
          1815 => x"82",
          1816 => x"82",
          1817 => x"88",
          1818 => x"39",
          1819 => x"2e",
          1820 => x"aa",
          1821 => x"80",
          1822 => x"44",
          1823 => x"78",
          1824 => x"08",
          1825 => x"88",
          1826 => x"53",
          1827 => x"82",
          1828 => x"80",
          1829 => x"38",
          1830 => x"70",
          1831 => x"51",
          1832 => x"38",
          1833 => x"82",
          1834 => x"80",
          1835 => x"64",
          1836 => x"51",
          1837 => x"11",
          1838 => x"3f",
          1839 => x"c0",
          1840 => x"ff",
          1841 => x"e0",
          1842 => x"59",
          1843 => x"64",
          1844 => x"11",
          1845 => x"3f",
          1846 => x"88",
          1847 => x"c5",
          1848 => x"fb",
          1849 => x"51",
          1850 => x"33",
          1851 => x"9f",
          1852 => x"fc",
          1853 => x"af",
          1854 => x"91",
          1855 => x"33",
          1856 => x"b1",
          1857 => x"87",
          1858 => x"f4",
          1859 => x"ae",
          1860 => x"f8",
          1861 => x"53",
          1862 => x"82",
          1863 => x"61",
          1864 => x"70",
          1865 => x"3d",
          1866 => x"51",
          1867 => x"df",
          1868 => x"54",
          1869 => x"9c",
          1870 => x"f8",
          1871 => x"79",
          1872 => x"f7",
          1873 => x"61",
          1874 => x"fe",
          1875 => x"df",
          1876 => x"2e",
          1877 => x"05",
          1878 => x"78",
          1879 => x"51",
          1880 => x"b5",
          1881 => x"05",
          1882 => x"08",
          1883 => x"fe",
          1884 => x"de",
          1885 => x"2e",
          1886 => x"61",
          1887 => x"11",
          1888 => x"3f",
          1889 => x"b0",
          1890 => x"c5",
          1891 => x"fb",
          1892 => x"51",
          1893 => x"33",
          1894 => x"9f",
          1895 => x"f0",
          1896 => x"86",
          1897 => x"8d",
          1898 => x"84",
          1899 => x"d4",
          1900 => x"39",
          1901 => x"84",
          1902 => x"98",
          1903 => x"52",
          1904 => x"3f",
          1905 => x"80",
          1906 => x"87",
          1907 => x"f5",
          1908 => x"51",
          1909 => x"2d",
          1910 => x"88",
          1911 => x"c6",
          1912 => x"f8",
          1913 => x"c7",
          1914 => x"39",
          1915 => x"3f",
          1916 => x"3f",
          1917 => x"78",
          1918 => x"52",
          1919 => x"98",
          1920 => x"2e",
          1921 => x"46",
          1922 => x"cc",
          1923 => x"06",
          1924 => x"38",
          1925 => x"3f",
          1926 => x"c1",
          1927 => x"38",
          1928 => x"2e",
          1929 => x"2e",
          1930 => x"f8",
          1931 => x"80",
          1932 => x"ff",
          1933 => x"b8",
          1934 => x"05",
          1935 => x"55",
          1936 => x"c7",
          1937 => x"51",
          1938 => x"54",
          1939 => x"3d",
          1940 => x"3f",
          1941 => x"57",
          1942 => x"80",
          1943 => x"3d",
          1944 => x"82",
          1945 => x"09",
          1946 => x"51",
          1947 => x"26",
          1948 => x"59",
          1949 => x"70",
          1950 => x"c3",
          1951 => x"07",
          1952 => x"09",
          1953 => x"51",
          1954 => x"f1",
          1955 => x"51",
          1956 => x"f5",
          1957 => x"34",
          1958 => x"55",
          1959 => x"93",
          1960 => x"75",
          1961 => x"73",
          1962 => x"98",
          1963 => x"9c",
          1964 => x"52",
          1965 => x"98",
          1966 => x"87",
          1967 => x"3f",
          1968 => x"0c",
          1969 => x"84",
          1970 => x"94",
          1971 => x"85",
          1972 => x"05",
          1973 => x"87",
          1974 => x"0c",
          1975 => x"3f",
          1976 => x"ff",
          1977 => x"ff",
          1978 => x"93",
          1979 => x"f0",
          1980 => x"76",
          1981 => x"54",
          1982 => x"33",
          1983 => x"86",
          1984 => x"33",
          1985 => x"86",
          1986 => x"52",
          1987 => x"38",
          1988 => x"33",
          1989 => x"81",
          1990 => x"ea",
          1991 => x"72",
          1992 => x"38",
          1993 => x"73",
          1994 => x"70",
          1995 => x"81",
          1996 => x"80",
          1997 => x"80",
          1998 => x"05",
          1999 => x"70",
          2000 => x"04",
          2001 => x"80",
          2002 => x"52",
          2003 => x"98",
          2004 => x"74",
          2005 => x"3d",
          2006 => x"11",
          2007 => x"70",
          2008 => x"33",
          2009 => x"26",
          2010 => x"83",
          2011 => x"85",
          2012 => x"26",
          2013 => x"85",
          2014 => x"88",
          2015 => x"e7",
          2016 => x"54",
          2017 => x"cc",
          2018 => x"0c",
          2019 => x"82",
          2020 => x"83",
          2021 => x"84",
          2022 => x"85",
          2023 => x"86",
          2024 => x"74",
          2025 => x"c0",
          2026 => x"98",
          2027 => x"98",
          2028 => x"0d",
          2029 => x"81",
          2030 => x"5e",
          2031 => x"08",
          2032 => x"98",
          2033 => x"87",
          2034 => x"1c",
          2035 => x"79",
          2036 => x"08",
          2037 => x"98",
          2038 => x"87",
          2039 => x"1c",
          2040 => x"ff",
          2041 => x"58",
          2042 => x"56",
          2043 => x"54",
          2044 => x"ff",
          2045 => x"94",
          2046 => x"3d",
          2047 => x"52",
          2048 => x"38",
          2049 => x"70",
          2050 => x"70",
          2051 => x"84",
          2052 => x"08",
          2053 => x"71",
          2054 => x"80",
          2055 => x"83",
          2056 => x"30",
          2057 => x"51",
          2058 => x"98",
          2059 => x"0d",
          2060 => x"53",
          2061 => x"98",
          2062 => x"07",
          2063 => x"25",
          2064 => x"85",
          2065 => x"9f",
          2066 => x"81",
          2067 => x"94",
          2068 => x"87",
          2069 => x"96",
          2070 => x"70",
          2071 => x"70",
          2072 => x"72",
          2073 => x"70",
          2074 => x"70",
          2075 => x"38",
          2076 => x"94",
          2077 => x"87",
          2078 => x"74",
          2079 => x"04",
          2080 => x"70",
          2081 => x"70",
          2082 => x"04",
          2083 => x"58",
          2084 => x"38",
          2085 => x"de",
          2086 => x"56",
          2087 => x"2e",
          2088 => x"72",
          2089 => x"55",
          2090 => x"73",
          2091 => x"72",
          2092 => x"06",
          2093 => x"73",
          2094 => x"72",
          2095 => x"53",
          2096 => x"2e",
          2097 => x"77",
          2098 => x"0c",
          2099 => x"79",
          2100 => x"06",
          2101 => x"fc",
          2102 => x"82",
          2103 => x"59",
          2104 => x"51",
          2105 => x"94",
          2106 => x"70",
          2107 => x"2e",
          2108 => x"06",
          2109 => x"32",
          2110 => x"2e",
          2111 => x"06",
          2112 => x"81",
          2113 => x"52",
          2114 => x"94",
          2115 => x"74",
          2116 => x"57",
          2117 => x"98",
          2118 => x"0d",
          2119 => x"06",
          2120 => x"72",
          2121 => x"94",
          2122 => x"81",
          2123 => x"e2",
          2124 => x"c0",
          2125 => x"38",
          2126 => x"70",
          2127 => x"51",
          2128 => x"82",
          2129 => x"e0",
          2130 => x"de",
          2131 => x"53",
          2132 => x"2e",
          2133 => x"71",
          2134 => x"51",
          2135 => x"a0",
          2136 => x"c0",
          2137 => x"38",
          2138 => x"70",
          2139 => x"51",
          2140 => x"0d",
          2141 => x"80",
          2142 => x"51",
          2143 => x"c0",
          2144 => x"87",
          2145 => x"0c",
          2146 => x"bc",
          2147 => x"de",
          2148 => x"82",
          2149 => x"08",
          2150 => x"ac",
          2151 => x"9e",
          2152 => x"c0",
          2153 => x"87",
          2154 => x"0c",
          2155 => x"dc",
          2156 => x"de",
          2157 => x"82",
          2158 => x"08",
          2159 => x"c0",
          2160 => x"87",
          2161 => x"0c",
          2162 => x"f4",
          2163 => x"80",
          2164 => x"84",
          2165 => x"80",
          2166 => x"de",
          2167 => x"90",
          2168 => x"52",
          2169 => x"52",
          2170 => x"87",
          2171 => x"0a",
          2172 => x"83",
          2173 => x"34",
          2174 => x"70",
          2175 => x"70",
          2176 => x"82",
          2177 => x"9e",
          2178 => x"51",
          2179 => x"81",
          2180 => x"0b",
          2181 => x"80",
          2182 => x"2e",
          2183 => x"fe",
          2184 => x"08",
          2185 => x"52",
          2186 => x"71",
          2187 => x"c0",
          2188 => x"06",
          2189 => x"38",
          2190 => x"80",
          2191 => x"81",
          2192 => x"80",
          2193 => x"df",
          2194 => x"90",
          2195 => x"52",
          2196 => x"52",
          2197 => x"87",
          2198 => x"06",
          2199 => x"38",
          2200 => x"87",
          2201 => x"06",
          2202 => x"82",
          2203 => x"9e",
          2204 => x"52",
          2205 => x"52",
          2206 => x"9e",
          2207 => x"84",
          2208 => x"86",
          2209 => x"08",
          2210 => x"80",
          2211 => x"df",
          2212 => x"70",
          2213 => x"88",
          2214 => x"0d",
          2215 => x"3f",
          2216 => x"2e",
          2217 => x"89",
          2218 => x"a5",
          2219 => x"73",
          2220 => x"08",
          2221 => x"82",
          2222 => x"82",
          2223 => x"94",
          2224 => x"d0",
          2225 => x"51",
          2226 => x"33",
          2227 => x"de",
          2228 => x"54",
          2229 => x"dc",
          2230 => x"80",
          2231 => x"82",
          2232 => x"c9",
          2233 => x"de",
          2234 => x"38",
          2235 => x"08",
          2236 => x"ff",
          2237 => x"54",
          2238 => x"84",
          2239 => x"88",
          2240 => x"73",
          2241 => x"33",
          2242 => x"f4",
          2243 => x"80",
          2244 => x"52",
          2245 => x"3f",
          2246 => x"2e",
          2247 => x"a3",
          2248 => x"73",
          2249 => x"51",
          2250 => x"33",
          2251 => x"ca",
          2252 => x"df",
          2253 => x"38",
          2254 => x"3f",
          2255 => x"2e",
          2256 => x"a3",
          2257 => x"a3",
          2258 => x"82",
          2259 => x"82",
          2260 => x"51",
          2261 => x"08",
          2262 => x"d4",
          2263 => x"d7",
          2264 => x"cc",
          2265 => x"de",
          2266 => x"75",
          2267 => x"98",
          2268 => x"31",
          2269 => x"82",
          2270 => x"82",
          2271 => x"aa",
          2272 => x"84",
          2273 => x"3f",
          2274 => x"29",
          2275 => x"98",
          2276 => x"85",
          2277 => x"73",
          2278 => x"08",
          2279 => x"ff",
          2280 => x"bd",
          2281 => x"54",
          2282 => x"90",
          2283 => x"ff",
          2284 => x"fe",
          2285 => x"05",
          2286 => x"84",
          2287 => x"08",
          2288 => x"82",
          2289 => x"cc",
          2290 => x"8b",
          2291 => x"82",
          2292 => x"84",
          2293 => x"04",
          2294 => x"04",
          2295 => x"84",
          2296 => x"2b",
          2297 => x"98",
          2298 => x"51",
          2299 => x"82",
          2300 => x"74",
          2301 => x"08",
          2302 => x"71",
          2303 => x"09",
          2304 => x"82",
          2305 => x"fb",
          2306 => x"05",
          2307 => x"80",
          2308 => x"52",
          2309 => x"fb",
          2310 => x"ae",
          2311 => x"51",
          2312 => x"05",
          2313 => x"06",
          2314 => x"b4",
          2315 => x"04",
          2316 => x"b7",
          2317 => x"33",
          2318 => x"82",
          2319 => x"59",
          2320 => x"38",
          2321 => x"e8",
          2322 => x"05",
          2323 => x"9d",
          2324 => x"0c",
          2325 => x"82",
          2326 => x"5a",
          2327 => x"78",
          2328 => x"82",
          2329 => x"82",
          2330 => x"55",
          2331 => x"82",
          2332 => x"38",
          2333 => x"2e",
          2334 => x"74",
          2335 => x"76",
          2336 => x"84",
          2337 => x"51",
          2338 => x"08",
          2339 => x"0d",
          2340 => x"53",
          2341 => x"2e",
          2342 => x"80",
          2343 => x"54",
          2344 => x"82",
          2345 => x"52",
          2346 => x"80",
          2347 => x"51",
          2348 => x"e4",
          2349 => x"0d",
          2350 => x"08",
          2351 => x"98",
          2352 => x"08",
          2353 => x"52",
          2354 => x"98",
          2355 => x"ff",
          2356 => x"55",
          2357 => x"9d",
          2358 => x"70",
          2359 => x"53",
          2360 => x"52",
          2361 => x"2e",
          2362 => x"3d",
          2363 => x"08",
          2364 => x"58",
          2365 => x"51",
          2366 => x"08",
          2367 => x"e4",
          2368 => x"3d",
          2369 => x"82",
          2370 => x"75",
          2371 => x"98",
          2372 => x"82",
          2373 => x"e0",
          2374 => x"55",
          2375 => x"70",
          2376 => x"78",
          2377 => x"38",
          2378 => x"53",
          2379 => x"98",
          2380 => x"e8",
          2381 => x"2e",
          2382 => x"79",
          2383 => x"ff",
          2384 => x"82",
          2385 => x"77",
          2386 => x"04",
          2387 => x"71",
          2388 => x"a0",
          2389 => x"33",
          2390 => x"38",
          2391 => x"56",
          2392 => x"06",
          2393 => x"80",
          2394 => x"05",
          2395 => x"3f",
          2396 => x"74",
          2397 => x"e0",
          2398 => x"33",
          2399 => x"82",
          2400 => x"3f",
          2401 => x"fc",
          2402 => x"3f",
          2403 => x"38",
          2404 => x"fd",
          2405 => x"ff",
          2406 => x"91",
          2407 => x"51",
          2408 => x"80",
          2409 => x"3d",
          2410 => x"08",
          2411 => x"5f",
          2412 => x"df",
          2413 => x"5b",
          2414 => x"e0",
          2415 => x"55",
          2416 => x"70",
          2417 => x"81",
          2418 => x"82",
          2419 => x"82",
          2420 => x"38",
          2421 => x"08",
          2422 => x"98",
          2423 => x"94",
          2424 => x"39",
          2425 => x"e4",
          2426 => x"70",
          2427 => x"e0",
          2428 => x"74",
          2429 => x"82",
          2430 => x"3f",
          2431 => x"82",
          2432 => x"e0",
          2433 => x"55",
          2434 => x"ff",
          2435 => x"81",
          2436 => x"93",
          2437 => x"ff",
          2438 => x"86",
          2439 => x"8c",
          2440 => x"84",
          2441 => x"80",
          2442 => x"08",
          2443 => x"78",
          2444 => x"06",
          2445 => x"70",
          2446 => x"98",
          2447 => x"05",
          2448 => x"70",
          2449 => x"51",
          2450 => x"56",
          2451 => x"74",
          2452 => x"29",
          2453 => x"51",
          2454 => x"76",
          2455 => x"3f",
          2456 => x"54",
          2457 => x"f7",
          2458 => x"81",
          2459 => x"70",
          2460 => x"51",
          2461 => x"53",
          2462 => x"82",
          2463 => x"73",
          2464 => x"80",
          2465 => x"74",
          2466 => x"70",
          2467 => x"98",
          2468 => x"70",
          2469 => x"5e",
          2470 => x"74",
          2471 => x"38",
          2472 => x"80",
          2473 => x"82",
          2474 => x"f7",
          2475 => x"78",
          2476 => x"54",
          2477 => x"84",
          2478 => x"08",
          2479 => x"7e",
          2480 => x"33",
          2481 => x"98",
          2482 => x"75",
          2483 => x"33",
          2484 => x"29",
          2485 => x"82",
          2486 => x"39",
          2487 => x"54",
          2488 => x"54",
          2489 => x"d8",
          2490 => x"81",
          2491 => x"82",
          2492 => x"29",
          2493 => x"82",
          2494 => x"74",
          2495 => x"08",
          2496 => x"ff",
          2497 => x"29",
          2498 => x"82",
          2499 => x"75",
          2500 => x"70",
          2501 => x"d8",
          2502 => x"25",
          2503 => x"52",
          2504 => x"81",
          2505 => x"70",
          2506 => x"51",
          2507 => x"ec",
          2508 => x"1b",
          2509 => x"82",
          2510 => x"fd",
          2511 => x"ff",
          2512 => x"c4",
          2513 => x"54",
          2514 => x"54",
          2515 => x"fc",
          2516 => x"3f",
          2517 => x"70",
          2518 => x"51",
          2519 => x"74",
          2520 => x"82",
          2521 => x"ff",
          2522 => x"29",
          2523 => x"82",
          2524 => x"75",
          2525 => x"52",
          2526 => x"f7",
          2527 => x"2c",
          2528 => x"57",
          2529 => x"fb",
          2530 => x"ce",
          2531 => x"80",
          2532 => x"d8",
          2533 => x"de",
          2534 => x"33",
          2535 => x"fb",
          2536 => x"9e",
          2537 => x"f6",
          2538 => x"ff",
          2539 => x"d8",
          2540 => x"81",
          2541 => x"3f",
          2542 => x"82",
          2543 => x"d8",
          2544 => x"3d",
          2545 => x"73",
          2546 => x"fc",
          2547 => x"3f",
          2548 => x"73",
          2549 => x"06",
          2550 => x"82",
          2551 => x"2e",
          2552 => x"82",
          2553 => x"98",
          2554 => x"55",
          2555 => x"54",
          2556 => x"fc",
          2557 => x"f6",
          2558 => x"80",
          2559 => x"d8",
          2560 => x"d5",
          2561 => x"51",
          2562 => x"33",
          2563 => x"f7",
          2564 => x"74",
          2565 => x"08",
          2566 => x"74",
          2567 => x"05",
          2568 => x"58",
          2569 => x"f7",
          2570 => x"81",
          2571 => x"56",
          2572 => x"82",
          2573 => x"73",
          2574 => x"33",
          2575 => x"f7",
          2576 => x"f7",
          2577 => x"26",
          2578 => x"dc",
          2579 => x"ee",
          2580 => x"34",
          2581 => x"9c",
          2582 => x"08",
          2583 => x"51",
          2584 => x"08",
          2585 => x"08",
          2586 => x"52",
          2587 => x"5b",
          2588 => x"df",
          2589 => x"74",
          2590 => x"9a",
          2591 => x"f7",
          2592 => x"ff",
          2593 => x"51",
          2594 => x"80",
          2595 => x"2e",
          2596 => x"91",
          2597 => x"81",
          2598 => x"55",
          2599 => x"ff",
          2600 => x"82",
          2601 => x"81",
          2602 => x"79",
          2603 => x"39",
          2604 => x"70",
          2605 => x"38",
          2606 => x"e0",
          2607 => x"e0",
          2608 => x"53",
          2609 => x"3f",
          2610 => x"5b",
          2611 => x"74",
          2612 => x"f7",
          2613 => x"3f",
          2614 => x"70",
          2615 => x"59",
          2616 => x"38",
          2617 => x"54",
          2618 => x"70",
          2619 => x"f4",
          2620 => x"73",
          2621 => x"fc",
          2622 => x"3f",
          2623 => x"73",
          2624 => x"f9",
          2625 => x"e0",
          2626 => x"84",
          2627 => x"84",
          2628 => x"82",
          2629 => x"74",
          2630 => x"82",
          2631 => x"34",
          2632 => x"08",
          2633 => x"15",
          2634 => x"84",
          2635 => x"70",
          2636 => x"58",
          2637 => x"73",
          2638 => x"70",
          2639 => x"f8",
          2640 => x"34",
          2641 => x"04",
          2642 => x"84",
          2643 => x"2a",
          2644 => x"51",
          2645 => x"83",
          2646 => x"a6",
          2647 => x"22",
          2648 => x"83",
          2649 => x"11",
          2650 => x"2b",
          2651 => x"71",
          2652 => x"2a",
          2653 => x"57",
          2654 => x"81",
          2655 => x"75",
          2656 => x"34",
          2657 => x"08",
          2658 => x"71",
          2659 => x"ff",
          2660 => x"05",
          2661 => x"2a",
          2662 => x"72",
          2663 => x"34",
          2664 => x"76",
          2665 => x"0d",
          2666 => x"08",
          2667 => x"83",
          2668 => x"12",
          2669 => x"07",
          2670 => x"05",
          2671 => x"88",
          2672 => x"56",
          2673 => x"13",
          2674 => x"84",
          2675 => x"2b",
          2676 => x"52",
          2677 => x"33",
          2678 => x"54",
          2679 => x"73",
          2680 => x"13",
          2681 => x"2b",
          2682 => x"88",
          2683 => x"73",
          2684 => x"0d",
          2685 => x"22",
          2686 => x"71",
          2687 => x"88",
          2688 => x"33",
          2689 => x"90",
          2690 => x"5a",
          2691 => x"80",
          2692 => x"82",
          2693 => x"81",
          2694 => x"2b",
          2695 => x"33",
          2696 => x"8f",
          2697 => x"53",
          2698 => x"2a",
          2699 => x"83",
          2700 => x"16",
          2701 => x"2b",
          2702 => x"55",
          2703 => x"71",
          2704 => x"06",
          2705 => x"52",
          2706 => x"88",
          2707 => x"e0",
          2708 => x"22",
          2709 => x"33",
          2710 => x"83",
          2711 => x"52",
          2712 => x"71",
          2713 => x"05",
          2714 => x"51",
          2715 => x"81",
          2716 => x"15",
          2717 => x"2b",
          2718 => x"52",
          2719 => x"33",
          2720 => x"54",
          2721 => x"72",
          2722 => x"14",
          2723 => x"88",
          2724 => x"54",
          2725 => x"7b",
          2726 => x"70",
          2727 => x"53",
          2728 => x"76",
          2729 => x"83",
          2730 => x"2b",
          2731 => x"33",
          2732 => x"53",
          2733 => x"59",
          2734 => x"80",
          2735 => x"81",
          2736 => x"33",
          2737 => x"76",
          2738 => x"58",
          2739 => x"ff",
          2740 => x"e0",
          2741 => x"85",
          2742 => x"88",
          2743 => x"84",
          2744 => x"e0",
          2745 => x"14",
          2746 => x"e0",
          2747 => x"75",
          2748 => x"18",
          2749 => x"2b",
          2750 => x"88",
          2751 => x"74",
          2752 => x"0d",
          2753 => x"e0",
          2754 => x"71",
          2755 => x"8c",
          2756 => x"0d",
          2757 => x"82",
          2758 => x"82",
          2759 => x"12",
          2760 => x"59",
          2761 => x"75",
          2762 => x"29",
          2763 => x"88",
          2764 => x"79",
          2765 => x"7f",
          2766 => x"77",
          2767 => x"85",
          2768 => x"33",
          2769 => x"57",
          2770 => x"ff",
          2771 => x"80",
          2772 => x"11",
          2773 => x"2b",
          2774 => x"52",
          2775 => x"83",
          2776 => x"26",
          2777 => x"2e",
          2778 => x"81",
          2779 => x"3f",
          2780 => x"79",
          2781 => x"e0",
          2782 => x"87",
          2783 => x"2b",
          2784 => x"7a",
          2785 => x"88",
          2786 => x"15",
          2787 => x"85",
          2788 => x"83",
          2789 => x"33",
          2790 => x"70",
          2791 => x"56",
          2792 => x"19",
          2793 => x"84",
          2794 => x"2b",
          2795 => x"55",
          2796 => x"76",
          2797 => x"70",
          2798 => x"12",
          2799 => x"2a",
          2800 => x"84",
          2801 => x"e0",
          2802 => x"82",
          2803 => x"fe",
          2804 => x"08",
          2805 => x"71",
          2806 => x"ed",
          2807 => x"82",
          2808 => x"ee",
          2809 => x"70",
          2810 => x"2e",
          2811 => x"3f",
          2812 => x"3f",
          2813 => x"39",
          2814 => x"3f",
          2815 => x"f5",
          2816 => x"ff",
          2817 => x"71",
          2818 => x"06",
          2819 => x"81",
          2820 => x"75",
          2821 => x"88",
          2822 => x"70",
          2823 => x"07",
          2824 => x"48",
          2825 => x"56",
          2826 => x"76",
          2827 => x"83",
          2828 => x"33",
          2829 => x"70",
          2830 => x"33",
          2831 => x"53",
          2832 => x"25",
          2833 => x"ff",
          2834 => x"81",
          2835 => x"2e",
          2836 => x"f6",
          2837 => x"58",
          2838 => x"74",
          2839 => x"3f",
          2840 => x"75",
          2841 => x"11",
          2842 => x"07",
          2843 => x"52",
          2844 => x"98",
          2845 => x"7c",
          2846 => x"08",
          2847 => x"87",
          2848 => x"84",
          2849 => x"5c",
          2850 => x"74",
          2851 => x"c9",
          2852 => x"11",
          2853 => x"07",
          2854 => x"52",
          2855 => x"98",
          2856 => x"7c",
          2857 => x"08",
          2858 => x"86",
          2859 => x"84",
          2860 => x"73",
          2861 => x"7b",
          2862 => x"e0",
          2863 => x"80",
          2864 => x"82",
          2865 => x"3f",
          2866 => x"7a",
          2867 => x"52",
          2868 => x"83",
          2869 => x"05",
          2870 => x"82",
          2871 => x"fc",
          2872 => x"54",
          2873 => x"55",
          2874 => x"38",
          2875 => x"08",
          2876 => x"e0",
          2877 => x"3d",
          2878 => x"52",
          2879 => x"94",
          2880 => x"0c",
          2881 => x"02",
          2882 => x"05",
          2883 => x"26",
          2884 => x"c0",
          2885 => x"74",
          2886 => x"73",
          2887 => x"51",
          2888 => x"98",
          2889 => x"82",
          2890 => x"38",
          2891 => x"ec",
          2892 => x"52",
          2893 => x"08",
          2894 => x"82",
          2895 => x"13",
          2896 => x"86",
          2897 => x"62",
          2898 => x"57",
          2899 => x"fe",
          2900 => x"06",
          2901 => x"71",
          2902 => x"80",
          2903 => x"c0",
          2904 => x"5a",
          2905 => x"0c",
          2906 => x"08",
          2907 => x"53",
          2908 => x"08",
          2909 => x"34",
          2910 => x"53",
          2911 => x"53",
          2912 => x"80",
          2913 => x"08",
          2914 => x"8c",
          2915 => x"78",
          2916 => x"0c",
          2917 => x"08",
          2918 => x"38",
          2919 => x"17",
          2920 => x"53",
          2921 => x"fc",
          2922 => x"7d",
          2923 => x"80",
          2924 => x"38",
          2925 => x"98",
          2926 => x"0d",
          2927 => x"05",
          2928 => x"80",
          2929 => x"e0",
          2930 => x"71",
          2931 => x"38",
          2932 => x"80",
          2933 => x"c0",
          2934 => x"5a",
          2935 => x"76",
          2936 => x"75",
          2937 => x"51",
          2938 => x"7a",
          2939 => x"81",
          2940 => x"06",
          2941 => x"87",
          2942 => x"38",
          2943 => x"80",
          2944 => x"99",
          2945 => x"8c",
          2946 => x"51",
          2947 => x"8d",
          2948 => x"84",
          2949 => x"2e",
          2950 => x"52",
          2951 => x"f8",
          2952 => x"71",
          2953 => x"53",
          2954 => x"0d",
          2955 => x"05",
          2956 => x"05",
          2957 => x"fe",
          2958 => x"53",
          2959 => x"0b",
          2960 => x"71",
          2961 => x"24",
          2962 => x"92",
          2963 => x"8d",
          2964 => x"80",
          2965 => x"70",
          2966 => x"52",
          2967 => x"98",
          2968 => x"c0",
          2969 => x"81",
          2970 => x"53",
          2971 => x"71",
          2972 => x"39",
          2973 => x"81",
          2974 => x"84",
          2975 => x"0c",
          2976 => x"74",
          2977 => x"2b",
          2978 => x"84",
          2979 => x"83",
          2980 => x"2b",
          2981 => x"70",
          2982 => x"07",
          2983 => x"56",
          2984 => x"3d",
          2985 => x"22",
          2986 => x"54",
          2987 => x"34",
          2988 => x"73",
          2989 => x"05",
          2990 => x"72",
          2991 => x"2a",
          2992 => x"34",
          2993 => x"83",
          2994 => x"75",
          2995 => x"92",
          2996 => x"73",
          2997 => x"51",
          2998 => x"3d",
          2999 => x"72",
          3000 => x"11",
          3001 => x"04",
          3002 => x"56",
          3003 => x"74",
          3004 => x"31",
          3005 => x"80",
          3006 => x"38",
          3007 => x"0d",
          3008 => x"51",
          3009 => x"81",
          3010 => x"38",
          3011 => x"3d",
          3012 => x"0c",
          3013 => x"70",
          3014 => x"55",
          3015 => x"e0",
          3016 => x"98",
          3017 => x"f9",
          3018 => x"ff",
          3019 => x"38",
          3020 => x"e0",
          3021 => x"3d",
          3022 => x"33",
          3023 => x"38",
          3024 => x"16",
          3025 => x"f9",
          3026 => x"2e",
          3027 => x"98",
          3028 => x"70",
          3029 => x"59",
          3030 => x"82",
          3031 => x"81",
          3032 => x"53",
          3033 => x"a5",
          3034 => x"e0",
          3035 => x"3d",
          3036 => x"74",
          3037 => x"51",
          3038 => x"57",
          3039 => x"54",
          3040 => x"33",
          3041 => x"08",
          3042 => x"57",
          3043 => x"98",
          3044 => x"0d",
          3045 => x"82",
          3046 => x"08",
          3047 => x"83",
          3048 => x"84",
          3049 => x"81",
          3050 => x"82",
          3051 => x"52",
          3052 => x"52",
          3053 => x"84",
          3054 => x"fb",
          3055 => x"52",
          3056 => x"94",
          3057 => x"fb",
          3058 => x"a4",
          3059 => x"08",
          3060 => x"55",
          3061 => x"f7",
          3062 => x"53",
          3063 => x"99",
          3064 => x"83",
          3065 => x"0c",
          3066 => x"77",
          3067 => x"55",
          3068 => x"8d",
          3069 => x"b0",
          3070 => x"e0",
          3071 => x"3d",
          3072 => x"57",
          3073 => x"9c",
          3074 => x"74",
          3075 => x"f5",
          3076 => x"81",
          3077 => x"83",
          3078 => x"76",
          3079 => x"16",
          3080 => x"96",
          3081 => x"38",
          3082 => x"33",
          3083 => x"08",
          3084 => x"fc",
          3085 => x"fe",
          3086 => x"11",
          3087 => x"81",
          3088 => x"51",
          3089 => x"ff",
          3090 => x"2a",
          3091 => x"fc",
          3092 => x"c6",
          3093 => x"05",
          3094 => x"e0",
          3095 => x"ae",
          3096 => x"05",
          3097 => x"e0",
          3098 => x"83",
          3099 => x"f8",
          3100 => x"0a",
          3101 => x"82",
          3102 => x"f8",
          3103 => x"56",
          3104 => x"38",
          3105 => x"38",
          3106 => x"9d",
          3107 => x"81",
          3108 => x"83",
          3109 => x"76",
          3110 => x"18",
          3111 => x"9e",
          3112 => x"e0",
          3113 => x"ff",
          3114 => x"81",
          3115 => x"80",
          3116 => x"f0",
          3117 => x"51",
          3118 => x"17",
          3119 => x"05",
          3120 => x"e0",
          3121 => x"81",
          3122 => x"b8",
          3123 => x"8f",
          3124 => x"f0",
          3125 => x"72",
          3126 => x"2a",
          3127 => x"fa",
          3128 => x"82",
          3129 => x"83",
          3130 => x"fe",
          3131 => x"e6",
          3132 => x"17",
          3133 => x"3f",
          3134 => x"98",
          3135 => x"77",
          3136 => x"b8",
          3137 => x"8b",
          3138 => x"06",
          3139 => x"3f",
          3140 => x"e0",
          3141 => x"3d",
          3142 => x"56",
          3143 => x"74",
          3144 => x"80",
          3145 => x"75",
          3146 => x"08",
          3147 => x"38",
          3148 => x"81",
          3149 => x"08",
          3150 => x"51",
          3151 => x"58",
          3152 => x"c7",
          3153 => x"d2",
          3154 => x"cf",
          3155 => x"fc",
          3156 => x"38",
          3157 => x"08",
          3158 => x"38",
          3159 => x"33",
          3160 => x"77",
          3161 => x"80",
          3162 => x"3d",
          3163 => x"71",
          3164 => x"90",
          3165 => x"38",
          3166 => x"81",
          3167 => x"f9",
          3168 => x"98",
          3169 => x"98",
          3170 => x"2e",
          3171 => x"e0",
          3172 => x"58",
          3173 => x"80",
          3174 => x"09",
          3175 => x"56",
          3176 => x"82",
          3177 => x"3f",
          3178 => x"2e",
          3179 => x"98",
          3180 => x"70",
          3181 => x"7c",
          3182 => x"51",
          3183 => x"e0",
          3184 => x"17",
          3185 => x"73",
          3186 => x"58",
          3187 => x"56",
          3188 => x"26",
          3189 => x"81",
          3190 => x"c6",
          3191 => x"b8",
          3192 => x"81",
          3193 => x"e0",
          3194 => x"09",
          3195 => x"70",
          3196 => x"80",
          3197 => x"06",
          3198 => x"39",
          3199 => x"f7",
          3200 => x"98",
          3201 => x"07",
          3202 => x"2e",
          3203 => x"75",
          3204 => x"3f",
          3205 => x"38",
          3206 => x"fe",
          3207 => x"74",
          3208 => x"0c",
          3209 => x"84",
          3210 => x"81",
          3211 => x"8c",
          3212 => x"39",
          3213 => x"98",
          3214 => x"0d",
          3215 => x"82",
          3216 => x"e0",
          3217 => x"74",
          3218 => x"08",
          3219 => x"59",
          3220 => x"70",
          3221 => x"84",
          3222 => x"58",
          3223 => x"75",
          3224 => x"51",
          3225 => x"80",
          3226 => x"32",
          3227 => x"2a",
          3228 => x"98",
          3229 => x"0d",
          3230 => x"74",
          3231 => x"74",
          3232 => x"74",
          3233 => x"73",
          3234 => x"27",
          3235 => x"9b",
          3236 => x"88",
          3237 => x"80",
          3238 => x"0c",
          3239 => x"89",
          3240 => x"38",
          3241 => x"82",
          3242 => x"08",
          3243 => x"e0",
          3244 => x"08",
          3245 => x"82",
          3246 => x"cb",
          3247 => x"3f",
          3248 => x"73",
          3249 => x"82",
          3250 => x"39",
          3251 => x"13",
          3252 => x"16",
          3253 => x"77",
          3254 => x"04",
          3255 => x"12",
          3256 => x"80",
          3257 => x"98",
          3258 => x"55",
          3259 => x"83",
          3260 => x"81",
          3261 => x"55",
          3262 => x"17",
          3263 => x"9b",
          3264 => x"ff",
          3265 => x"81",
          3266 => x"e6",
          3267 => x"55",
          3268 => x"80",
          3269 => x"08",
          3270 => x"08",
          3271 => x"38",
          3272 => x"84",
          3273 => x"52",
          3274 => x"98",
          3275 => x"08",
          3276 => x"82",
          3277 => x"81",
          3278 => x"b0",
          3279 => x"51",
          3280 => x"a0",
          3281 => x"75",
          3282 => x"08",
          3283 => x"77",
          3284 => x"55",
          3285 => x"0d",
          3286 => x"08",
          3287 => x"fc",
          3288 => x"82",
          3289 => x"e0",
          3290 => x"78",
          3291 => x"08",
          3292 => x"38",
          3293 => x"70",
          3294 => x"2e",
          3295 => x"82",
          3296 => x"81",
          3297 => x"2e",
          3298 => x"2e",
          3299 => x"82",
          3300 => x"51",
          3301 => x"54",
          3302 => x"9b",
          3303 => x"83",
          3304 => x"0c",
          3305 => x"76",
          3306 => x"82",
          3307 => x"76",
          3308 => x"2e",
          3309 => x"51",
          3310 => x"90",
          3311 => x"98",
          3312 => x"0d",
          3313 => x"54",
          3314 => x"3f",
          3315 => x"2e",
          3316 => x"2a",
          3317 => x"86",
          3318 => x"54",
          3319 => x"71",
          3320 => x"05",
          3321 => x"06",
          3322 => x"e4",
          3323 => x"3d",
          3324 => x"40",
          3325 => x"ff",
          3326 => x"2e",
          3327 => x"7d",
          3328 => x"08",
          3329 => x"38",
          3330 => x"73",
          3331 => x"8b",
          3332 => x"06",
          3333 => x"e0",
          3334 => x"09",
          3335 => x"e0",
          3336 => x"81",
          3337 => x"07",
          3338 => x"08",
          3339 => x"2e",
          3340 => x"75",
          3341 => x"81",
          3342 => x"06",
          3343 => x"81",
          3344 => x"38",
          3345 => x"70",
          3346 => x"5d",
          3347 => x"81",
          3348 => x"73",
          3349 => x"8c",
          3350 => x"cc",
          3351 => x"ff",
          3352 => x"33",
          3353 => x"05",
          3354 => x"d2",
          3355 => x"a4",
          3356 => x"ff",
          3357 => x"73",
          3358 => x"10",
          3359 => x"81",
          3360 => x"ff",
          3361 => x"17",
          3362 => x"33",
          3363 => x"54",
          3364 => x"81",
          3365 => x"53",
          3366 => x"ff",
          3367 => x"53",
          3368 => x"74",
          3369 => x"08",
          3370 => x"a7",
          3371 => x"39",
          3372 => x"82",
          3373 => x"08",
          3374 => x"38",
          3375 => x"7a",
          3376 => x"04",
          3377 => x"59",
          3378 => x"82",
          3379 => x"08",
          3380 => x"5c",
          3381 => x"08",
          3382 => x"e0",
          3383 => x"83",
          3384 => x"57",
          3385 => x"f6",
          3386 => x"81",
          3387 => x"34",
          3388 => x"74",
          3389 => x"74",
          3390 => x"38",
          3391 => x"f7",
          3392 => x"70",
          3393 => x"a1",
          3394 => x"51",
          3395 => x"17",
          3396 => x"1c",
          3397 => x"75",
          3398 => x"38",
          3399 => x"09",
          3400 => x"08",
          3401 => x"82",
          3402 => x"55",
          3403 => x"bf",
          3404 => x"81",
          3405 => x"33",
          3406 => x"e0",
          3407 => x"79",
          3408 => x"26",
          3409 => x"a0",
          3410 => x"1e",
          3411 => x"55",
          3412 => x"98",
          3413 => x"38",
          3414 => x"ff",
          3415 => x"1b",
          3416 => x"76",
          3417 => x"51",
          3418 => x"73",
          3419 => x"70",
          3420 => x"1c",
          3421 => x"39",
          3422 => x"7b",
          3423 => x"82",
          3424 => x"73",
          3425 => x"81",
          3426 => x"a0",
          3427 => x"b0",
          3428 => x"9e",
          3429 => x"1a",
          3430 => x"3f",
          3431 => x"98",
          3432 => x"82",
          3433 => x"ee",
          3434 => x"33",
          3435 => x"55",
          3436 => x"08",
          3437 => x"2e",
          3438 => x"70",
          3439 => x"53",
          3440 => x"53",
          3441 => x"cb",
          3442 => x"2e",
          3443 => x"1b",
          3444 => x"56",
          3445 => x"e3",
          3446 => x"38",
          3447 => x"ff",
          3448 => x"38",
          3449 => x"59",
          3450 => x"10",
          3451 => x"70",
          3452 => x"80",
          3453 => x"32",
          3454 => x"db",
          3455 => x"84",
          3456 => x"07",
          3457 => x"38",
          3458 => x"16",
          3459 => x"56",
          3460 => x"17",
          3461 => x"27",
          3462 => x"2e",
          3463 => x"54",
          3464 => x"80",
          3465 => x"74",
          3466 => x"15",
          3467 => x"19",
          3468 => x"3d",
          3469 => x"81",
          3470 => x"26",
          3471 => x"33",
          3472 => x"75",
          3473 => x"3f",
          3474 => x"1b",
          3475 => x"38",
          3476 => x"f0",
          3477 => x"e0",
          3478 => x"82",
          3479 => x"ab",
          3480 => x"70",
          3481 => x"5e",
          3482 => x"8d",
          3483 => x"3f",
          3484 => x"52",
          3485 => x"98",
          3486 => x"9e",
          3487 => x"81",
          3488 => x"08",
          3489 => x"dd",
          3490 => x"e0",
          3491 => x"51",
          3492 => x"81",
          3493 => x"7b",
          3494 => x"08",
          3495 => x"38",
          3496 => x"81",
          3497 => x"17",
          3498 => x"e0",
          3499 => x"98",
          3500 => x"3f",
          3501 => x"55",
          3502 => x"74",
          3503 => x"51",
          3504 => x"33",
          3505 => x"85",
          3506 => x"57",
          3507 => x"ff",
          3508 => x"70",
          3509 => x"80",
          3510 => x"0b",
          3511 => x"ef",
          3512 => x"82",
          3513 => x"19",
          3514 => x"08",
          3515 => x"e0",
          3516 => x"ae",
          3517 => x"52",
          3518 => x"8b",
          3519 => x"51",
          3520 => x"1b",
          3521 => x"16",
          3522 => x"55",
          3523 => x"0d",
          3524 => x"90",
          3525 => x"57",
          3526 => x"52",
          3527 => x"98",
          3528 => x"c9",
          3529 => x"e1",
          3530 => x"82",
          3531 => x"08",
          3532 => x"17",
          3533 => x"38",
          3534 => x"ee",
          3535 => x"82",
          3536 => x"73",
          3537 => x"82",
          3538 => x"3d",
          3539 => x"71",
          3540 => x"19",
          3541 => x"e2",
          3542 => x"bb",
          3543 => x"08",
          3544 => x"72",
          3545 => x"14",
          3546 => x"7a",
          3547 => x"83",
          3548 => x"ff",
          3549 => x"39",
          3550 => x"31",
          3551 => x"90",
          3552 => x"3f",
          3553 => x"06",
          3554 => x"81",
          3555 => x"53",
          3556 => x"82",
          3557 => x"70",
          3558 => x"07",
          3559 => x"38",
          3560 => x"81",
          3561 => x"1d",
          3562 => x"54",
          3563 => x"70",
          3564 => x"51",
          3565 => x"0b",
          3566 => x"58",
          3567 => x"33",
          3568 => x"2e",
          3569 => x"06",
          3570 => x"32",
          3571 => x"51",
          3572 => x"72",
          3573 => x"81",
          3574 => x"76",
          3575 => x"57",
          3576 => x"17",
          3577 => x"34",
          3578 => x"38",
          3579 => x"34",
          3580 => x"89",
          3581 => x"2e",
          3582 => x"55",
          3583 => x"55",
          3584 => x"08",
          3585 => x"27",
          3586 => x"39",
          3587 => x"53",
          3588 => x"70",
          3589 => x"76",
          3590 => x"81",
          3591 => x"55",
          3592 => x"94",
          3593 => x"9c",
          3594 => x"72",
          3595 => x"1c",
          3596 => x"34",
          3597 => x"d9",
          3598 => x"0c",
          3599 => x"e0",
          3600 => x"51",
          3601 => x"84",
          3602 => x"3d",
          3603 => x"64",
          3604 => x"2e",
          3605 => x"2e",
          3606 => x"7f",
          3607 => x"39",
          3608 => x"56",
          3609 => x"06",
          3610 => x"32",
          3611 => x"51",
          3612 => x"1f",
          3613 => x"9f",
          3614 => x"1f",
          3615 => x"3f",
          3616 => x"39",
          3617 => x"5b",
          3618 => x"51",
          3619 => x"ff",
          3620 => x"0b",
          3621 => x"78",
          3622 => x"2a",
          3623 => x"59",
          3624 => x"06",
          3625 => x"27",
          3626 => x"56",
          3627 => x"ae",
          3628 => x"75",
          3629 => x"3f",
          3630 => x"78",
          3631 => x"10",
          3632 => x"59",
          3633 => x"61",
          3634 => x"2e",
          3635 => x"73",
          3636 => x"25",
          3637 => x"38",
          3638 => x"57",
          3639 => x"38",
          3640 => x"38",
          3641 => x"81",
          3642 => x"54",
          3643 => x"c1",
          3644 => x"09",
          3645 => x"54",
          3646 => x"56",
          3647 => x"38",
          3648 => x"57",
          3649 => x"e9",
          3650 => x"1f",
          3651 => x"a8",
          3652 => x"74",
          3653 => x"70",
          3654 => x"58",
          3655 => x"73",
          3656 => x"38",
          3657 => x"74",
          3658 => x"90",
          3659 => x"39",
          3660 => x"06",
          3661 => x"81",
          3662 => x"1b",
          3663 => x"2e",
          3664 => x"ff",
          3665 => x"81",
          3666 => x"78",
          3667 => x"05",
          3668 => x"9d",
          3669 => x"ff",
          3670 => x"fe",
          3671 => x"2e",
          3672 => x"a0",
          3673 => x"80",
          3674 => x"1a",
          3675 => x"75",
          3676 => x"2e",
          3677 => x"70",
          3678 => x"2e",
          3679 => x"76",
          3680 => x"73",
          3681 => x"5b",
          3682 => x"07",
          3683 => x"55",
          3684 => x"8b",
          3685 => x"8b",
          3686 => x"26",
          3687 => x"8b",
          3688 => x"5f",
          3689 => x"af",
          3690 => x"52",
          3691 => x"e0",
          3692 => x"87",
          3693 => x"73",
          3694 => x"06",
          3695 => x"81",
          3696 => x"54",
          3697 => x"07",
          3698 => x"18",
          3699 => x"73",
          3700 => x"39",
          3701 => x"82",
          3702 => x"e0",
          3703 => x"df",
          3704 => x"ff",
          3705 => x"38",
          3706 => x"54",
          3707 => x"07",
          3708 => x"58",
          3709 => x"75",
          3710 => x"39",
          3711 => x"2e",
          3712 => x"a0",
          3713 => x"06",
          3714 => x"06",
          3715 => x"2e",
          3716 => x"83",
          3717 => x"82",
          3718 => x"06",
          3719 => x"06",
          3720 => x"90",
          3721 => x"06",
          3722 => x"76",
          3723 => x"7d",
          3724 => x"08",
          3725 => x"98",
          3726 => x"98",
          3727 => x"e8",
          3728 => x"76",
          3729 => x"2e",
          3730 => x"80",
          3731 => x"ab",
          3732 => x"74",
          3733 => x"56",
          3734 => x"06",
          3735 => x"33",
          3736 => x"55",
          3737 => x"1e",
          3738 => x"05",
          3739 => x"e0",
          3740 => x"39",
          3741 => x"0d",
          3742 => x"7b",
          3743 => x"55",
          3744 => x"75",
          3745 => x"26",
          3746 => x"70",
          3747 => x"06",
          3748 => x"70",
          3749 => x"89",
          3750 => x"ff",
          3751 => x"2e",
          3752 => x"98",
          3753 => x"76",
          3754 => x"81",
          3755 => x"53",
          3756 => x"13",
          3757 => x"9f",
          3758 => x"e0",
          3759 => x"72",
          3760 => x"72",
          3761 => x"ff",
          3762 => x"70",
          3763 => x"9f",
          3764 => x"80",
          3765 => x"59",
          3766 => x"8b",
          3767 => x"76",
          3768 => x"82",
          3769 => x"98",
          3770 => x"0d",
          3771 => x"ff",
          3772 => x"51",
          3773 => x"98",
          3774 => x"51",
          3775 => x"83",
          3776 => x"82",
          3777 => x"e3",
          3778 => x"57",
          3779 => x"83",
          3780 => x"70",
          3781 => x"51",
          3782 => x"2e",
          3783 => x"82",
          3784 => x"cf",
          3785 => x"82",
          3786 => x"85",
          3787 => x"16",
          3788 => x"08",
          3789 => x"83",
          3790 => x"0c",
          3791 => x"61",
          3792 => x"58",
          3793 => x"e1",
          3794 => x"56",
          3795 => x"87",
          3796 => x"29",
          3797 => x"53",
          3798 => x"38",
          3799 => x"74",
          3800 => x"38",
          3801 => x"82",
          3802 => x"81",
          3803 => x"80",
          3804 => x"70",
          3805 => x"86",
          3806 => x"34",
          3807 => x"33",
          3808 => x"33",
          3809 => x"08",
          3810 => x"55",
          3811 => x"80",
          3812 => x"81",
          3813 => x"b8",
          3814 => x"fd",
          3815 => x"ff",
          3816 => x"76",
          3817 => x"8d",
          3818 => x"90",
          3819 => x"56",
          3820 => x"72",
          3821 => x"51",
          3822 => x"57",
          3823 => x"ff",
          3824 => x"25",
          3825 => x"11",
          3826 => x"71",
          3827 => x"f0",
          3828 => x"74",
          3829 => x"90",
          3830 => x"3f",
          3831 => x"57",
          3832 => x"54",
          3833 => x"83",
          3834 => x"38",
          3835 => x"84",
          3836 => x"38",
          3837 => x"38",
          3838 => x"38",
          3839 => x"82",
          3840 => x"53",
          3841 => x"84",
          3842 => x"ec",
          3843 => x"ff",
          3844 => x"14",
          3845 => x"08",
          3846 => x"14",
          3847 => x"33",
          3848 => x"54",
          3849 => x"98",
          3850 => x"29",
          3851 => x"72",
          3852 => x"38",
          3853 => x"2e",
          3854 => x"80",
          3855 => x"e0",
          3856 => x"88",
          3857 => x"56",
          3858 => x"51",
          3859 => x"83",
          3860 => x"80",
          3861 => x"e0",
          3862 => x"c8",
          3863 => x"ff",
          3864 => x"2e",
          3865 => x"14",
          3866 => x"75",
          3867 => x"52",
          3868 => x"3f",
          3869 => x"98",
          3870 => x"e0",
          3871 => x"26",
          3872 => x"f5",
          3873 => x"f5",
          3874 => x"8d",
          3875 => x"82",
          3876 => x"16",
          3877 => x"7a",
          3878 => x"83",
          3879 => x"e2",
          3880 => x"98",
          3881 => x"56",
          3882 => x"38",
          3883 => x"82",
          3884 => x"82",
          3885 => x"80",
          3886 => x"15",
          3887 => x"8d",
          3888 => x"76",
          3889 => x"13",
          3890 => x"15",
          3891 => x"94",
          3892 => x"ff",
          3893 => x"2e",
          3894 => x"e8",
          3895 => x"98",
          3896 => x"81",
          3897 => x"81",
          3898 => x"82",
          3899 => x"e0",
          3900 => x"14",
          3901 => x"08",
          3902 => x"d4",
          3903 => x"38",
          3904 => x"e0",
          3905 => x"2e",
          3906 => x"14",
          3907 => x"08",
          3908 => x"81",
          3909 => x"c5",
          3910 => x"15",
          3911 => x"3f",
          3912 => x"76",
          3913 => x"05",
          3914 => x"86",
          3915 => x"15",
          3916 => x"56",
          3917 => x"0d",
          3918 => x"55",
          3919 => x"53",
          3920 => x"52",
          3921 => x"22",
          3922 => x"2e",
          3923 => x"33",
          3924 => x"98",
          3925 => x"71",
          3926 => x"53",
          3927 => x"e0",
          3928 => x"3d",
          3929 => x"89",
          3930 => x"3f",
          3931 => x"08",
          3932 => x"84",
          3933 => x"55",
          3934 => x"74",
          3935 => x"38",
          3936 => x"54",
          3937 => x"89",
          3938 => x"e4",
          3939 => x"82",
          3940 => x"ea",
          3941 => x"eb",
          3942 => x"80",
          3943 => x"70",
          3944 => x"3d",
          3945 => x"82",
          3946 => x"08",
          3947 => x"8c",
          3948 => x"82",
          3949 => x"08",
          3950 => x"70",
          3951 => x"83",
          3952 => x"73",
          3953 => x"2e",
          3954 => x"06",
          3955 => x"82",
          3956 => x"b2",
          3957 => x"b8",
          3958 => x"51",
          3959 => x"55",
          3960 => x"74",
          3961 => x"81",
          3962 => x"af",
          3963 => x"3f",
          3964 => x"b2",
          3965 => x"f4",
          3966 => x"34",
          3967 => x"85",
          3968 => x"c2",
          3969 => x"15",
          3970 => x"7a",
          3971 => x"75",
          3972 => x"86",
          3973 => x"e0",
          3974 => x"74",
          3975 => x"70",
          3976 => x"56",
          3977 => x"82",
          3978 => x"06",
          3979 => x"75",
          3980 => x"38",
          3981 => x"7a",
          3982 => x"08",
          3983 => x"55",
          3984 => x"77",
          3985 => x"73",
          3986 => x"07",
          3987 => x"0c",
          3988 => x"52",
          3989 => x"08",
          3990 => x"63",
          3991 => x"82",
          3992 => x"8c",
          3993 => x"17",
          3994 => x"34",
          3995 => x"9c",
          3996 => x"77",
          3997 => x"73",
          3998 => x"98",
          3999 => x"e0",
          4000 => x"22",
          4001 => x"a8",
          4002 => x"3f",
          4003 => x"98",
          4004 => x"82",
          4005 => x"06",
          4006 => x"56",
          4007 => x"51",
          4008 => x"70",
          4009 => x"76",
          4010 => x"83",
          4011 => x"38",
          4012 => x"82",
          4013 => x"8e",
          4014 => x"08",
          4015 => x"79",
          4016 => x"0c",
          4017 => x"60",
          4018 => x"80",
          4019 => x"78",
          4020 => x"08",
          4021 => x"91",
          4022 => x"38",
          4023 => x"33",
          4024 => x"2e",
          4025 => x"91",
          4026 => x"81",
          4027 => x"a3",
          4028 => x"31",
          4029 => x"5c",
          4030 => x"19",
          4031 => x"74",
          4032 => x"ff",
          4033 => x"79",
          4034 => x"08",
          4035 => x"78",
          4036 => x"08",
          4037 => x"74",
          4038 => x"1a",
          4039 => x"c3",
          4040 => x"2e",
          4041 => x"1a",
          4042 => x"2e",
          4043 => x"11",
          4044 => x"85",
          4045 => x"76",
          4046 => x"ff",
          4047 => x"fe",
          4048 => x"56",
          4049 => x"08",
          4050 => x"38",
          4051 => x"16",
          4052 => x"51",
          4053 => x"56",
          4054 => x"19",
          4055 => x"31",
          4056 => x"7b",
          4057 => x"c0",
          4058 => x"ff",
          4059 => x"ff",
          4060 => x"ff",
          4061 => x"08",
          4062 => x"08",
          4063 => x"f0",
          4064 => x"0c",
          4065 => x"60",
          4066 => x"80",
          4067 => x"77",
          4068 => x"08",
          4069 => x"91",
          4070 => x"38",
          4071 => x"33",
          4072 => x"56",
          4073 => x"ab",
          4074 => x"34",
          4075 => x"91",
          4076 => x"94",
          4077 => x"76",
          4078 => x"80",
          4079 => x"70",
          4080 => x"82",
          4081 => x"77",
          4082 => x"38",
          4083 => x"74",
          4084 => x"18",
          4085 => x"82",
          4086 => x"08",
          4087 => x"2e",
          4088 => x"95",
          4089 => x"08",
          4090 => x"55",
          4091 => x"09",
          4092 => x"bd",
          4093 => x"ed",
          4094 => x"ff",
          4095 => x"80",
          4096 => x"08",
          4097 => x"80",
          4098 => x"8a",
          4099 => x"27",
          4100 => x"54",
          4101 => x"51",
          4102 => x"08",
          4103 => x"78",
          4104 => x"38",
          4105 => x"31",
          4106 => x"51",
          4107 => x"0b",
          4108 => x"80",
          4109 => x"08",
          4110 => x"f6",
          4111 => x"38",
          4112 => x"9c",
          4113 => x"06",
          4114 => x"76",
          4115 => x"08",
          4116 => x"82",
          4117 => x"53",
          4118 => x"06",
          4119 => x"3f",
          4120 => x"7b",
          4121 => x"76",
          4122 => x"1c",
          4123 => x"5c",
          4124 => x"74",
          4125 => x"18",
          4126 => x"19",
          4127 => x"0c",
          4128 => x"7a",
          4129 => x"56",
          4130 => x"57",
          4131 => x"90",
          4132 => x"06",
          4133 => x"ee",
          4134 => x"ff",
          4135 => x"57",
          4136 => x"a4",
          4137 => x"55",
          4138 => x"08",
          4139 => x"a5",
          4140 => x"51",
          4141 => x"0a",
          4142 => x"3f",
          4143 => x"c6",
          4144 => x"34",
          4145 => x"e0",
          4146 => x"06",
          4147 => x"82",
          4148 => x"fc",
          4149 => x"d4",
          4150 => x"e0",
          4151 => x"05",
          4152 => x"e0",
          4153 => x"87",
          4154 => x"72",
          4155 => x"04",
          4156 => x"89",
          4157 => x"98",
          4158 => x"08",
          4159 => x"82",
          4160 => x"ee",
          4161 => x"05",
          4162 => x"82",
          4163 => x"08",
          4164 => x"94",
          4165 => x"82",
          4166 => x"08",
          4167 => x"70",
          4168 => x"89",
          4169 => x"b2",
          4170 => x"2a",
          4171 => x"80",
          4172 => x"52",
          4173 => x"08",
          4174 => x"98",
          4175 => x"38",
          4176 => x"94",
          4177 => x"80",
          4178 => x"5b",
          4179 => x"df",
          4180 => x"3d",
          4181 => x"08",
          4182 => x"38",
          4183 => x"98",
          4184 => x"58",
          4185 => x"2e",
          4186 => x"3d",
          4187 => x"e0",
          4188 => x"82",
          4189 => x"7b",
          4190 => x"98",
          4191 => x"d8",
          4192 => x"51",
          4193 => x"80",
          4194 => x"c3",
          4195 => x"82",
          4196 => x"52",
          4197 => x"98",
          4198 => x"38",
          4199 => x"c8",
          4200 => x"2e",
          4201 => x"e8",
          4202 => x"e0",
          4203 => x"84",
          4204 => x"57",
          4205 => x"80",
          4206 => x"51",
          4207 => x"11",
          4208 => x"73",
          4209 => x"05",
          4210 => x"56",
          4211 => x"54",
          4212 => x"80",
          4213 => x"55",
          4214 => x"ff",
          4215 => x"74",
          4216 => x"18",
          4217 => x"af",
          4218 => x"2e",
          4219 => x"80",
          4220 => x"74",
          4221 => x"70",
          4222 => x"08",
          4223 => x"73",
          4224 => x"1a",
          4225 => x"38",
          4226 => x"38",
          4227 => x"74",
          4228 => x"05",
          4229 => x"ba",
          4230 => x"ff",
          4231 => x"57",
          4232 => x"81",
          4233 => x"81",
          4234 => x"38",
          4235 => x"0c",
          4236 => x"0d",
          4237 => x"71",
          4238 => x"e0",
          4239 => x"82",
          4240 => x"82",
          4241 => x"76",
          4242 => x"81",
          4243 => x"72",
          4244 => x"54",
          4245 => x"78",
          4246 => x"22",
          4247 => x"78",
          4248 => x"51",
          4249 => x"08",
          4250 => x"53",
          4251 => x"08",
          4252 => x"75",
          4253 => x"31",
          4254 => x"b2",
          4255 => x"38",
          4256 => x"3f",
          4257 => x"98",
          4258 => x"e0",
          4259 => x"82",
          4260 => x"98",
          4261 => x"38",
          4262 => x"77",
          4263 => x"0c",
          4264 => x"81",
          4265 => x"2e",
          4266 => x"bb",
          4267 => x"82",
          4268 => x"98",
          4269 => x"51",
          4270 => x"08",
          4271 => x"74",
          4272 => x"14",
          4273 => x"0c",
          4274 => x"94",
          4275 => x"72",
          4276 => x"51",
          4277 => x"08",
          4278 => x"82",
          4279 => x"16",
          4280 => x"2a",
          4281 => x"15",
          4282 => x"90",
          4283 => x"33",
          4284 => x"34",
          4285 => x"2e",
          4286 => x"85",
          4287 => x"72",
          4288 => x"04",
          4289 => x"75",
          4290 => x"89",
          4291 => x"05",
          4292 => x"08",
          4293 => x"38",
          4294 => x"d4",
          4295 => x"82",
          4296 => x"16",
          4297 => x"74",
          4298 => x"84",
          4299 => x"73",
          4300 => x"52",
          4301 => x"98",
          4302 => x"14",
          4303 => x"51",
          4304 => x"08",
          4305 => x"85",
          4306 => x"2e",
          4307 => x"73",
          4308 => x"04",
          4309 => x"05",
          4310 => x"82",
          4311 => x"98",
          4312 => x"fb",
          4313 => x"05",
          4314 => x"3f",
          4315 => x"98",
          4316 => x"82",
          4317 => x"bb",
          4318 => x"80",
          4319 => x"73",
          4320 => x"08",
          4321 => x"09",
          4322 => x"39",
          4323 => x"52",
          4324 => x"73",
          4325 => x"98",
          4326 => x"07",
          4327 => x"06",
          4328 => x"98",
          4329 => x"0d",
          4330 => x"53",
          4331 => x"82",
          4332 => x"08",
          4333 => x"a6",
          4334 => x"e0",
          4335 => x"05",
          4336 => x"80",
          4337 => x"76",
          4338 => x"51",
          4339 => x"0c",
          4340 => x"63",
          4341 => x"ec",
          4342 => x"3f",
          4343 => x"98",
          4344 => x"73",
          4345 => x"13",
          4346 => x"26",
          4347 => x"39",
          4348 => x"81",
          4349 => x"33",
          4350 => x"06",
          4351 => x"76",
          4352 => x"af",
          4353 => x"2e",
          4354 => x"2e",
          4355 => x"70",
          4356 => x"7a",
          4357 => x"54",
          4358 => x"80",
          4359 => x"98",
          4360 => x"52",
          4361 => x"8e",
          4362 => x"e0",
          4363 => x"33",
          4364 => x"54",
          4365 => x"38",
          4366 => x"82",
          4367 => x"70",
          4368 => x"59",
          4369 => x"51",
          4370 => x"08",
          4371 => x"25",
          4372 => x"75",
          4373 => x"ff",
          4374 => x"94",
          4375 => x"56",
          4376 => x"e0",
          4377 => x"3d",
          4378 => x"70",
          4379 => x"98",
          4380 => x"aa",
          4381 => x"a2",
          4382 => x"70",
          4383 => x"73",
          4384 => x"08",
          4385 => x"82",
          4386 => x"08",
          4387 => x"ff",
          4388 => x"74",
          4389 => x"98",
          4390 => x"c6",
          4391 => x"09",
          4392 => x"e0",
          4393 => x"85",
          4394 => x"38",
          4395 => x"15",
          4396 => x"53",
          4397 => x"ff",
          4398 => x"56",
          4399 => x"17",
          4400 => x"18",
          4401 => x"91",
          4402 => x"98",
          4403 => x"0d",
          4404 => x"52",
          4405 => x"e0",
          4406 => x"81",
          4407 => x"52",
          4408 => x"3f",
          4409 => x"98",
          4410 => x"05",
          4411 => x"51",
          4412 => x"38",
          4413 => x"81",
          4414 => x"70",
          4415 => x"81",
          4416 => x"ba",
          4417 => x"84",
          4418 => x"73",
          4419 => x"82",
          4420 => x"81",
          4421 => x"08",
          4422 => x"54",
          4423 => x"08",
          4424 => x"38",
          4425 => x"ff",
          4426 => x"55",
          4427 => x"55",
          4428 => x"84",
          4429 => x"80",
          4430 => x"82",
          4431 => x"30",
          4432 => x"25",
          4433 => x"38",
          4434 => x"75",
          4435 => x"82",
          4436 => x"78",
          4437 => x"98",
          4438 => x"a2",
          4439 => x"53",
          4440 => x"3d",
          4441 => x"08",
          4442 => x"38",
          4443 => x"52",
          4444 => x"08",
          4445 => x"88",
          4446 => x"08",
          4447 => x"38",
          4448 => x"2a",
          4449 => x"81",
          4450 => x"3d",
          4451 => x"82",
          4452 => x"e0",
          4453 => x"e0",
          4454 => x"83",
          4455 => x"ff",
          4456 => x"54",
          4457 => x"82",
          4458 => x"b2",
          4459 => x"82",
          4460 => x"53",
          4461 => x"c6",
          4462 => x"34",
          4463 => x"34",
          4464 => x"19",
          4465 => x"78",
          4466 => x"3f",
          4467 => x"d8",
          4468 => x"54",
          4469 => x"53",
          4470 => x"b7",
          4471 => x"15",
          4472 => x"82",
          4473 => x"08",
          4474 => x"64",
          4475 => x"75",
          4476 => x"9d",
          4477 => x"34",
          4478 => x"78",
          4479 => x"98",
          4480 => x"52",
          4481 => x"82",
          4482 => x"d8",
          4483 => x"d1",
          4484 => x"fc",
          4485 => x"3f",
          4486 => x"98",
          4487 => x"3d",
          4488 => x"c8",
          4489 => x"82",
          4490 => x"81",
          4491 => x"86",
          4492 => x"a5",
          4493 => x"05",
          4494 => x"77",
          4495 => x"a2",
          4496 => x"51",
          4497 => x"55",
          4498 => x"a1",
          4499 => x"38",
          4500 => x"88",
          4501 => x"08",
          4502 => x"38",
          4503 => x"e0",
          4504 => x"81",
          4505 => x"3d",
          4506 => x"ff",
          4507 => x"8b",
          4508 => x"2a",
          4509 => x"89",
          4510 => x"17",
          4511 => x"34",
          4512 => x"81",
          4513 => x"80",
          4514 => x"38",
          4515 => x"3f",
          4516 => x"ff",
          4517 => x"98",
          4518 => x"e0",
          4519 => x"9e",
          4520 => x"d8",
          4521 => x"08",
          4522 => x"73",
          4523 => x"63",
          4524 => x"9d",
          4525 => x"34",
          4526 => x"38",
          4527 => x"98",
          4528 => x"38",
          4529 => x"e0",
          4530 => x"0c",
          4531 => x"02",
          4532 => x"80",
          4533 => x"96",
          4534 => x"d1",
          4535 => x"82",
          4536 => x"5a",
          4537 => x"c5",
          4538 => x"82",
          4539 => x"cf",
          4540 => x"55",
          4541 => x"71",
          4542 => x"74",
          4543 => x"8b",
          4544 => x"15",
          4545 => x"82",
          4546 => x"98",
          4547 => x"0d",
          4548 => x"05",
          4549 => x"82",
          4550 => x"08",
          4551 => x"94",
          4552 => x"82",
          4553 => x"08",
          4554 => x"81",
          4555 => x"38",
          4556 => x"90",
          4557 => x"ff",
          4558 => x"83",
          4559 => x"3f",
          4560 => x"e0",
          4561 => x"3d",
          4562 => x"99",
          4563 => x"cf",
          4564 => x"e0",
          4565 => x"08",
          4566 => x"80",
          4567 => x"06",
          4568 => x"38",
          4569 => x"3d",
          4570 => x"82",
          4571 => x"08",
          4572 => x"ff",
          4573 => x"57",
          4574 => x"e0",
          4575 => x"5b",
          4576 => x"18",
          4577 => x"81",
          4578 => x"8b",
          4579 => x"75",
          4580 => x"1b",
          4581 => x"2e",
          4582 => x"09",
          4583 => x"80",
          4584 => x"25",
          4585 => x"38",
          4586 => x"11",
          4587 => x"82",
          4588 => x"08",
          4589 => x"80",
          4590 => x"80",
          4591 => x"a7",
          4592 => x"9b",
          4593 => x"0c",
          4594 => x"0d",
          4595 => x"3d",
          4596 => x"cd",
          4597 => x"e0",
          4598 => x"08",
          4599 => x"8a",
          4600 => x"3f",
          4601 => x"9f",
          4602 => x"9d",
          4603 => x"e0",
          4604 => x"c4",
          4605 => x"c0",
          4606 => x"08",
          4607 => x"08",
          4608 => x"2e",
          4609 => x"51",
          4610 => x"08",
          4611 => x"38",
          4612 => x"8a",
          4613 => x"e7",
          4614 => x"74",
          4615 => x"05",
          4616 => x"70",
          4617 => x"70",
          4618 => x"fe",
          4619 => x"55",
          4620 => x"75",
          4621 => x"55",
          4622 => x"a0",
          4623 => x"16",
          4624 => x"42",
          4625 => x"ff",
          4626 => x"54",
          4627 => x"81",
          4628 => x"82",
          4629 => x"08",
          4630 => x"54",
          4631 => x"e0",
          4632 => x"80",
          4633 => x"80",
          4634 => x"ab",
          4635 => x"82",
          4636 => x"82",
          4637 => x"99",
          4638 => x"15",
          4639 => x"ff",
          4640 => x"83",
          4641 => x"3f",
          4642 => x"74",
          4643 => x"04",
          4644 => x"05",
          4645 => x"05",
          4646 => x"b9",
          4647 => x"e0",
          4648 => x"33",
          4649 => x"2e",
          4650 => x"90",
          4651 => x"70",
          4652 => x"38",
          4653 => x"82",
          4654 => x"7e",
          4655 => x"55",
          4656 => x"cb",
          4657 => x"70",
          4658 => x"08",
          4659 => x"5d",
          4660 => x"9c",
          4661 => x"57",
          4662 => x"52",
          4663 => x"15",
          4664 => x"26",
          4665 => x"08",
          4666 => x"98",
          4667 => x"e0",
          4668 => x"75",
          4669 => x"93",
          4670 => x"2e",
          4671 => x"58",
          4672 => x"38",
          4673 => x"b4",
          4674 => x"09",
          4675 => x"53",
          4676 => x"3f",
          4677 => x"98",
          4678 => x"ff",
          4679 => x"84",
          4680 => x"12",
          4681 => x"78",
          4682 => x"90",
          4683 => x"90",
          4684 => x"94",
          4685 => x"91",
          4686 => x"84",
          4687 => x"16",
          4688 => x"0c",
          4689 => x"6c",
          4690 => x"33",
          4691 => x"d1",
          4692 => x"98",
          4693 => x"98",
          4694 => x"70",
          4695 => x"38",
          4696 => x"82",
          4697 => x"11",
          4698 => x"41",
          4699 => x"ac",
          4700 => x"06",
          4701 => x"74",
          4702 => x"81",
          4703 => x"cc",
          4704 => x"52",
          4705 => x"e0",
          4706 => x"80",
          4707 => x"26",
          4708 => x"74",
          4709 => x"80",
          4710 => x"92",
          4711 => x"38",
          4712 => x"2e",
          4713 => x"78",
          4714 => x"2b",
          4715 => x"38",
          4716 => x"77",
          4717 => x"dc",
          4718 => x"81",
          4719 => x"ff",
          4720 => x"98",
          4721 => x"51",
          4722 => x"08",
          4723 => x"74",
          4724 => x"8b",
          4725 => x"b2",
          4726 => x"8b",
          4727 => x"92",
          4728 => x"ba",
          4729 => x"82",
          4730 => x"3d",
          4731 => x"ff",
          4732 => x"98",
          4733 => x"70",
          4734 => x"51",
          4735 => x"55",
          4736 => x"38",
          4737 => x"ff",
          4738 => x"78",
          4739 => x"81",
          4740 => x"80",
          4741 => x"74",
          4742 => x"06",
          4743 => x"62",
          4744 => x"74",
          4745 => x"7d",
          4746 => x"38",
          4747 => x"81",
          4748 => x"74",
          4749 => x"98",
          4750 => x"82",
          4751 => x"80",
          4752 => x"38",
          4753 => x"3f",
          4754 => x"87",
          4755 => x"5c",
          4756 => x"80",
          4757 => x"0a",
          4758 => x"39",
          4759 => x"81",
          4760 => x"74",
          4761 => x"98",
          4762 => x"82",
          4763 => x"80",
          4764 => x"38",
          4765 => x"3f",
          4766 => x"57",
          4767 => x"96",
          4768 => x"10",
          4769 => x"72",
          4770 => x"ff",
          4771 => x"46",
          4772 => x"70",
          4773 => x"06",
          4774 => x"41",
          4775 => x"38",
          4776 => x"39",
          4777 => x"70",
          4778 => x"76",
          4779 => x"7d",
          4780 => x"55",
          4781 => x"08",
          4782 => x"9b",
          4783 => x"f5",
          4784 => x"38",
          4785 => x"38",
          4786 => x"81",
          4787 => x"0b",
          4788 => x"78",
          4789 => x"c0",
          4790 => x"39",
          4791 => x"8f",
          4792 => x"e0",
          4793 => x"78",
          4794 => x"80",
          4795 => x"39",
          4796 => x"06",
          4797 => x"27",
          4798 => x"56",
          4799 => x"80",
          4800 => x"8b",
          4801 => x"ff",
          4802 => x"1b",
          4803 => x"1c",
          4804 => x"8e",
          4805 => x"0b",
          4806 => x"30",
          4807 => x"51",
          4808 => x"3f",
          4809 => x"90",
          4810 => x"93",
          4811 => x"39",
          4812 => x"fc",
          4813 => x"52",
          4814 => x"81",
          4815 => x"c6",
          4816 => x"8d",
          4817 => x"06",
          4818 => x"52",
          4819 => x"3f",
          4820 => x"bc",
          4821 => x"8d",
          4822 => x"ff",
          4823 => x"51",
          4824 => x"80",
          4825 => x"1c",
          4826 => x"80",
          4827 => x"b2",
          4828 => x"fc",
          4829 => x"96",
          4830 => x"80",
          4831 => x"1c",
          4832 => x"ab",
          4833 => x"d4",
          4834 => x"59",
          4835 => x"53",
          4836 => x"3f",
          4837 => x"9c",
          4838 => x"80",
          4839 => x"7a",
          4840 => x"84",
          4841 => x"8c",
          4842 => x"52",
          4843 => x"8a",
          4844 => x"51",
          4845 => x"83",
          4846 => x"82",
          4847 => x"e4",
          4848 => x"ff",
          4849 => x"53",
          4850 => x"3f",
          4851 => x"7f",
          4852 => x"80",
          4853 => x"60",
          4854 => x"81",
          4855 => x"ff",
          4856 => x"51",
          4857 => x"88",
          4858 => x"f8",
          4859 => x"55",
          4860 => x"3f",
          4861 => x"83",
          4862 => x"7a",
          4863 => x"82",
          4864 => x"80",
          4865 => x"51",
          4866 => x"78",
          4867 => x"18",
          4868 => x"79",
          4869 => x"55",
          4870 => x"74",
          4871 => x"7f",
          4872 => x"98",
          4873 => x"78",
          4874 => x"57",
          4875 => x"67",
          4876 => x"57",
          4877 => x"64",
          4878 => x"53",
          4879 => x"3f",
          4880 => x"c4",
          4881 => x"83",
          4882 => x"98",
          4883 => x"85",
          4884 => x"2a",
          4885 => x"84",
          4886 => x"89",
          4887 => x"51",
          4888 => x"55",
          4889 => x"34",
          4890 => x"16",
          4891 => x"56",
          4892 => x"93",
          4893 => x"82",
          4894 => x"56",
          4895 => x"08",
          4896 => x"1b",
          4897 => x"83",
          4898 => x"81",
          4899 => x"ff",
          4900 => x"98",
          4901 => x"7f",
          4902 => x"82",
          4903 => x"8e",
          4904 => x"82",
          4905 => x"98",
          4906 => x"0d",
          4907 => x"ff",
          4908 => x"b4",
          4909 => x"81",
          4910 => x"94",
          4911 => x"9c",
          4912 => x"2e",
          4913 => x"58",
          4914 => x"09",
          4915 => x"78",
          4916 => x"82",
          4917 => x"f7",
          4918 => x"05",
          4919 => x"81",
          4920 => x"e7",
          4921 => x"24",
          4922 => x"8c",
          4923 => x"16",
          4924 => x"3d",
          4925 => x"52",
          4926 => x"76",
          4927 => x"2a",
          4928 => x"84",
          4929 => x"8b",
          4930 => x"84",
          4931 => x"a7",
          4932 => x"53",
          4933 => x"dc",
          4934 => x"84",
          4935 => x"87",
          4936 => x"ff",
          4937 => x"3d",
          4938 => x"80",
          4939 => x"86",
          4940 => x"0d",
          4941 => x"05",
          4942 => x"54",
          4943 => x"fe",
          4944 => x"98",
          4945 => x"02",
          4946 => x"80",
          4947 => x"72",
          4948 => x"39",
          4949 => x"83",
          4950 => x"70",
          4951 => x"22",
          4952 => x"12",
          4953 => x"71",
          4954 => x"82",
          4955 => x"e1",
          4956 => x"06",
          4957 => x"85",
          4958 => x"92",
          4959 => x"22",
          4960 => x"26",
          4961 => x"83",
          4962 => x"70",
          4963 => x"82",
          4964 => x"72",
          4965 => x"04",
          4966 => x"ff",
          4967 => x"ff",
          4968 => x"9f",
          4969 => x"e0",
          4970 => x"70",
          4971 => x"07",
          4972 => x"75",
          4973 => x"2a",
          4974 => x"52",
          4975 => x"38",
          4976 => x"84",
          4977 => x"08",
          4978 => x"70",
          4979 => x"71",
          4980 => x"51",
          4981 => x"39",
          4982 => x"51",
          4983 => x"88",
          4984 => x"51",
          4985 => x"83",
          4986 => x"fe",
          4987 => x"f1",
          4988 => x"0c",
          4989 => x"ff",
          4990 => x"ff",
          4991 => x"01",
          4992 => x"8c",
          4993 => x"9a",
          4994 => x"a8",
          4995 => x"b6",
          4996 => x"c4",
          4997 => x"d1",
          4998 => x"dd",
          4999 => x"e9",
          5000 => x"f5",
          5001 => x"81",
          5002 => x"8d",
          5003 => x"99",
          5004 => x"79",
          5005 => x"e2",
          5006 => x"4c",
          5007 => x"b3",
          5008 => x"2b",
          5009 => x"34",
          5010 => x"8a",
          5011 => x"52",
          5012 => x"4c",
          5013 => x"2b",
          5014 => x"e2",
          5015 => x"9f",
          5016 => x"b0",
          5017 => x"ba",
          5018 => x"c4",
          5019 => x"65",
          5020 => x"4e",
          5021 => x"4e",
          5022 => x"4e",
          5023 => x"4e",
          5024 => x"4e",
          5025 => x"4e",
          5026 => x"ac",
          5027 => x"4e",
          5028 => x"4e",
          5029 => x"4e",
          5030 => x"4e",
          5031 => x"4e",
          5032 => x"4e",
          5033 => x"4e",
          5034 => x"4e",
          5035 => x"4e",
          5036 => x"4e",
          5037 => x"4e",
          5038 => x"4e",
          5039 => x"4e",
          5040 => x"4e",
          5041 => x"4e",
          5042 => x"4e",
          5043 => x"4e",
          5044 => x"4e",
          5045 => x"4e",
          5046 => x"4e",
          5047 => x"4a",
          5048 => x"4e",
          5049 => x"4e",
          5050 => x"4e",
          5051 => x"4e",
          5052 => x"4e",
          5053 => x"73",
          5054 => x"e3",
          5055 => x"4e",
          5056 => x"4e",
          5057 => x"cc",
          5058 => x"4e",
          5059 => x"2b",
          5060 => x"4e",
          5061 => x"4e",
          5062 => x"4e",
          5063 => x"4a",
          5064 => x"00",
          5065 => x"00",
          5066 => x"00",
          5067 => x"00",
          5068 => x"00",
          5069 => x"00",
          5070 => x"00",
          5071 => x"00",
          5072 => x"00",
          5073 => x"00",
          5074 => x"00",
          5075 => x"00",
          5076 => x"6c",
          5077 => x"00",
          5078 => x"00",
          5079 => x"00",
          5080 => x"00",
          5081 => x"00",
          5082 => x"00",
          5083 => x"00",
          5084 => x"6b",
          5085 => x"00",
          5086 => x"6c",
          5087 => x"00",
          5088 => x"74",
          5089 => x"00",
          5090 => x"20",
          5091 => x"00",
          5092 => x"20",
          5093 => x"00",
          5094 => x"20",
          5095 => x"65",
          5096 => x"65",
          5097 => x"65",
          5098 => x"65",
          5099 => x"79",
          5100 => x"2e",
          5101 => x"65",
          5102 => x"20",
          5103 => x"2e",
          5104 => x"69",
          5105 => x"20",
          5106 => x"65",
          5107 => x"76",
          5108 => x"72",
          5109 => x"61",
          5110 => x"00",
          5111 => x"74",
          5112 => x"64",
          5113 => x"63",
          5114 => x"6c",
          5115 => x"79",
          5116 => x"75",
          5117 => x"69",
          5118 => x"6d",
          5119 => x"74",
          5120 => x"65",
          5121 => x"65",
          5122 => x"63",
          5123 => x"64",
          5124 => x"65",
          5125 => x"6b",
          5126 => x"75",
          5127 => x"74",
          5128 => x"2e",
          5129 => x"20",
          5130 => x"65",
          5131 => x"2e",
          5132 => x"61",
          5133 => x"69",
          5134 => x"74",
          5135 => x"63",
          5136 => x"00",
          5137 => x"20",
          5138 => x"00",
          5139 => x"74",
          5140 => x"74",
          5141 => x"74",
          5142 => x"0a",
          5143 => x"64",
          5144 => x"6c",
          5145 => x"00",
          5146 => x"00",
          5147 => x"20",
          5148 => x"58",
          5149 => x"00",
          5150 => x"00",
          5151 => x"25",
          5152 => x"31",
          5153 => x"00",
          5154 => x"00",
          5155 => x"65",
          5156 => x"20",
          5157 => x"2a",
          5158 => x"20",
          5159 => x"70",
          5160 => x"65",
          5161 => x"65",
          5162 => x"72",
          5163 => x"20",
          5164 => x"70",
          5165 => x"54",
          5166 => x"74",
          5167 => x"00",
          5168 => x"52",
          5169 => x"75",
          5170 => x"54",
          5171 => x"74",
          5172 => x"00",
          5173 => x"58",
          5174 => x"75",
          5175 => x"54",
          5176 => x"74",
          5177 => x"00",
          5178 => x"58",
          5179 => x"75",
          5180 => x"74",
          5181 => x"74",
          5182 => x"00",
          5183 => x"67",
          5184 => x"2e",
          5185 => x"6f",
          5186 => x"74",
          5187 => x"5f",
          5188 => x"00",
          5189 => x"6c",
          5190 => x"6e",
          5191 => x"65",
          5192 => x"64",
          5193 => x"61",
          5194 => x"20",
          5195 => x"79",
          5196 => x"00",
          5197 => x"67",
          5198 => x"00",
          5199 => x"2e",
          5200 => x"70",
          5201 => x"2e",
          5202 => x"6c",
          5203 => x"2d",
          5204 => x"25",
          5205 => x"00",
          5206 => x"6d",
          5207 => x"6d",
          5208 => x"00",
          5209 => x"30",
          5210 => x"00",
          5211 => x"30",
          5212 => x"6c",
          5213 => x"2d",
          5214 => x"63",
          5215 => x"6f",
          5216 => x"38",
          5217 => x"00",
          5218 => x"20",
          5219 => x"25",
          5220 => x"2e",
          5221 => x"6c",
          5222 => x"65",
          5223 => x"28",
          5224 => x"00",
          5225 => x"69",
          5226 => x"69",
          5227 => x"2e",
          5228 => x"64",
          5229 => x"69",
          5230 => x"00",
          5231 => x"00",
          5232 => x"25",
          5233 => x"00",
          5234 => x"25",
          5235 => x"5c",
          5236 => x"20",
          5237 => x"2e",
          5238 => x"6f",
          5239 => x"75",
          5240 => x"61",
          5241 => x"6f",
          5242 => x"6d",
          5243 => x"00",
          5244 => x"2e",
          5245 => x"62",
          5246 => x"74",
          5247 => x"2e",
          5248 => x"25",
          5249 => x"3a",
          5250 => x"64",
          5251 => x"20",
          5252 => x"72",
          5253 => x"00",
          5254 => x"53",
          5255 => x"69",
          5256 => x"65",
          5257 => x"6d",
          5258 => x"65",
          5259 => x"20",
          5260 => x"4d",
          5261 => x"3a",
          5262 => x"00",
          5263 => x"41",
          5264 => x"25",
          5265 => x"58",
          5266 => x"20",
          5267 => x"41",
          5268 => x"3a",
          5269 => x"00",
          5270 => x"4d",
          5271 => x"25",
          5272 => x"58",
          5273 => x"20",
          5274 => x"20",
          5275 => x"3a",
          5276 => x"00",
          5277 => x"43",
          5278 => x"44",
          5279 => x"3d",
          5280 => x"00",
          5281 => x"45",
          5282 => x"54",
          5283 => x"3d",
          5284 => x"00",
          5285 => x"52",
          5286 => x"43",
          5287 => x"3d",
          5288 => x"00",
          5289 => x"48",
          5290 => x"53",
          5291 => x"20",
          5292 => x"00",
          5293 => x"54",
          5294 => x"20",
          5295 => x"20",
          5296 => x"72",
          5297 => x"00",
          5298 => x"20",
          5299 => x"65",
          5300 => x"64",
          5301 => x"25",
          5302 => x"00",
          5303 => x"20",
          5304 => x"53",
          5305 => x"64",
          5306 => x"25",
          5307 => x"00",
          5308 => x"63",
          5309 => x"20",
          5310 => x"20",
          5311 => x"25",
          5312 => x"00",
          5313 => x"00",
          5314 => x"20",
          5315 => x"20",
          5316 => x"20",
          5317 => x"25",
          5318 => x"00",
          5319 => x"74",
          5320 => x"6b",
          5321 => x"20",
          5322 => x"25",
          5323 => x"48",
          5324 => x"20",
          5325 => x"6c",
          5326 => x"71",
          5327 => x"20",
          5328 => x"30",
          5329 => x"00",
          5330 => x"68",
          5331 => x"52",
          5332 => x"6b",
          5333 => x"25",
          5334 => x"48",
          5335 => x"6c",
          5336 => x"69",
          5337 => x"78",
          5338 => x"00",
          5339 => x"00",
          5340 => x"00",
          5341 => x"00",
          5342 => x"40",
          5343 => x"03",
          5344 => x"00",
          5345 => x"38",
          5346 => x"05",
          5347 => x"00",
          5348 => x"30",
          5349 => x"07",
          5350 => x"00",
          5351 => x"28",
          5352 => x"08",
          5353 => x"00",
          5354 => x"20",
          5355 => x"09",
          5356 => x"00",
          5357 => x"18",
          5358 => x"0d",
          5359 => x"00",
          5360 => x"10",
          5361 => x"0e",
          5362 => x"00",
          5363 => x"08",
          5364 => x"0f",
          5365 => x"00",
          5366 => x"00",
          5367 => x"11",
          5368 => x"00",
          5369 => x"f8",
          5370 => x"13",
          5371 => x"00",
          5372 => x"f0",
          5373 => x"15",
          5374 => x"00",
          5375 => x"00",
          5376 => x"7e",
          5377 => x"00",
          5378 => x"7e",
          5379 => x"00",
          5380 => x"00",
          5381 => x"00",
          5382 => x"00",
          5383 => x"00",
          5384 => x"00",
          5385 => x"00",
          5386 => x"00",
          5387 => x"6c",
          5388 => x"00",
          5389 => x"74",
          5390 => x"20",
          5391 => x"74",
          5392 => x"65",
          5393 => x"2e",
          5394 => x"6e",
          5395 => x"2f",
          5396 => x"68",
          5397 => x"66",
          5398 => x"73",
          5399 => x"00",
          5400 => x"3c",
          5401 => x"00",
          5402 => x"00",
          5403 => x"33",
          5404 => x"4d",
          5405 => x"00",
          5406 => x"20",
          5407 => x"32",
          5408 => x"4e",
          5409 => x"46",
          5410 => x"00",
          5411 => x"00",
          5412 => x"00",
          5413 => x"12",
          5414 => x"00",
          5415 => x"80",
          5416 => x"8f",
          5417 => x"55",
          5418 => x"9f",
          5419 => x"a7",
          5420 => x"af",
          5421 => x"b7",
          5422 => x"bf",
          5423 => x"c7",
          5424 => x"cf",
          5425 => x"d7",
          5426 => x"df",
          5427 => x"e7",
          5428 => x"ef",
          5429 => x"f7",
          5430 => x"ff",
          5431 => x"2f",
          5432 => x"7c",
          5433 => x"04",
          5434 => x"00",
          5435 => x"02",
          5436 => x"20",
          5437 => x"fc",
          5438 => x"e0",
          5439 => x"eb",
          5440 => x"ec",
          5441 => x"e6",
          5442 => x"f2",
          5443 => x"d6",
          5444 => x"a5",
          5445 => x"ed",
          5446 => x"d1",
          5447 => x"10",
          5448 => x"a1",
          5449 => x"92",
          5450 => x"61",
          5451 => x"63",
          5452 => x"5c",
          5453 => x"34",
          5454 => x"3c",
          5455 => x"54",
          5456 => x"50",
          5457 => x"64",
          5458 => x"52",
          5459 => x"18",
          5460 => x"8c",
          5461 => x"df",
          5462 => x"c3",
          5463 => x"98",
          5464 => x"c6",
          5465 => x"b1",
          5466 => x"21",
          5467 => x"19",
          5468 => x"b2",
          5469 => x"1a",
          5470 => x"07",
          5471 => x"00",
          5472 => x"39",
          5473 => x"79",
          5474 => x"43",
          5475 => x"84",
          5476 => x"87",
          5477 => x"8b",
          5478 => x"90",
          5479 => x"94",
          5480 => x"98",
          5481 => x"9c",
          5482 => x"a0",
          5483 => x"a4",
          5484 => x"a7",
          5485 => x"ac",
          5486 => x"af",
          5487 => x"b3",
          5488 => x"b8",
          5489 => x"bc",
          5490 => x"c0",
          5491 => x"c4",
          5492 => x"c8",
          5493 => x"ca",
          5494 => x"01",
          5495 => x"f3",
          5496 => x"f4",
          5497 => x"12",
          5498 => x"3b",
          5499 => x"3f",
          5500 => x"46",
          5501 => x"81",
          5502 => x"8a",
          5503 => x"90",
          5504 => x"5f",
          5505 => x"94",
          5506 => x"67",
          5507 => x"62",
          5508 => x"9c",
          5509 => x"73",
          5510 => x"77",
          5511 => x"7b",
          5512 => x"7f",
          5513 => x"a9",
          5514 => x"87",
          5515 => x"b2",
          5516 => x"8f",
          5517 => x"7b",
          5518 => x"ff",
          5519 => x"88",
          5520 => x"11",
          5521 => x"a3",
          5522 => x"03",
          5523 => x"d8",
          5524 => x"f9",
          5525 => x"f6",
          5526 => x"fa",
          5527 => x"50",
          5528 => x"8a",
          5529 => x"cf",
          5530 => x"44",
          5531 => x"00",
          5532 => x"00",
          5533 => x"00",
          5534 => x"20",
          5535 => x"40",
          5536 => x"59",
          5537 => x"5d",
          5538 => x"08",
          5539 => x"bb",
          5540 => x"cb",
          5541 => x"f9",
          5542 => x"fb",
          5543 => x"08",
          5544 => x"04",
          5545 => x"bc",
          5546 => x"d0",
          5547 => x"e5",
          5548 => x"01",
          5549 => x"32",
          5550 => x"01",
          5551 => x"30",
          5552 => x"67",
          5553 => x"80",
          5554 => x"41",
          5555 => x"00",
          5556 => x"00",
          5557 => x"00",
          5558 => x"00",
          5559 => x"00",
          5560 => x"00",
          5561 => x"00",
          5562 => x"00",
          5563 => x"00",
          5564 => x"00",
          5565 => x"00",
          5566 => x"00",
          5567 => x"00",
          5568 => x"00",
          5569 => x"00",
          5570 => x"00",
          5571 => x"00",
          5572 => x"00",
          5573 => x"00",
          5574 => x"00",
          5575 => x"00",
          5576 => x"00",
          5577 => x"00",
          5578 => x"00",
          5579 => x"00",
          5580 => x"00",
          5581 => x"00",
          5582 => x"00",
          5583 => x"00",
          5584 => x"00",
          5585 => x"00",
          5586 => x"00",
          5587 => x"00",
          5588 => x"00",
          5589 => x"00",
          5590 => x"00",
          5591 => x"00",
          5592 => x"00",
          5593 => x"00",
          5594 => x"00",
          5595 => x"00",
          5596 => x"00",
          5597 => x"00",
          5598 => x"00",
          5599 => x"00",
          5600 => x"00",
          5601 => x"00",
          5602 => x"00",
          5603 => x"00",
          5604 => x"00",
          5605 => x"00",
          5606 => x"00",
          5607 => x"00",
          5608 => x"00",
          5609 => x"00",
          5610 => x"00",
          5611 => x"00",
          5612 => x"00",
          5613 => x"00",
          5614 => x"00",
          5615 => x"01",
          5616 => x"01",
          5617 => x"00",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"48",
          5630 => x"50",
          5631 => x"58",
          5632 => x"00",
          5633 => x"02",
          5634 => x"00",
        others => X"00"
    );

    shared variable RAM5 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"88",
             5 => x"88",
             6 => x"00",
             7 => x"00",
             8 => x"06",
             9 => x"2a",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"05",
            14 => x"ff",
            15 => x"04",
            16 => x"73",
            17 => x"73",
            18 => x"04",
            19 => x"00",
            20 => x"07",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"81",
            25 => x"0a",
            26 => x"81",
            27 => x"00",
            28 => x"07",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"00",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"51",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"05",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"06",
            49 => x"ff",
            50 => x"00",
            51 => x"00",
            52 => x"73",
            53 => x"83",
            54 => x"0c",
            55 => x"00",
            56 => x"09",
            57 => x"06",
            58 => x"00",
            59 => x"00",
            60 => x"09",
            61 => x"81",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"53",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"09",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"06",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"82",
            81 => x"05",
            82 => x"04",
            83 => x"00",
            84 => x"75",
            85 => x"50",
            86 => x"0c",
            87 => x"00",
            88 => x"75",
            89 => x"50",
            90 => x"0c",
            91 => x"00",
            92 => x"06",
            93 => x"71",
            94 => x"05",
            95 => x"00",
            96 => x"06",
            97 => x"54",
            98 => x"ff",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"05",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"53",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"0b",
           133 => x"0b",
           134 => x"a6",
           135 => x"0b",
           136 => x"0b",
           137 => x"e6",
           138 => x"0b",
           139 => x"0b",
           140 => x"a8",
           141 => x"0b",
           142 => x"0b",
           143 => x"eb",
           144 => x"0b",
           145 => x"0b",
           146 => x"af",
           147 => x"0b",
           148 => x"0b",
           149 => x"f3",
           150 => x"0b",
           151 => x"0b",
           152 => x"b7",
           153 => x"0b",
           154 => x"0b",
           155 => x"fb",
           156 => x"0b",
           157 => x"0b",
           158 => x"bf",
           159 => x"0b",
           160 => x"0b",
           161 => x"83",
           162 => x"0b",
           163 => x"0b",
           164 => x"c7",
           165 => x"0b",
           166 => x"0b",
           167 => x"8b",
           168 => x"0b",
           169 => x"0b",
           170 => x"cf",
           171 => x"0b",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"e0",
           193 => x"e0",
           194 => x"82",
           195 => x"e0",
           196 => x"82",
           197 => x"e0",
           198 => x"82",
           199 => x"e0",
           200 => x"82",
           201 => x"e0",
           202 => x"82",
           203 => x"e0",
           204 => x"82",
           205 => x"82",
           206 => x"04",
           207 => x"2d",
           208 => x"90",
           209 => x"2d",
           210 => x"90",
           211 => x"2d",
           212 => x"90",
           213 => x"2d",
           214 => x"90",
           215 => x"e7",
           216 => x"80",
           217 => x"ff",
           218 => x"c0",
           219 => x"81",
           220 => x"80",
           221 => x"0c",
           222 => x"08",
           223 => x"a4",
           224 => x"a4",
           225 => x"e0",
           226 => x"e0",
           227 => x"82",
           228 => x"82",
           229 => x"04",
           230 => x"2d",
           231 => x"90",
           232 => x"8c",
           233 => x"80",
           234 => x"88",
           235 => x"c0",
           236 => x"82",
           237 => x"80",
           238 => x"0c",
           239 => x"08",
           240 => x"a4",
           241 => x"a4",
           242 => x"e0",
           243 => x"e0",
           244 => x"82",
           245 => x"82",
           246 => x"04",
           247 => x"2d",
           248 => x"90",
           249 => x"9d",
           250 => x"80",
           251 => x"98",
           252 => x"c0",
           253 => x"82",
           254 => x"80",
           255 => x"0c",
           256 => x"08",
           257 => x"a4",
           258 => x"a4",
           259 => x"e0",
           260 => x"e0",
           261 => x"82",
           262 => x"82",
           263 => x"04",
           264 => x"2d",
           265 => x"90",
           266 => x"a4",
           267 => x"80",
           268 => x"9d",
           269 => x"c0",
           270 => x"82",
           271 => x"80",
           272 => x"0c",
           273 => x"08",
           274 => x"a4",
           275 => x"a4",
           276 => x"e0",
           277 => x"e0",
           278 => x"82",
           279 => x"82",
           280 => x"04",
           281 => x"2d",
           282 => x"90",
           283 => x"8b",
           284 => x"80",
           285 => x"b6",
           286 => x"c0",
           287 => x"81",
           288 => x"80",
           289 => x"0c",
           290 => x"08",
           291 => x"a4",
           292 => x"a4",
           293 => x"e0",
           294 => x"e0",
           295 => x"82",
           296 => x"82",
           297 => x"04",
           298 => x"2d",
           299 => x"90",
           300 => x"c7",
           301 => x"80",
           302 => x"b3",
           303 => x"c0",
           304 => x"81",
           305 => x"80",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"04",
           311 => x"83",
           312 => x"10",
           313 => x"51",
           314 => x"06",
           315 => x"10",
           316 => x"ed",
           317 => x"e0",
           318 => x"38",
           319 => x"0b",
           320 => x"51",
           321 => x"a4",
           322 => x"3d",
           323 => x"70",
           324 => x"82",
           325 => x"82",
           326 => x"82",
           327 => x"3f",
           328 => x"a4",
           329 => x"08",
           330 => x"0c",
           331 => x"a4",
           332 => x"82",
           333 => x"e0",
           334 => x"33",
           335 => x"51",
           336 => x"82",
           337 => x"83",
           338 => x"a4",
           339 => x"82",
           340 => x"05",
           341 => x"80",
           342 => x"0c",
           343 => x"82",
           344 => x"e0",
           345 => x"80",
           346 => x"08",
           347 => x"82",
           348 => x"a0",
           349 => x"82",
           350 => x"82",
           351 => x"2e",
           352 => x"82",
           353 => x"d2",
           354 => x"08",
           355 => x"53",
           356 => x"08",
           357 => x"a4",
           358 => x"08",
           359 => x"a4",
           360 => x"82",
           361 => x"80",
           362 => x"05",
           363 => x"05",
           364 => x"05",
           365 => x"0d",
           366 => x"a4",
           367 => x"3d",
           368 => x"e5",
           369 => x"05",
           370 => x"0c",
           371 => x"e8",
           372 => x"05",
           373 => x"0c",
           374 => x"54",
           375 => x"53",
           376 => x"53",
           377 => x"98",
           378 => x"05",
           379 => x"08",
           380 => x"05",
           381 => x"a4",
           382 => x"98",
           383 => x"a4",
           384 => x"82",
           385 => x"e0",
           386 => x"a4",
           387 => x"08",
           388 => x"08",
           389 => x"08",
           390 => x"82",
           391 => x"08",
           392 => x"f8",
           393 => x"51",
           394 => x"0c",
           395 => x"e0",
           396 => x"82",
           397 => x"e0",
           398 => x"0b",
           399 => x"88",
           400 => x"2a",
           401 => x"51",
           402 => x"38",
           403 => x"05",
           404 => x"08",
           405 => x"72",
           406 => x"72",
           407 => x"95",
           408 => x"05",
           409 => x"8c",
           410 => x"05",
           411 => x"80",
           412 => x"08",
           413 => x"81",
           414 => x"05",
           415 => x"38",
           416 => x"53",
           417 => x"c5",
           418 => x"33",
           419 => x"51",
           420 => x"08",
           421 => x"81",
           422 => x"53",
           423 => x"a4",
           424 => x"07",
           425 => x"e4",
           426 => x"a4",
           427 => x"70",
           428 => x"11",
           429 => x"55",
           430 => x"05",
           431 => x"33",
           432 => x"33",
           433 => x"72",
           434 => x"82",
           435 => x"98",
           436 => x"72",
           437 => x"82",
           438 => x"e0",
           439 => x"2a",
           440 => x"fd",
           441 => x"05",
           442 => x"70",
           443 => x"51",
           444 => x"ec",
           445 => x"a4",
           446 => x"70",
           447 => x"2e",
           448 => x"05",
           449 => x"51",
           450 => x"82",
           451 => x"e0",
           452 => x"82",
           453 => x"82",
           454 => x"d8",
           455 => x"08",
           456 => x"b9",
           457 => x"53",
           458 => x"05",
           459 => x"82",
           460 => x"e0",
           461 => x"07",
           462 => x"e4",
           463 => x"a4",
           464 => x"07",
           465 => x"e4",
           466 => x"a4",
           467 => x"07",
           468 => x"e4",
           469 => x"a4",
           470 => x"51",
           471 => x"05",
           472 => x"e8",
           473 => x"a4",
           474 => x"51",
           475 => x"05",
           476 => x"e0",
           477 => x"a4",
           478 => x"53",
           479 => x"23",
           480 => x"f8",
           481 => x"a4",
           482 => x"08",
           483 => x"a4",
           484 => x"53",
           485 => x"34",
           486 => x"ff",
           487 => x"08",
           488 => x"e0",
           489 => x"a4",
           490 => x"e0",
           491 => x"82",
           492 => x"e0",
           493 => x"2a",
           494 => x"72",
           495 => x"08",
           496 => x"72",
           497 => x"fc",
           498 => x"82",
           499 => x"a4",
           500 => x"e0",
           501 => x"8a",
           502 => x"82",
           503 => x"e0",
           504 => x"e0",
           505 => x"31",
           506 => x"ec",
           507 => x"a4",
           508 => x"08",
           509 => x"a4",
           510 => x"e0",
           511 => x"a4",
           512 => x"70",
           513 => x"80",
           514 => x"e8",
           515 => x"98",
           516 => x"05",
           517 => x"e0",
           518 => x"08",
           519 => x"a4",
           520 => x"3f",
           521 => x"e0",
           522 => x"a4",
           523 => x"a4",
           524 => x"54",
           525 => x"05",
           526 => x"08",
           527 => x"81",
           528 => x"a4",
           529 => x"08",
           530 => x"84",
           531 => x"0c",
           532 => x"05",
           533 => x"08",
           534 => x"90",
           535 => x"08",
           536 => x"a4",
           537 => x"a4",
           538 => x"08",
           539 => x"fc",
           540 => x"e0",
           541 => x"07",
           542 => x"e4",
           543 => x"05",
           544 => x"05",
           545 => x"22",
           546 => x"82",
           547 => x"af",
           548 => x"f4",
           549 => x"08",
           550 => x"51",
           551 => x"05",
           552 => x"08",
           553 => x"a4",
           554 => x"08",
           555 => x"81",
           556 => x"a4",
           557 => x"08",
           558 => x"84",
           559 => x"0c",
           560 => x"05",
           561 => x"08",
           562 => x"90",
           563 => x"08",
           564 => x"a4",
           565 => x"a4",
           566 => x"08",
           567 => x"e4",
           568 => x"72",
           569 => x"82",
           570 => x"f0",
           571 => x"05",
           572 => x"22",
           573 => x"71",
           574 => x"ca",
           575 => x"75",
           576 => x"08",
           577 => x"82",
           578 => x"33",
           579 => x"82",
           580 => x"72",
           581 => x"05",
           582 => x"53",
           583 => x"34",
           584 => x"05",
           585 => x"53",
           586 => x"34",
           587 => x"53",
           588 => x"73",
           589 => x"08",
           590 => x"05",
           591 => x"22",
           592 => x"05",
           593 => x"e0",
           594 => x"fc",
           595 => x"fc",
           596 => x"b2",
           597 => x"08",
           598 => x"74",
           599 => x"e0",
           600 => x"a4",
           601 => x"51",
           602 => x"e0",
           603 => x"51",
           604 => x"05",
           605 => x"22",
           606 => x"51",
           607 => x"82",
           608 => x"90",
           609 => x"0c",
           610 => x"90",
           611 => x"0c",
           612 => x"51",
           613 => x"95",
           614 => x"08",
           615 => x"08",
           616 => x"a4",
           617 => x"72",
           618 => x"82",
           619 => x"e0",
           620 => x"a4",
           621 => x"70",
           622 => x"2e",
           623 => x"e8",
           624 => x"2c",
           625 => x"57",
           626 => x"38",
           627 => x"70",
           628 => x"a4",
           629 => x"e0",
           630 => x"e0",
           631 => x"31",
           632 => x"e8",
           633 => x"05",
           634 => x"51",
           635 => x"82",
           636 => x"88",
           637 => x"70",
           638 => x"72",
           639 => x"22",
           640 => x"e0",
           641 => x"82",
           642 => x"88",
           643 => x"70",
           644 => x"72",
           645 => x"22",
           646 => x"e0",
           647 => x"a4",
           648 => x"06",
           649 => x"a4",
           650 => x"54",
           651 => x"23",
           652 => x"53",
           653 => x"a4",
           654 => x"8a",
           655 => x"08",
           656 => x"81",
           657 => x"91",
           658 => x"08",
           659 => x"c7",
           660 => x"22",
           661 => x"51",
           662 => x"e0",
           663 => x"51",
           664 => x"a4",
           665 => x"70",
           666 => x"2e",
           667 => x"05",
           668 => x"82",
           669 => x"86",
           670 => x"72",
           671 => x"08",
           672 => x"df",
           673 => x"22",
           674 => x"94",
           675 => x"08",
           676 => x"33",
           677 => x"08",
           678 => x"81",
           679 => x"b0",
           680 => x"22",
           681 => x"a4",
           682 => x"70",
           683 => x"90",
           684 => x"08",
           685 => x"39",
           686 => x"70",
           687 => x"53",
           688 => x"a4",
           689 => x"54",
           690 => x"34",
           691 => x"53",
           692 => x"a4",
           693 => x"88",
           694 => x"08",
           695 => x"81",
           696 => x"82",
           697 => x"11",
           698 => x"ec",
           699 => x"2c",
           700 => x"82",
           701 => x"a0",
           702 => x"e0",
           703 => x"80",
           704 => x"82",
           705 => x"82",
           706 => x"87",
           707 => x"a4",
           708 => x"f3",
           709 => x"82",
           710 => x"11",
           711 => x"f4",
           712 => x"53",
           713 => x"38",
           714 => x"52",
           715 => x"70",
           716 => x"05",
           717 => x"fc",
           718 => x"b7",
           719 => x"33",
           720 => x"06",
           721 => x"f4",
           722 => x"82",
           723 => x"83",
           724 => x"ff",
           725 => x"08",
           726 => x"08",
           727 => x"86",
           728 => x"05",
           729 => x"fc",
           730 => x"a4",
           731 => x"2e",
           732 => x"05",
           733 => x"05",
           734 => x"f0",
           735 => x"05",
           736 => x"3f",
           737 => x"05",
           738 => x"51",
           739 => x"38",
           740 => x"ff",
           741 => x"08",
           742 => x"90",
           743 => x"38",
           744 => x"52",
           745 => x"82",
           746 => x"82",
           747 => x"85",
           748 => x"08",
           749 => x"e0",
           750 => x"a5",
           751 => x"0b",
           752 => x"80",
           753 => x"23",
           754 => x"05",
           755 => x"f4",
           756 => x"a4",
           757 => x"a4",
           758 => x"3f",
           759 => x"88",
           760 => x"e0",
           761 => x"82",
           762 => x"e0",
           763 => x"a4",
           764 => x"82",
           765 => x"fb",
           766 => x"8c",
           767 => x"88",
           768 => x"e0",
           769 => x"54",
           770 => x"04",
           771 => x"a4",
           772 => x"e0",
           773 => x"fc",
           774 => x"70",
           775 => x"51",
           776 => x"ff",
           777 => x"0c",
           778 => x"88",
           779 => x"a4",
           780 => x"e0",
           781 => x"82",
           782 => x"81",
           783 => x"38",
           784 => x"08",
           785 => x"33",
           786 => x"2d",
           787 => x"2e",
           788 => x"a4",
           789 => x"82",
           790 => x"53",
           791 => x"72",
           792 => x"80",
           793 => x"a4",
           794 => x"08",
           795 => x"08",
           796 => x"08",
           797 => x"87",
           798 => x"82",
           799 => x"0c",
           800 => x"a4",
           801 => x"08",
           802 => x"81",
           803 => x"51",
           804 => x"8d",
           805 => x"f4",
           806 => x"a4",
           807 => x"82",
           808 => x"05",
           809 => x"53",
           810 => x"34",
           811 => x"2e",
           812 => x"05",
           813 => x"08",
           814 => x"33",
           815 => x"2d",
           816 => x"2e",
           817 => x"a4",
           818 => x"82",
           819 => x"82",
           820 => x"82",
           821 => x"e0",
           822 => x"a4",
           823 => x"82",
           824 => x"fb",
           825 => x"88",
           826 => x"98",
           827 => x"84",
           828 => x"82",
           829 => x"0c",
           830 => x"8c",
           831 => x"2a",
           832 => x"51",
           833 => x"38",
           834 => x"05",
           835 => x"08",
           836 => x"82",
           837 => x"53",
           838 => x"e0",
           839 => x"a4",
           840 => x"14",
           841 => x"82",
           842 => x"08",
           843 => x"08",
           844 => x"73",
           845 => x"a4",
           846 => x"81",
           847 => x"08",
           848 => x"08",
           849 => x"39",
           850 => x"82",
           851 => x"82",
           852 => x"81",
           853 => x"54",
           854 => x"53",
           855 => x"8c",
           856 => x"8c",
           857 => x"05",
           858 => x"05",
           859 => x"82",
           860 => x"e0",
           861 => x"98",
           862 => x"0c",
           863 => x"e0",
           864 => x"a4",
           865 => x"70",
           866 => x"51",
           867 => x"0b",
           868 => x"83",
           869 => x"05",
           870 => x"70",
           871 => x"80",
           872 => x"08",
           873 => x"88",
           874 => x"70",
           875 => x"14",
           876 => x"08",
           877 => x"0c",
           878 => x"84",
           879 => x"f8",
           880 => x"39",
           881 => x"85",
           882 => x"06",
           883 => x"80",
           884 => x"05",
           885 => x"a4",
           886 => x"e0",
           887 => x"82",
           888 => x"e0",
           889 => x"85",
           890 => x"71",
           891 => x"a4",
           892 => x"82",
           893 => x"08",
           894 => x"39",
           895 => x"82",
           896 => x"94",
           897 => x"e0",
           898 => x"fc",
           899 => x"fc",
           900 => x"82",
           901 => x"e0",
           902 => x"a4",
           903 => x"82",
           904 => x"82",
           905 => x"2e",
           906 => x"a4",
           907 => x"71",
           908 => x"93",
           909 => x"08",
           910 => x"08",
           911 => x"f4",
           912 => x"ec",
           913 => x"82",
           914 => x"39",
           915 => x"8c",
           916 => x"82",
           917 => x"81",
           918 => x"f8",
           919 => x"a4",
           920 => x"0c",
           921 => x"04",
           922 => x"a4",
           923 => x"08",
           924 => x"fc",
           925 => x"05",
           926 => x"0c",
           927 => x"80",
           928 => x"08",
           929 => x"fc",
           930 => x"e0",
           931 => x"a4",
           932 => x"e0",
           933 => x"81",
           934 => x"05",
           935 => x"08",
           936 => x"0c",
           937 => x"82",
           938 => x"82",
           939 => x"e0",
           940 => x"82",
           941 => x"e0",
           942 => x"82",
           943 => x"e0",
           944 => x"81",
           945 => x"05",
           946 => x"fc",
           947 => x"05",
           948 => x"f8",
           949 => x"05",
           950 => x"08",
           951 => x"ae",
           952 => x"08",
           953 => x"05",
           954 => x"08",
           955 => x"05",
           956 => x"08",
           957 => x"08",
           958 => x"e0",
           959 => x"82",
           960 => x"e0",
           961 => x"71",
           962 => x"05",
           963 => x"fc",
           964 => x"a4",
           965 => x"98",
           966 => x"a4",
           967 => x"82",
           968 => x"e0",
           969 => x"a4",
           970 => x"08",
           971 => x"e0",
           972 => x"82",
           973 => x"81",
           974 => x"83",
           975 => x"fc",
           976 => x"08",
           977 => x"fc",
           978 => x"05",
           979 => x"51",
           980 => x"04",
           981 => x"a4",
           982 => x"08",
           983 => x"fc",
           984 => x"05",
           985 => x"08",
           986 => x"a4",
           987 => x"08",
           988 => x"34",
           989 => x"81",
           990 => x"0c",
           991 => x"2e",
           992 => x"a4",
           993 => x"98",
           994 => x"a4",
           995 => x"82",
           996 => x"e0",
           997 => x"a4",
           998 => x"08",
           999 => x"f8",
          1000 => x"05",
          1001 => x"e0",
          1002 => x"82",
          1003 => x"e0",
          1004 => x"82",
          1005 => x"e0",
          1006 => x"ba",
          1007 => x"08",
          1008 => x"f8",
          1009 => x"08",
          1010 => x"fc",
          1011 => x"82",
          1012 => x"05",
          1013 => x"ff",
          1014 => x"05",
          1015 => x"85",
          1016 => x"82",
          1017 => x"0c",
          1018 => x"90",
          1019 => x"82",
          1020 => x"71",
          1021 => x"08",
          1022 => x"05",
          1023 => x"08",
          1024 => x"54",
          1025 => x"80",
          1026 => x"05",
          1027 => x"08",
          1028 => x"a4",
          1029 => x"06",
          1030 => x"82",
          1031 => x"9b",
          1032 => x"08",
          1033 => x"05",
          1034 => x"08",
          1035 => x"82",
          1036 => x"2e",
          1037 => x"88",
          1038 => x"8d",
          1039 => x"fc",
          1040 => x"a4",
          1041 => x"e0",
          1042 => x"a4",
          1043 => x"52",
          1044 => x"a4",
          1045 => x"e0",
          1046 => x"82",
          1047 => x"33",
          1048 => x"08",
          1049 => x"53",
          1050 => x"08",
          1051 => x"fc",
          1052 => x"3d",
          1053 => x"e0",
          1054 => x"fa",
          1055 => x"05",
          1056 => x"05",
          1057 => x"98",
          1058 => x"05",
          1059 => x"08",
          1060 => x"ec",
          1061 => x"82",
          1062 => x"82",
          1063 => x"38",
          1064 => x"05",
          1065 => x"fc",
          1066 => x"05",
          1067 => x"e0",
          1068 => x"e0",
          1069 => x"e0",
          1070 => x"a2",
          1071 => x"e0",
          1072 => x"e0",
          1073 => x"98",
          1074 => x"0c",
          1075 => x"e0",
          1076 => x"a4",
          1077 => x"08",
          1078 => x"8c",
          1079 => x"e0",
          1080 => x"39",
          1081 => x"52",
          1082 => x"05",
          1083 => x"f8",
          1084 => x"51",
          1085 => x"a4",
          1086 => x"e0",
          1087 => x"a4",
          1088 => x"38",
          1089 => x"f8",
          1090 => x"08",
          1091 => x"f8",
          1092 => x"05",
          1093 => x"fc",
          1094 => x"fc",
          1095 => x"3d",
          1096 => x"e0",
          1097 => x"fe",
          1098 => x"05",
          1099 => x"0c",
          1100 => x"80",
          1101 => x"08",
          1102 => x"a4",
          1103 => x"08",
          1104 => x"a4",
          1105 => x"08",
          1106 => x"82",
          1107 => x"70",
          1108 => x"52",
          1109 => x"08",
          1110 => x"a4",
          1111 => x"82",
          1112 => x"82",
          1113 => x"82",
          1114 => x"08",
          1115 => x"0d",
          1116 => x"52",
          1117 => x"51",
          1118 => x"82",
          1119 => x"82",
          1120 => x"08",
          1121 => x"0d",
          1122 => x"05",
          1123 => x"08",
          1124 => x"08",
          1125 => x"82",
          1126 => x"08",
          1127 => x"e0",
          1128 => x"a4",
          1129 => x"08",
          1130 => x"82",
          1131 => x"83",
          1132 => x"e0",
          1133 => x"82",
          1134 => x"97",
          1135 => x"08",
          1136 => x"31",
          1137 => x"82",
          1138 => x"e0",
          1139 => x"a4",
          1140 => x"71",
          1141 => x"27",
          1142 => x"08",
          1143 => x"e0",
          1144 => x"52",
          1145 => x"08",
          1146 => x"e0",
          1147 => x"e0",
          1148 => x"af",
          1149 => x"08",
          1150 => x"05",
          1151 => x"08",
          1152 => x"2a",
          1153 => x"82",
          1154 => x"e0",
          1155 => x"e0",
          1156 => x"82",
          1157 => x"80",
          1158 => x"0c",
          1159 => x"80",
          1160 => x"08",
          1161 => x"08",
          1162 => x"a4",
          1163 => x"73",
          1164 => x"0c",
          1165 => x"10",
          1166 => x"08",
          1167 => x"0c",
          1168 => x"82",
          1169 => x"ff",
          1170 => x"08",
          1171 => x"a4",
          1172 => x"08",
          1173 => x"a4",
          1174 => x"08",
          1175 => x"ec",
          1176 => x"f4",
          1177 => x"08",
          1178 => x"f8",
          1179 => x"08",
          1180 => x"51",
          1181 => x"e0",
          1182 => x"82",
          1183 => x"82",
          1184 => x"e0",
          1185 => x"e0",
          1186 => x"82",
          1187 => x"e0",
          1188 => x"a4",
          1189 => x"82",
          1190 => x"e0",
          1191 => x"a4",
          1192 => x"08",
          1193 => x"51",
          1194 => x"a4",
          1195 => x"0b",
          1196 => x"82",
          1197 => x"e0",
          1198 => x"82",
          1199 => x"82",
          1200 => x"2a",
          1201 => x"82",
          1202 => x"e0",
          1203 => x"a4",
          1204 => x"06",
          1205 => x"82",
          1206 => x"39",
          1207 => x"05",
          1208 => x"08",
          1209 => x"88",
          1210 => x"08",
          1211 => x"08",
          1212 => x"05",
          1213 => x"08",
          1214 => x"05",
          1215 => x"82",
          1216 => x"f0",
          1217 => x"0b",
          1218 => x"8a",
          1219 => x"e8",
          1220 => x"05",
          1221 => x"0c",
          1222 => x"05",
          1223 => x"05",
          1224 => x"fc",
          1225 => x"05",
          1226 => x"08",
          1227 => x"0c",
          1228 => x"8c",
          1229 => x"0b",
          1230 => x"8a",
          1231 => x"e4",
          1232 => x"05",
          1233 => x"0c",
          1234 => x"05",
          1235 => x"05",
          1236 => x"fc",
          1237 => x"05",
          1238 => x"08",
          1239 => x"0c",
          1240 => x"05",
          1241 => x"05",
          1242 => x"81",
          1243 => x"e0",
          1244 => x"70",
          1245 => x"51",
          1246 => x"0d",
          1247 => x"a4",
          1248 => x"3d",
          1249 => x"08",
          1250 => x"08",
          1251 => x"08",
          1252 => x"08",
          1253 => x"08",
          1254 => x"51",
          1255 => x"a4",
          1256 => x"82",
          1257 => x"e0",
          1258 => x"e0",
          1259 => x"3f",
          1260 => x"98",
          1261 => x"a4",
          1262 => x"82",
          1263 => x"0b",
          1264 => x"82",
          1265 => x"2e",
          1266 => x"05",
          1267 => x"98",
          1268 => x"05",
          1269 => x"08",
          1270 => x"e4",
          1271 => x"05",
          1272 => x"a4",
          1273 => x"3f",
          1274 => x"08",
          1275 => x"a4",
          1276 => x"82",
          1277 => x"e0",
          1278 => x"e0",
          1279 => x"a4",
          1280 => x"08",
          1281 => x"fc",
          1282 => x"e0",
          1283 => x"38",
          1284 => x"70",
          1285 => x"52",
          1286 => x"fc",
          1287 => x"e0",
          1288 => x"81",
          1289 => x"a4",
          1290 => x"82",
          1291 => x"05",
          1292 => x"82",
          1293 => x"e0",
          1294 => x"e0",
          1295 => x"a4",
          1296 => x"08",
          1297 => x"08",
          1298 => x"a4",
          1299 => x"82",
          1300 => x"e0",
          1301 => x"81",
          1302 => x"05",
          1303 => x"05",
          1304 => x"88",
          1305 => x"82",
          1306 => x"e0",
          1307 => x"82",
          1308 => x"82",
          1309 => x"e0",
          1310 => x"a4",
          1311 => x"82",
          1312 => x"05",
          1313 => x"ec",
          1314 => x"05",
          1315 => x"f0",
          1316 => x"05",
          1317 => x"08",
          1318 => x"08",
          1319 => x"05",
          1320 => x"08",
          1321 => x"05",
          1322 => x"53",
          1323 => x"08",
          1324 => x"08",
          1325 => x"08",
          1326 => x"8c",
          1327 => x"82",
          1328 => x"0c",
          1329 => x"a4",
          1330 => x"08",
          1331 => x"fc",
          1332 => x"f8",
          1333 => x"05",
          1334 => x"08",
          1335 => x"0c",
          1336 => x"82",
          1337 => x"70",
          1338 => x"31",
          1339 => x"82",
          1340 => x"e0",
          1341 => x"82",
          1342 => x"82",
          1343 => x"e0",
          1344 => x"a4",
          1345 => x"a4",
          1346 => x"08",
          1347 => x"08",
          1348 => x"ac",
          1349 => x"e0",
          1350 => x"82",
          1351 => x"70",
          1352 => x"87",
          1353 => x"82",
          1354 => x"0c",
          1355 => x"a4",
          1356 => x"08",
          1357 => x"82",
          1358 => x"08",
          1359 => x"e0",
          1360 => x"ff",
          1361 => x"06",
          1362 => x"05",
          1363 => x"53",
          1364 => x"05",
          1365 => x"06",
          1366 => x"08",
          1367 => x"88",
          1368 => x"0c",
          1369 => x"e0",
          1370 => x"a4",
          1371 => x"2e",
          1372 => x"e0",
          1373 => x"81",
          1374 => x"72",
          1375 => x"34",
          1376 => x"82",
          1377 => x"e0",
          1378 => x"2e",
          1379 => x"05",
          1380 => x"cd",
          1381 => x"f4",
          1382 => x"05",
          1383 => x"70",
          1384 => x"a4",
          1385 => x"82",
          1386 => x"34",
          1387 => x"70",
          1388 => x"51",
          1389 => x"f8",
          1390 => x"a4",
          1391 => x"26",
          1392 => x"08",
          1393 => x"e0",
          1394 => x"73",
          1395 => x"f8",
          1396 => x"38",
          1397 => x"08",
          1398 => x"0b",
          1399 => x"b2",
          1400 => x"33",
          1401 => x"e0",
          1402 => x"b9",
          1403 => x"82",
          1404 => x"a5",
          1405 => x"f4",
          1406 => x"08",
          1407 => x"f8",
          1408 => x"cf",
          1409 => x"33",
          1410 => x"82",
          1411 => x"11",
          1412 => x"f8",
          1413 => x"05",
          1414 => x"e0",
          1415 => x"a4",
          1416 => x"27",
          1417 => x"05",
          1418 => x"e0",
          1419 => x"a4",
          1420 => x"26",
          1421 => x"08",
          1422 => x"e0",
          1423 => x"a4",
          1424 => x"74",
          1425 => x"a4",
          1426 => x"82",
          1427 => x"82",
          1428 => x"82",
          1429 => x"12",
          1430 => x"82",
          1431 => x"08",
          1432 => x"51",
          1433 => x"a4",
          1434 => x"82",
          1435 => x"72",
          1436 => x"08",
          1437 => x"08",
          1438 => x"8c",
          1439 => x"05",
          1440 => x"e0",
          1441 => x"a4",
          1442 => x"0c",
          1443 => x"04",
          1444 => x"a4",
          1445 => x"e0",
          1446 => x"a4",
          1447 => x"0c",
          1448 => x"70",
          1449 => x"82",
          1450 => x"81",
          1451 => x"81",
          1452 => x"88",
          1453 => x"0c",
          1454 => x"f8",
          1455 => x"81",
          1456 => x"a4",
          1457 => x"08",
          1458 => x"71",
          1459 => x"82",
          1460 => x"e0",
          1461 => x"b0",
          1462 => x"82",
          1463 => x"08",
          1464 => x"53",
          1465 => x"05",
          1466 => x"33",
          1467 => x"82",
          1468 => x"e2",
          1469 => x"e8",
          1470 => x"80",
          1471 => x"08",
          1472 => x"88",
          1473 => x"0c",
          1474 => x"e0",
          1475 => x"39",
          1476 => x"05",
          1477 => x"08",
          1478 => x"08",
          1479 => x"08",
          1480 => x"e0",
          1481 => x"a0",
          1482 => x"a4",
          1483 => x"82",
          1484 => x"af",
          1485 => x"08",
          1486 => x"83",
          1487 => x"a4",
          1488 => x"88",
          1489 => x"34",
          1490 => x"05",
          1491 => x"82",
          1492 => x"72",
          1493 => x"0b",
          1494 => x"82",
          1495 => x"08",
          1496 => x"a4",
          1497 => x"08",
          1498 => x"81",
          1499 => x"05",
          1500 => x"38",
          1501 => x"e0",
          1502 => x"08",
          1503 => x"f8",
          1504 => x"82",
          1505 => x"e0",
          1506 => x"73",
          1507 => x"f8",
          1508 => x"82",
          1509 => x"e0",
          1510 => x"89",
          1511 => x"a4",
          1512 => x"82",
          1513 => x"e0",
          1514 => x"72",
          1515 => x"e0",
          1516 => x"39",
          1517 => x"70",
          1518 => x"29",
          1519 => x"70",
          1520 => x"0c",
          1521 => x"70",
          1522 => x"51",
          1523 => x"e0",
          1524 => x"39",
          1525 => x"53",
          1526 => x"a4",
          1527 => x"a4",
          1528 => x"08",
          1529 => x"fc",
          1530 => x"82",
          1531 => x"e0",
          1532 => x"98",
          1533 => x"0c",
          1534 => x"70",
          1535 => x"df",
          1536 => x"85",
          1537 => x"33",
          1538 => x"86",
          1539 => x"57",
          1540 => x"70",
          1541 => x"e0",
          1542 => x"75",
          1543 => x"3f",
          1544 => x"16",
          1545 => x"38",
          1546 => x"54",
          1547 => x"73",
          1548 => x"04",
          1549 => x"04",
          1550 => x"26",
          1551 => x"b7",
          1552 => x"bd",
          1553 => x"f0",
          1554 => x"51",
          1555 => x"80",
          1556 => x"e4",
          1557 => x"39",
          1558 => x"82",
          1559 => x"be",
          1560 => x"84",
          1561 => x"51",
          1562 => x"39",
          1563 => x"bf",
          1564 => x"51",
          1565 => x"39",
          1566 => x"c0",
          1567 => x"51",
          1568 => x"39",
          1569 => x"83",
          1570 => x"79",
          1571 => x"38",
          1572 => x"90",
          1573 => x"a4",
          1574 => x"51",
          1575 => x"54",
          1576 => x"51",
          1577 => x"04",
          1578 => x"80",
          1579 => x"78",
          1580 => x"57",
          1581 => x"26",
          1582 => x"70",
          1583 => x"74",
          1584 => x"8c",
          1585 => x"3f",
          1586 => x"98",
          1587 => x"87",
          1588 => x"08",
          1589 => x"80",
          1590 => x"d5",
          1591 => x"e0",
          1592 => x"80",
          1593 => x"59",
          1594 => x"51",
          1595 => x"78",
          1596 => x"2a",
          1597 => x"80",
          1598 => x"87",
          1599 => x"fe",
          1600 => x"98",
          1601 => x"0d",
          1602 => x"58",
          1603 => x"7a",
          1604 => x"08",
          1605 => x"76",
          1606 => x"fb",
          1607 => x"e0",
          1608 => x"2d",
          1609 => x"78",
          1610 => x"3d",
          1611 => x"63",
          1612 => x"73",
          1613 => x"5e",
          1614 => x"3f",
          1615 => x"53",
          1616 => x"90",
          1617 => x"86",
          1618 => x"58",
          1619 => x"ae",
          1620 => x"ae",
          1621 => x"81",
          1622 => x"7b",
          1623 => x"74",
          1624 => x"72",
          1625 => x"ae",
          1626 => x"51",
          1627 => x"80",
          1628 => x"27",
          1629 => x"c4",
          1630 => x"82",
          1631 => x"84",
          1632 => x"72",
          1633 => x"82",
          1634 => x"89",
          1635 => x"ed",
          1636 => x"08",
          1637 => x"fc",
          1638 => x"d5",
          1639 => x"c6",
          1640 => x"80",
          1641 => x"56",
          1642 => x"81",
          1643 => x"06",
          1644 => x"73",
          1645 => x"fc",
          1646 => x"fb",
          1647 => x"3f",
          1648 => x"c1",
          1649 => x"78",
          1650 => x"3f",
          1651 => x"98",
          1652 => x"81",
          1653 => x"3f",
          1654 => x"98",
          1655 => x"9b",
          1656 => x"75",
          1657 => x"51",
          1658 => x"9b",
          1659 => x"72",
          1660 => x"72",
          1661 => x"04",
          1662 => x"55",
          1663 => x"f8",
          1664 => x"85",
          1665 => x"d8",
          1666 => x"90",
          1667 => x"c2",
          1668 => x"80",
          1669 => x"3d",
          1670 => x"96",
          1671 => x"51",
          1672 => x"9a",
          1673 => x"72",
          1674 => x"71",
          1675 => x"a1",
          1676 => x"3f",
          1677 => x"2a",
          1678 => x"2e",
          1679 => x"82",
          1680 => x"51",
          1681 => x"81",
          1682 => x"38",
          1683 => x"ec",
          1684 => x"d9",
          1685 => x"51",
          1686 => x"51",
          1687 => x"99",
          1688 => x"72",
          1689 => x"71",
          1690 => x"a9",
          1691 => x"3f",
          1692 => x"2a",
          1693 => x"2e",
          1694 => x"82",
          1695 => x"51",
          1696 => x"81",
          1697 => x"38",
          1698 => x"bc",
          1699 => x"e1",
          1700 => x"51",
          1701 => x"51",
          1702 => x"98",
          1703 => x"a4",
          1704 => x"3d",
          1705 => x"33",
          1706 => x"51",
          1707 => x"9c",
          1708 => x"82",
          1709 => x"81",
          1710 => x"30",
          1711 => x"25",
          1712 => x"0b",
          1713 => x"82",
          1714 => x"09",
          1715 => x"53",
          1716 => x"3f",
          1717 => x"38",
          1718 => x"3f",
          1719 => x"97",
          1720 => x"db",
          1721 => x"33",
          1722 => x"8c",
          1723 => x"75",
          1724 => x"e0",
          1725 => x"3d",
          1726 => x"82",
          1727 => x"51",
          1728 => x"08",
          1729 => x"09",
          1730 => x"83",
          1731 => x"d1",
          1732 => x"e1",
          1733 => x"e0",
          1734 => x"c4",
          1735 => x"41",
          1736 => x"c5",
          1737 => x"f8",
          1738 => x"3d",
          1739 => x"82",
          1740 => x"2c",
          1741 => x"a5",
          1742 => x"78",
          1743 => x"24",
          1744 => x"38",
          1745 => x"dc",
          1746 => x"38",
          1747 => x"78",
          1748 => x"39",
          1749 => x"78",
          1750 => x"c3",
          1751 => x"2e",
          1752 => x"81",
          1753 => x"83",
          1754 => x"89",
          1755 => x"85",
          1756 => x"b5",
          1757 => x"05",
          1758 => x"08",
          1759 => x"fe",
          1760 => x"ec",
          1761 => x"2e",
          1762 => x"11",
          1763 => x"3f",
          1764 => x"e0",
          1765 => x"ff",
          1766 => x"79",
          1767 => x"78",
          1768 => x"7a",
          1769 => x"3d",
          1770 => x"51",
          1771 => x"80",
          1772 => x"fc",
          1773 => x"b0",
          1774 => x"fd",
          1775 => x"53",
          1776 => x"82",
          1777 => x"38",
          1778 => x"3f",
          1779 => x"38",
          1780 => x"33",
          1781 => x"39",
          1782 => x"84",
          1783 => x"98",
          1784 => x"3d",
          1785 => x"51",
          1786 => x"80",
          1787 => x"f8",
          1788 => x"b8",
          1789 => x"fc",
          1790 => x"a4",
          1791 => x"a8",
          1792 => x"5a",
          1793 => x"55",
          1794 => x"82",
          1795 => x"81",
          1796 => x"39",
          1797 => x"39",
          1798 => x"84",
          1799 => x"98",
          1800 => x"33",
          1801 => x"de",
          1802 => x"de",
          1803 => x"38",
          1804 => x"82",
          1805 => x"88",
          1806 => x"39",
          1807 => x"2e",
          1808 => x"9a",
          1809 => x"80",
          1810 => x"45",
          1811 => x"80",
          1812 => x"53",
          1813 => x"82",
          1814 => x"de",
          1815 => x"38",
          1816 => x"39",
          1817 => x"2e",
          1818 => x"bb",
          1819 => x"80",
          1820 => x"44",
          1821 => x"78",
          1822 => x"08",
          1823 => x"59",
          1824 => x"d8",
          1825 => x"08",
          1826 => x"11",
          1827 => x"3f",
          1828 => x"38",
          1829 => x"83",
          1830 => x"30",
          1831 => x"06",
          1832 => x"88",
          1833 => x"43",
          1834 => x"3f",
          1835 => x"52",
          1836 => x"bc",
          1837 => x"80",
          1838 => x"a8",
          1839 => x"f9",
          1840 => x"53",
          1841 => x"82",
          1842 => x"64",
          1843 => x"34",
          1844 => x"fc",
          1845 => x"f0",
          1846 => x"f9",
          1847 => x"82",
          1848 => x"82",
          1849 => x"79",
          1850 => x"79",
          1851 => x"38",
          1852 => x"fe",
          1853 => x"e6",
          1854 => x"2e",
          1855 => x"05",
          1856 => x"ff",
          1857 => x"bc",
          1858 => x"fe",
          1859 => x"e0",
          1860 => x"2e",
          1861 => x"11",
          1862 => x"3f",
          1863 => x"38",
          1864 => x"79",
          1865 => x"b5",
          1866 => x"05",
          1867 => x"08",
          1868 => x"22",
          1869 => x"9f",
          1870 => x"80",
          1871 => x"3f",
          1872 => x"2e",
          1873 => x"38",
          1874 => x"3d",
          1875 => x"51",
          1876 => x"80",
          1877 => x"c2",
          1878 => x"23",
          1879 => x"d4",
          1880 => x"39",
          1881 => x"84",
          1882 => x"98",
          1883 => x"3d",
          1884 => x"51",
          1885 => x"80",
          1886 => x"59",
          1887 => x"f0",
          1888 => x"c7",
          1889 => x"f6",
          1890 => x"82",
          1891 => x"82",
          1892 => x"79",
          1893 => x"79",
          1894 => x"38",
          1895 => x"fe",
          1896 => x"de",
          1897 => x"2e",
          1898 => x"61",
          1899 => x"c5",
          1900 => x"aa",
          1901 => x"ff",
          1902 => x"e0",
          1903 => x"64",
          1904 => x"85",
          1905 => x"ff",
          1906 => x"e3",
          1907 => x"2e",
          1908 => x"90",
          1909 => x"78",
          1910 => x"f5",
          1911 => x"82",
          1912 => x"f4",
          1913 => x"b8",
          1914 => x"e9",
          1915 => x"b8",
          1916 => x"ce",
          1917 => x"59",
          1918 => x"f8",
          1919 => x"e0",
          1920 => x"80",
          1921 => x"08",
          1922 => x"83",
          1923 => x"7f",
          1924 => x"d2",
          1925 => x"8a",
          1926 => x"81",
          1927 => x"b2",
          1928 => x"81",
          1929 => x"83",
          1930 => x"c6",
          1931 => x"54",
          1932 => x"3d",
          1933 => x"3f",
          1934 => x"b0",
          1935 => x"7b",
          1936 => x"82",
          1937 => x"05",
          1938 => x"7b",
          1939 => x"b5",
          1940 => x"cd",
          1941 => x"c8",
          1942 => x"90",
          1943 => x"b5",
          1944 => x"3f",
          1945 => x"08",
          1946 => x"25",
          1947 => x"83",
          1948 => x"06",
          1949 => x"1b",
          1950 => x"fe",
          1951 => x"32",
          1952 => x"2e",
          1953 => x"a4",
          1954 => x"b1",
          1955 => x"b4",
          1956 => x"39",
          1957 => x"c8",
          1958 => x"54",
          1959 => x"cb",
          1960 => x"2b",
          1961 => x"52",
          1962 => x"e0",
          1963 => x"94",
          1964 => x"80",
          1965 => x"e0",
          1966 => x"53",
          1967 => x"d4",
          1968 => x"75",
          1969 => x"94",
          1970 => x"c0",
          1971 => x"81",
          1972 => x"99",
          1973 => x"0b",
          1974 => x"72",
          1975 => x"aa",
          1976 => x"51",
          1977 => x"51",
          1978 => x"51",
          1979 => x"3f",
          1980 => x"0d",
          1981 => x"52",
          1982 => x"72",
          1983 => x"06",
          1984 => x"72",
          1985 => x"06",
          1986 => x"72",
          1987 => x"9f",
          1988 => x"72",
          1989 => x"38",
          1990 => x"73",
          1991 => x"80",
          1992 => x"83",
          1993 => x"38",
          1994 => x"54",
          1995 => x"38",
          1996 => x"70",
          1997 => x"70",
          1998 => x"81",
          1999 => x"51",
          2000 => x"0d",
          2001 => x"08",
          2002 => x"05",
          2003 => x"e0",
          2004 => x"39",
          2005 => x"86",
          2006 => x"82",
          2007 => x"52",
          2008 => x"13",
          2009 => x"9e",
          2010 => x"51",
          2011 => x"38",
          2012 => x"bb",
          2013 => x"51",
          2014 => x"38",
          2015 => x"87",
          2016 => x"22",
          2017 => x"80",
          2018 => x"9c",
          2019 => x"0c",
          2020 => x"0c",
          2021 => x"0c",
          2022 => x"0c",
          2023 => x"0c",
          2024 => x"0c",
          2025 => x"87",
          2026 => x"c0",
          2027 => x"e0",
          2028 => x"3d",
          2029 => x"5d",
          2030 => x"08",
          2031 => x"b8",
          2032 => x"c0",
          2033 => x"34",
          2034 => x"84",
          2035 => x"5a",
          2036 => x"a8",
          2037 => x"c0",
          2038 => x"23",
          2039 => x"8a",
          2040 => x"ff",
          2041 => x"06",
          2042 => x"33",
          2043 => x"33",
          2044 => x"ff",
          2045 => x"ff",
          2046 => x"fd",
          2047 => x"80",
          2048 => x"83",
          2049 => x"30",
          2050 => x"51",
          2051 => x"3f",
          2052 => x"98",
          2053 => x"52",
          2054 => x"38",
          2055 => x"06",
          2056 => x"70",
          2057 => x"51",
          2058 => x"e0",
          2059 => x"3d",
          2060 => x"2b",
          2061 => x"e0",
          2062 => x"74",
          2063 => x"80",
          2064 => x"0c",
          2065 => x"02",
          2066 => x"70",
          2067 => x"c0",
          2068 => x"38",
          2069 => x"70",
          2070 => x"52",
          2071 => x"2a",
          2072 => x"38",
          2073 => x"51",
          2074 => x"2a",
          2075 => x"be",
          2076 => x"c0",
          2077 => x"38",
          2078 => x"0c",
          2079 => x"0d",
          2080 => x"33",
          2081 => x"52",
          2082 => x"0d",
          2083 => x"33",
          2084 => x"87",
          2085 => x"82",
          2086 => x"58",
          2087 => x"80",
          2088 => x"53",
          2089 => x"06",
          2090 => x"38",
          2091 => x"53",
          2092 => x"81",
          2093 => x"38",
          2094 => x"53",
          2095 => x"06",
          2096 => x"80",
          2097 => x"54",
          2098 => x"98",
          2099 => x"0d",
          2100 => x"ff",
          2101 => x"80",
          2102 => x"15",
          2103 => x"06",
          2104 => x"84",
          2105 => x"c0",
          2106 => x"2a",
          2107 => x"80",
          2108 => x"81",
          2109 => x"81",
          2110 => x"80",
          2111 => x"81",
          2112 => x"74",
          2113 => x"80",
          2114 => x"c0",
          2115 => x"17",
          2116 => x"53",
          2117 => x"e0",
          2118 => x"3d",
          2119 => x"ff",
          2120 => x"51",
          2121 => x"94",
          2122 => x"70",
          2123 => x"2e",
          2124 => x"87",
          2125 => x"86",
          2126 => x"08",
          2127 => x"0c",
          2128 => x"3f",
          2129 => x"82",
          2130 => x"82",
          2131 => x"52",
          2132 => x"80",
          2133 => x"52",
          2134 => x"06",
          2135 => x"2e",
          2136 => x"87",
          2137 => x"86",
          2138 => x"08",
          2139 => x"53",
          2140 => x"3d",
          2141 => x"9e",
          2142 => x"51",
          2143 => x"87",
          2144 => x"0c",
          2145 => x"b8",
          2146 => x"de",
          2147 => x"82",
          2148 => x"08",
          2149 => x"a0",
          2150 => x"9e",
          2151 => x"c0",
          2152 => x"87",
          2153 => x"0c",
          2154 => x"d8",
          2155 => x"de",
          2156 => x"82",
          2157 => x"08",
          2158 => x"80",
          2159 => x"87",
          2160 => x"0c",
          2161 => x"f0",
          2162 => x"de",
          2163 => x"34",
          2164 => x"70",
          2165 => x"70",
          2166 => x"82",
          2167 => x"9e",
          2168 => x"51",
          2169 => x"81",
          2170 => x"0b",
          2171 => x"80",
          2172 => x"2e",
          2173 => x"fb",
          2174 => x"08",
          2175 => x"52",
          2176 => x"71",
          2177 => x"c0",
          2178 => x"06",
          2179 => x"38",
          2180 => x"80",
          2181 => x"90",
          2182 => x"80",
          2183 => x"de",
          2184 => x"90",
          2185 => x"52",
          2186 => x"52",
          2187 => x"87",
          2188 => x"80",
          2189 => x"83",
          2190 => x"34",
          2191 => x"70",
          2192 => x"70",
          2193 => x"82",
          2194 => x"9e",
          2195 => x"51",
          2196 => x"81",
          2197 => x"0b",
          2198 => x"80",
          2199 => x"83",
          2200 => x"34",
          2201 => x"80",
          2202 => x"70",
          2203 => x"c0",
          2204 => x"51",
          2205 => x"81",
          2206 => x"c0",
          2207 => x"70",
          2208 => x"df",
          2209 => x"90",
          2210 => x"70",
          2211 => x"82",
          2212 => x"08",
          2213 => x"df",
          2214 => x"3d",
          2215 => x"cd",
          2216 => x"80",
          2217 => x"ff",
          2218 => x"ff",
          2219 => x"54",
          2220 => x"d4",
          2221 => x"52",
          2222 => x"3f",
          2223 => x"2e",
          2224 => x"de",
          2225 => x"f8",
          2226 => x"fc",
          2227 => x"82",
          2228 => x"11",
          2229 => x"88",
          2230 => x"73",
          2231 => x"08",
          2232 => x"82",
          2233 => x"82",
          2234 => x"94",
          2235 => x"c8",
          2236 => x"51",
          2237 => x"33",
          2238 => x"df",
          2239 => x"ff",
          2240 => x"54",
          2241 => x"88",
          2242 => x"87",
          2243 => x"73",
          2244 => x"33",
          2245 => x"dd",
          2246 => x"80",
          2247 => x"ff",
          2248 => x"54",
          2249 => x"dc",
          2250 => x"80",
          2251 => x"82",
          2252 => x"82",
          2253 => x"89",
          2254 => x"a0",
          2255 => x"80",
          2256 => x"ff",
          2257 => x"ff",
          2258 => x"52",
          2259 => x"3f",
          2260 => x"b8",
          2261 => x"e4",
          2262 => x"86",
          2263 => x"a2",
          2264 => x"82",
          2265 => x"82",
          2266 => x"52",
          2267 => x"e0",
          2268 => x"71",
          2269 => x"52",
          2270 => x"3f",
          2271 => x"2e",
          2272 => x"bd",
          2273 => x"c4",
          2274 => x"c0",
          2275 => x"e0",
          2276 => x"ff",
          2277 => x"54",
          2278 => x"f4",
          2279 => x"51",
          2280 => x"08",
          2281 => x"54",
          2282 => x"cd",
          2283 => x"51",
          2284 => x"04",
          2285 => x"ff",
          2286 => x"71",
          2287 => x"71",
          2288 => x"39",
          2289 => x"cd",
          2290 => x"51",
          2291 => x"39",
          2292 => x"3f",
          2293 => x"0c",
          2294 => x"0c",
          2295 => x"96",
          2296 => x"98",
          2297 => x"70",
          2298 => x"2b",
          2299 => x"0b",
          2300 => x"71",
          2301 => x"11",
          2302 => x"33",
          2303 => x"2e",
          2304 => x"72",
          2305 => x"04",
          2306 => x"a3",
          2307 => x"72",
          2308 => x"08",
          2309 => x"82",
          2310 => x"a3",
          2311 => x"88",
          2312 => x"ff",
          2313 => x"ff",
          2314 => x"83",
          2315 => x"0d",
          2316 => x"05",
          2317 => x"05",
          2318 => x"29",
          2319 => x"59",
          2320 => x"86",
          2321 => x"df",
          2322 => x"90",
          2323 => x"5a",
          2324 => x"75",
          2325 => x"29",
          2326 => x"56",
          2327 => x"53",
          2328 => x"3f",
          2329 => x"74",
          2330 => x"06",
          2331 => x"0b",
          2332 => x"b6",
          2333 => x"80",
          2334 => x"55",
          2335 => x"54",
          2336 => x"ec",
          2337 => x"8a",
          2338 => x"e4",
          2339 => x"3d",
          2340 => x"90",
          2341 => x"80",
          2342 => x"3f",
          2343 => x"54",
          2344 => x"0b",
          2345 => x"08",
          2346 => x"51",
          2347 => x"08",
          2348 => x"df",
          2349 => x"3d",
          2350 => x"e4",
          2351 => x"e0",
          2352 => x"e4",
          2353 => x"70",
          2354 => x"e0",
          2355 => x"51",
          2356 => x"08",
          2357 => x"25",
          2358 => x"05",
          2359 => x"75",
          2360 => x"dc",
          2361 => x"ff",
          2362 => x"a6",
          2363 => x"3d",
          2364 => x"70",
          2365 => x"08",
          2366 => x"98",
          2367 => x"df",
          2368 => x"8b",
          2369 => x"3f",
          2370 => x"38",
          2371 => x"e0",
          2372 => x"0b",
          2373 => x"82",
          2374 => x"55",
          2375 => x"30",
          2376 => x"55",
          2377 => x"ac",
          2378 => x"08",
          2379 => x"e0",
          2380 => x"d0",
          2381 => x"77",
          2382 => x"52",
          2383 => x"51",
          2384 => x"54",
          2385 => x"58",
          2386 => x"0d",
          2387 => x"5c",
          2388 => x"73",
          2389 => x"78",
          2390 => x"98",
          2391 => x"33",
          2392 => x"81",
          2393 => x"38",
          2394 => x"ec",
          2395 => x"da",
          2396 => x"52",
          2397 => x"82",
          2398 => x"15",
          2399 => x"74",
          2400 => x"e6",
          2401 => x"3d",
          2402 => x"88",
          2403 => x"9a",
          2404 => x"51",
          2405 => x"81",
          2406 => x"54",
          2407 => x"06",
          2408 => x"38",
          2409 => x"8c",
          2410 => x"3d",
          2411 => x"59",
          2412 => x"82",
          2413 => x"55",
          2414 => x"df",
          2415 => x"81",
          2416 => x"81",
          2417 => x"2e",
          2418 => x"3f",
          2419 => x"0c",
          2420 => x"92",
          2421 => x"98",
          2422 => x"e0",
          2423 => x"d1",
          2424 => x"f7",
          2425 => x"df",
          2426 => x"3d",
          2427 => x"82",
          2428 => x"08",
          2429 => x"38",
          2430 => x"c2",
          2431 => x"0b",
          2432 => x"82",
          2433 => x"55",
          2434 => x"81",
          2435 => x"3f",
          2436 => x"54",
          2437 => x"74",
          2438 => x"38",
          2439 => x"76",
          2440 => x"2e",
          2441 => x"5d",
          2442 => x"98",
          2443 => x"59",
          2444 => x"ff",
          2445 => x"2b",
          2446 => x"70",
          2447 => x"2c",
          2448 => x"05",
          2449 => x"51",
          2450 => x"81",
          2451 => x"77",
          2452 => x"0a",
          2453 => x"2c",
          2454 => x"38",
          2455 => x"83",
          2456 => x"06",
          2457 => x"82",
          2458 => x"74",
          2459 => x"05",
          2460 => x"56",
          2461 => x"76",
          2462 => x"3f",
          2463 => x"54",
          2464 => x"75",
          2465 => x"55",
          2466 => x"2b",
          2467 => x"70",
          2468 => x"11",
          2469 => x"33",
          2470 => x"55",
          2471 => x"90",
          2472 => x"0c",
          2473 => x"0b",
          2474 => x"82",
          2475 => x"34",
          2476 => x"7e",
          2477 => x"73",
          2478 => x"73",
          2479 => x"73",
          2480 => x"d8",
          2481 => x"74",
          2482 => x"73",
          2483 => x"73",
          2484 => x"0a",
          2485 => x"2c",
          2486 => x"df",
          2487 => x"56",
          2488 => x"1a",
          2489 => x"f7",
          2490 => x"38",
          2491 => x"34",
          2492 => x"0a",
          2493 => x"2c",
          2494 => x"56",
          2495 => x"fc",
          2496 => x"54",
          2497 => x"0a",
          2498 => x"2c",
          2499 => x"73",
          2500 => x"33",
          2501 => x"f7",
          2502 => x"77",
          2503 => x"08",
          2504 => x"74",
          2505 => x"05",
          2506 => x"56",
          2507 => x"fb",
          2508 => x"81",
          2509 => x"52",
          2510 => x"81",
          2511 => x"81",
          2512 => x"fb",
          2513 => x"05",
          2514 => x"15",
          2515 => x"fb",
          2516 => x"bf",
          2517 => x"2b",
          2518 => x"57",
          2519 => x"38",
          2520 => x"34",
          2521 => x"51",
          2522 => x"0a",
          2523 => x"2c",
          2524 => x"75",
          2525 => x"08",
          2526 => x"82",
          2527 => x"98",
          2528 => x"56",
          2529 => x"82",
          2530 => x"95",
          2531 => x"81",
          2532 => x"f7",
          2533 => x"25",
          2534 => x"d8",
          2535 => x"82",
          2536 => x"95",
          2537 => x"51",
          2538 => x"81",
          2539 => x"f7",
          2540 => x"38",
          2541 => x"f1",
          2542 => x"0b",
          2543 => x"f7",
          2544 => x"af",
          2545 => x"54",
          2546 => x"fb",
          2547 => x"c7",
          2548 => x"54",
          2549 => x"ff",
          2550 => x"33",
          2551 => x"75",
          2552 => x"73",
          2553 => x"70",
          2554 => x"51",
          2555 => x"1a",
          2556 => x"fb",
          2557 => x"93",
          2558 => x"81",
          2559 => x"f7",
          2560 => x"24",
          2561 => x"a0",
          2562 => x"dc",
          2563 => x"82",
          2564 => x"74",
          2565 => x"fc",
          2566 => x"3f",
          2567 => x"0a",
          2568 => x"33",
          2569 => x"38",
          2570 => x"70",
          2571 => x"59",
          2572 => x"38",
          2573 => x"54",
          2574 => x"70",
          2575 => x"82",
          2576 => x"82",
          2577 => x"75",
          2578 => x"f7",
          2579 => x"51",
          2580 => x"dc",
          2581 => x"f7",
          2582 => x"dc",
          2583 => x"74",
          2584 => x"98",
          2585 => x"98",
          2586 => x"74",
          2587 => x"93",
          2588 => x"82",
          2589 => x"54",
          2590 => x"ff",
          2591 => x"82",
          2592 => x"81",
          2593 => x"79",
          2594 => x"54",
          2595 => x"80",
          2596 => x"9a",
          2597 => x"09",
          2598 => x"08",
          2599 => x"51",
          2600 => x"08",
          2601 => x"08",
          2602 => x"52",
          2603 => x"c3",
          2604 => x"05",
          2605 => x"ab",
          2606 => x"82",
          2607 => x"82",
          2608 => x"05",
          2609 => x"8a",
          2610 => x"06",
          2611 => x"34",
          2612 => x"82",
          2613 => x"e0",
          2614 => x"33",
          2615 => x"33",
          2616 => x"85",
          2617 => x"14",
          2618 => x"1a",
          2619 => x"3f",
          2620 => x"54",
          2621 => x"fb",
          2622 => x"ef",
          2623 => x"54",
          2624 => x"39",
          2625 => x"82",
          2626 => x"e0",
          2627 => x"52",
          2628 => x"3f",
          2629 => x"77",
          2630 => x"34",
          2631 => x"15",
          2632 => x"88",
          2633 => x"87",
          2634 => x"e0",
          2635 => x"07",
          2636 => x"2a",
          2637 => x"34",
          2638 => x"22",
          2639 => x"05",
          2640 => x"15",
          2641 => x"0d",
          2642 => x"51",
          2643 => x"83",
          2644 => x"06",
          2645 => x"0c",
          2646 => x"02",
          2647 => x"05",
          2648 => x"71",
          2649 => x"73",
          2650 => x"88",
          2651 => x"22",
          2652 => x"88",
          2653 => x"5b",
          2654 => x"70",
          2655 => x"14",
          2656 => x"15",
          2657 => x"88",
          2658 => x"33",
          2659 => x"8f",
          2660 => x"71",
          2661 => x"88",
          2662 => x"34",
          2663 => x"12",
          2664 => x"71",
          2665 => x"3d",
          2666 => x"88",
          2667 => x"70",
          2668 => x"87",
          2669 => x"2b",
          2670 => x"72",
          2671 => x"71",
          2672 => x"56",
          2673 => x"85",
          2674 => x"14",
          2675 => x"8b",
          2676 => x"57",
          2677 => x"13",
          2678 => x"2a",
          2679 => x"34",
          2680 => x"08",
          2681 => x"88",
          2682 => x"70",
          2683 => x"71",
          2684 => x"3d",
          2685 => x"05",
          2686 => x"2b",
          2687 => x"71",
          2688 => x"70",
          2689 => x"71",
          2690 => x"52",
          2691 => x"25",
          2692 => x"3f",
          2693 => x"33",
          2694 => x"83",
          2695 => x"12",
          2696 => x"2b",
          2697 => x"51",
          2698 => x"88",
          2699 => x"73",
          2700 => x"70",
          2701 => x"8b",
          2702 => x"57",
          2703 => x"33",
          2704 => x"ff",
          2705 => x"58",
          2706 => x"34",
          2707 => x"82",
          2708 => x"05",
          2709 => x"11",
          2710 => x"71",
          2711 => x"56",
          2712 => x"33",
          2713 => x"a2",
          2714 => x"53",
          2715 => x"70",
          2716 => x"70",
          2717 => x"8b",
          2718 => x"57",
          2719 => x"13",
          2720 => x"2a",
          2721 => x"34",
          2722 => x"08",
          2723 => x"71",
          2724 => x"52",
          2725 => x"0d",
          2726 => x"2a",
          2727 => x"57",
          2728 => x"08",
          2729 => x"33",
          2730 => x"83",
          2731 => x"12",
          2732 => x"07",
          2733 => x"55",
          2734 => x"82",
          2735 => x"3f",
          2736 => x"15",
          2737 => x"07",
          2738 => x"55",
          2739 => x"81",
          2740 => x"82",
          2741 => x"33",
          2742 => x"70",
          2743 => x"72",
          2744 => x"82",
          2745 => x"86",
          2746 => x"82",
          2747 => x"34",
          2748 => x"08",
          2749 => x"88",
          2750 => x"70",
          2751 => x"74",
          2752 => x"3d",
          2753 => x"82",
          2754 => x"3f",
          2755 => x"fe",
          2756 => x"3d",
          2757 => x"3f",
          2758 => x"06",
          2759 => x"85",
          2760 => x"5f",
          2761 => x"59",
          2762 => x"88",
          2763 => x"71",
          2764 => x"06",
          2765 => x"70",
          2766 => x"55",
          2767 => x"2e",
          2768 => x"15",
          2769 => x"07",
          2770 => x"ff",
          2771 => x"56",
          2772 => x"08",
          2773 => x"88",
          2774 => x"51",
          2775 => x"2e",
          2776 => x"78",
          2777 => x"80",
          2778 => x"09",
          2779 => x"f2",
          2780 => x"53",
          2781 => x"82",
          2782 => x"33",
          2783 => x"83",
          2784 => x"05",
          2785 => x"70",
          2786 => x"84",
          2787 => x"76",
          2788 => x"75",
          2789 => x"11",
          2790 => x"07",
          2791 => x"5a",
          2792 => x"87",
          2793 => x"1c",
          2794 => x"8b",
          2795 => x"5a",
          2796 => x"34",
          2797 => x"08",
          2798 => x"85",
          2799 => x"88",
          2800 => x"73",
          2801 => x"82",
          2802 => x"73",
          2803 => x"04",
          2804 => x"88",
          2805 => x"53",
          2806 => x"fc",
          2807 => x"72",
          2808 => x"04",
          2809 => x"80",
          2810 => x"60",
          2811 => x"a8",
          2812 => x"b8",
          2813 => x"c7",
          2814 => x"92",
          2815 => x"51",
          2816 => x"83",
          2817 => x"7d",
          2818 => x"ff",
          2819 => x"33",
          2820 => x"70",
          2821 => x"70",
          2822 => x"1a",
          2823 => x"2b",
          2824 => x"53",
          2825 => x"5c",
          2826 => x"38",
          2827 => x"70",
          2828 => x"16",
          2829 => x"07",
          2830 => x"12",
          2831 => x"07",
          2832 => x"80",
          2833 => x"83",
          2834 => x"27",
          2835 => x"7b",
          2836 => x"51",
          2837 => x"06",
          2838 => x"7a",
          2839 => x"aa",
          2840 => x"7a",
          2841 => x"82",
          2842 => x"2b",
          2843 => x"80",
          2844 => x"e0",
          2845 => x"54",
          2846 => x"88",
          2847 => x"ff",
          2848 => x"14",
          2849 => x"59",
          2850 => x"7a",
          2851 => x"f5",
          2852 => x"82",
          2853 => x"2b",
          2854 => x"80",
          2855 => x"e0",
          2856 => x"54",
          2857 => x"88",
          2858 => x"ff",
          2859 => x"14",
          2860 => x"5c",
          2861 => x"39",
          2862 => x"82",
          2863 => x"08",
          2864 => x"52",
          2865 => x"8a",
          2866 => x"58",
          2867 => x"7a",
          2868 => x"19",
          2869 => x"84",
          2870 => x"73",
          2871 => x"04",
          2872 => x"52",
          2873 => x"08",
          2874 => x"8e",
          2875 => x"98",
          2876 => x"82",
          2877 => x"ff",
          2878 => x"81",
          2879 => x"e0",
          2880 => x"98",
          2881 => x"0d",
          2882 => x"9f",
          2883 => x"81",
          2884 => x"87",
          2885 => x"54",
          2886 => x"54",
          2887 => x"11",
          2888 => x"c0",
          2889 => x"70",
          2890 => x"8a",
          2891 => x"70",
          2892 => x"06",
          2893 => x"8c",
          2894 => x"71",
          2895 => x"94",
          2896 => x"0c",
          2897 => x"60",
          2898 => x"33",
          2899 => x"5a",
          2900 => x"81",
          2901 => x"38",
          2902 => x"92",
          2903 => x"87",
          2904 => x"57",
          2905 => x"8c",
          2906 => x"75",
          2907 => x"51",
          2908 => x"7b",
          2909 => x"5d",
          2910 => x"06",
          2911 => x"81",
          2912 => x"72",
          2913 => x"8c",
          2914 => x"98",
          2915 => x"38",
          2916 => x"76",
          2917 => x"72",
          2918 => x"f7",
          2919 => x"80",
          2920 => x"5a",
          2921 => x"73",
          2922 => x"38",
          2923 => x"fc",
          2924 => x"83",
          2925 => x"e0",
          2926 => x"3d",
          2927 => x"bf",
          2928 => x"59",
          2929 => x"82",
          2930 => x"52",
          2931 => x"b1",
          2932 => x"92",
          2933 => x"87",
          2934 => x"56",
          2935 => x"0c",
          2936 => x"58",
          2937 => x"06",
          2938 => x"38",
          2939 => x"0c",
          2940 => x"81",
          2941 => x"38",
          2942 => x"d0",
          2943 => x"71",
          2944 => x"2e",
          2945 => x"92",
          2946 => x"06",
          2947 => x"59",
          2948 => x"06",
          2949 => x"80",
          2950 => x"06",
          2951 => x"fe",
          2952 => x"52",
          2953 => x"71",
          2954 => x"3d",
          2955 => x"84",
          2956 => x"a7",
          2957 => x"fa",
          2958 => x"06",
          2959 => x"85",
          2960 => x"56",
          2961 => x"76",
          2962 => x"c0",
          2963 => x"2e",
          2964 => x"2e",
          2965 => x"08",
          2966 => x"51",
          2967 => x"c0",
          2968 => x"87",
          2969 => x"38",
          2970 => x"14",
          2971 => x"52",
          2972 => x"92",
          2973 => x"39",
          2974 => x"39",
          2975 => x"98",
          2976 => x"0d",
          2977 => x"88",
          2978 => x"51",
          2979 => x"75",
          2980 => x"90",
          2981 => x"33",
          2982 => x"71",
          2983 => x"54",
          2984 => x"ff",
          2985 => x"05",
          2986 => x"05",
          2987 => x"72",
          2988 => x"0d",
          2989 => x"81",
          2990 => x"70",
          2991 => x"88",
          2992 => x"54",
          2993 => x"34",
          2994 => x"76",
          2995 => x"2e",
          2996 => x"33",
          2997 => x"11",
          2998 => x"fe",
          2999 => x"53",
          3000 => x"ff",
          3001 => x"0d",
          3002 => x"56",
          3003 => x"33",
          3004 => x"71",
          3005 => x"72",
          3006 => x"e2",
          3007 => x"3d",
          3008 => x"54",
          3009 => x"38",
          3010 => x"f3",
          3011 => x"84",
          3012 => x"98",
          3013 => x"08",
          3014 => x"54",
          3015 => x"82",
          3016 => x"2e",
          3017 => x"80",
          3018 => x"83",
          3019 => x"86",
          3020 => x"82",
          3021 => x"f7",
          3022 => x"17",
          3023 => x"d6",
          3024 => x"b8",
          3025 => x"59",
          3026 => x"7a",
          3027 => x"e0",
          3028 => x"08",
          3029 => x"08",
          3030 => x"38",
          3031 => x"09",
          3032 => x"18",
          3033 => x"f9",
          3034 => x"82",
          3035 => x"fa",
          3036 => x"57",
          3037 => x"75",
          3038 => x"08",
          3039 => x"81",
          3040 => x"16",
          3041 => x"98",
          3042 => x"81",
          3043 => x"e0",
          3044 => x"3d",
          3045 => x"3f",
          3046 => x"98",
          3047 => x"74",
          3048 => x"38",
          3049 => x"09",
          3050 => x"53",
          3051 => x"70",
          3052 => x"d5",
          3053 => x"3f",
          3054 => x"51",
          3055 => x"f2",
          3056 => x"3f",
          3057 => x"51",
          3058 => x"84",
          3059 => x"17",
          3060 => x"79",
          3061 => x"51",
          3062 => x"80",
          3063 => x"f9",
          3064 => x"2e",
          3065 => x"98",
          3066 => x"0d",
          3067 => x"05",
          3068 => x"27",
          3069 => x"29",
          3070 => x"82",
          3071 => x"f9",
          3072 => x"54",
          3073 => x"76",
          3074 => x"ff",
          3075 => x"80",
          3076 => x"72",
          3077 => x"72",
          3078 => x"39",
          3079 => x"a8",
          3080 => x"fd",
          3081 => x"9f",
          3082 => x"11",
          3083 => x"18",
          3084 => x"53",
          3085 => x"80",
          3086 => x"b8",
          3087 => x"79",
          3088 => x"58",
          3089 => x"9f",
          3090 => x"88",
          3091 => x"51",
          3092 => x"80",
          3093 => x"74",
          3094 => x"82",
          3095 => x"58",
          3096 => x"08",
          3097 => x"82",
          3098 => x"2b",
          3099 => x"51",
          3100 => x"f0",
          3101 => x"77",
          3102 => x"04",
          3103 => x"58",
          3104 => x"9e",
          3105 => x"96",
          3106 => x"81",
          3107 => x"72",
          3108 => x"72",
          3109 => x"39",
          3110 => x"a8",
          3111 => x"fb",
          3112 => x"82",
          3113 => x"83",
          3114 => x"78",
          3115 => x"76",
          3116 => x"9f",
          3117 => x"07",
          3118 => x"83",
          3119 => x"08",
          3120 => x"82",
          3121 => x"08",
          3122 => x"16",
          3123 => x"76",
          3124 => x"81",
          3125 => x"53",
          3126 => x"88",
          3127 => x"51",
          3128 => x"59",
          3129 => x"77",
          3130 => x"83",
          3131 => x"f6",
          3132 => x"a8",
          3133 => x"ef",
          3134 => x"e0",
          3135 => x"06",
          3136 => x"18",
          3137 => x"f6",
          3138 => x"0a",
          3139 => x"c5",
          3140 => x"82",
          3141 => x"f8",
          3142 => x"59",
          3143 => x"38",
          3144 => x"73",
          3145 => x"52",
          3146 => x"98",
          3147 => x"f2",
          3148 => x"39",
          3149 => x"98",
          3150 => x"78",
          3151 => x"08",
          3152 => x"80",
          3153 => x"2e",
          3154 => x"2e",
          3155 => x"51",
          3156 => x"c5",
          3157 => x"18",
          3158 => x"90",
          3159 => x"16",
          3160 => x"34",
          3161 => x"38",
          3162 => x"8a",
          3163 => x"7e",
          3164 => x"38",
          3165 => x"88",
          3166 => x"38",
          3167 => x"51",
          3168 => x"e0",
          3169 => x"e0",
          3170 => x"ff",
          3171 => x"82",
          3172 => x"79",
          3173 => x"73",
          3174 => x"2e",
          3175 => x"1a",
          3176 => x"38",
          3177 => x"af",
          3178 => x"81",
          3179 => x"e0",
          3180 => x"09",
          3181 => x"70",
          3182 => x"51",
          3183 => x"82",
          3184 => x"90",
          3185 => x"38",
          3186 => x"73",
          3187 => x"77",
          3188 => x"76",
          3189 => x"26",
          3190 => x"f8",
          3191 => x"2e",
          3192 => x"08",
          3193 => x"82",
          3194 => x"08",
          3195 => x"25",
          3196 => x"73",
          3197 => x"81",
          3198 => x"f5",
          3199 => x"f9",
          3200 => x"e0",
          3201 => x"08",
          3202 => x"80",
          3203 => x"38",
          3204 => x"d0",
          3205 => x"a5",
          3206 => x"08",
          3207 => x"74",
          3208 => x"18",
          3209 => x"73",
          3210 => x"74",
          3211 => x"55",
          3212 => x"85",
          3213 => x"e0",
          3214 => x"3d",
          3215 => x"3f",
          3216 => x"82",
          3217 => x"52",
          3218 => x"98",
          3219 => x"0c",
          3220 => x"15",
          3221 => x"56",
          3222 => x"22",
          3223 => x"54",
          3224 => x"33",
          3225 => x"08",
          3226 => x"76",
          3227 => x"9f",
          3228 => x"e0",
          3229 => x"3d",
          3230 => x"57",
          3231 => x"38",
          3232 => x"38",
          3233 => x"54",
          3234 => x"73",
          3235 => x"73",
          3236 => x"0b",
          3237 => x"27",
          3238 => x"18",
          3239 => x"70",
          3240 => x"b2",
          3241 => x"3f",
          3242 => x"98",
          3243 => x"82",
          3244 => x"16",
          3245 => x"38",
          3246 => x"55",
          3247 => x"d5",
          3248 => x"0c",
          3249 => x"53",
          3250 => x"85",
          3251 => x"2a",
          3252 => x"06",
          3253 => x"58",
          3254 => x"0d",
          3255 => x"90",
          3256 => x"f0",
          3257 => x"0b",
          3258 => x"84",
          3259 => x"76",
          3260 => x"38",
          3261 => x"08",
          3262 => x"88",
          3263 => x"81",
          3264 => x"22",
          3265 => x"72",
          3266 => x"f3",
          3267 => x"82",
          3268 => x"27",
          3269 => x"98",
          3270 => x"16",
          3271 => x"ca",
          3272 => x"0c",
          3273 => x"08",
          3274 => x"e0",
          3275 => x"98",
          3276 => x"55",
          3277 => x"38",
          3278 => x"2e",
          3279 => x"75",
          3280 => x"08",
          3281 => x"52",
          3282 => x"98",
          3283 => x"0c",
          3284 => x"80",
          3285 => x"3d",
          3286 => x"71",
          3287 => x"51",
          3288 => x"54",
          3289 => x"82",
          3290 => x"52",
          3291 => x"98",
          3292 => x"d2",
          3293 => x"08",
          3294 => x"e5",
          3295 => x"58",
          3296 => x"38",
          3297 => x"80",
          3298 => x"7a",
          3299 => x"39",
          3300 => x"76",
          3301 => x"08",
          3302 => x"ff",
          3303 => x"06",
          3304 => x"98",
          3305 => x"0d",
          3306 => x"3f",
          3307 => x"06",
          3308 => x"83",
          3309 => x"14",
          3310 => x"08",
          3311 => x"e0",
          3312 => x"3d",
          3313 => x"06",
          3314 => x"af",
          3315 => x"83",
          3316 => x"90",
          3317 => x"3f",
          3318 => x"75",
          3319 => x"2a",
          3320 => x"81",
          3321 => x"ff",
          3322 => x"72",
          3323 => x"85",
          3324 => x"62",
          3325 => x"81",
          3326 => x"80",
          3327 => x"52",
          3328 => x"98",
          3329 => x"eb",
          3330 => x"55",
          3331 => x"39",
          3332 => x"ff",
          3333 => x"82",
          3334 => x"2e",
          3335 => x"82",
          3336 => x"09",
          3337 => x"73",
          3338 => x"98",
          3339 => x"88",
          3340 => x"56",
          3341 => x"5c",
          3342 => x"81",
          3343 => x"70",
          3344 => x"92",
          3345 => x"06",
          3346 => x"56",
          3347 => x"06",
          3348 => x"7c",
          3349 => x"38",
          3350 => x"e8",
          3351 => x"ff",
          3352 => x"74",
          3353 => x"f3",
          3354 => x"82",
          3355 => x"e8",
          3356 => x"ff",
          3357 => x"38",
          3358 => x"73",
          3359 => x"23",
          3360 => x"ff",
          3361 => x"81",
          3362 => x"74",
          3363 => x"51",
          3364 => x"73",
          3365 => x"1a",
          3366 => x"81",
          3367 => x"ff",
          3368 => x"38",
          3369 => x"98",
          3370 => x"2e",
          3371 => x"a0",
          3372 => x"3f",
          3373 => x"98",
          3374 => x"84",
          3375 => x"0c",
          3376 => x"0d",
          3377 => x"40",
          3378 => x"3f",
          3379 => x"98",
          3380 => x"5f",
          3381 => x"19",
          3382 => x"82",
          3383 => x"08",
          3384 => x"33",
          3385 => x"82",
          3386 => x"70",
          3387 => x"1a",
          3388 => x"38",
          3389 => x"54",
          3390 => x"b2",
          3391 => x"81",
          3392 => x"2a",
          3393 => x"82",
          3394 => x"06",
          3395 => x"8d",
          3396 => x"90",
          3397 => x"5e",
          3398 => x"b9",
          3399 => x"2e",
          3400 => x"1f",
          3401 => x"3f",
          3402 => x"06",
          3403 => x"70",
          3404 => x"56",
          3405 => x"1b",
          3406 => x"82",
          3407 => x"56",
          3408 => x"fe",
          3409 => x"e1",
          3410 => x"10",
          3411 => x"59",
          3412 => x"e0",
          3413 => x"c1",
          3414 => x"ff",
          3415 => x"81",
          3416 => x"38",
          3417 => x"06",
          3418 => x"38",
          3419 => x"1d",
          3420 => x"ff",
          3421 => x"84",
          3422 => x"39",
          3423 => x"3f",
          3424 => x"54",
          3425 => x"33",
          3426 => x"53",
          3427 => x"e5",
          3428 => x"2e",
          3429 => x"ac",
          3430 => x"81",
          3431 => x"e0",
          3432 => x"77",
          3433 => x"04",
          3434 => x"12",
          3435 => x"86",
          3436 => x"1d",
          3437 => x"80",
          3438 => x"16",
          3439 => x"8c",
          3440 => x"70",
          3441 => x"80",
          3442 => x"80",
          3443 => x"ab",
          3444 => x"7b",
          3445 => x"51",
          3446 => x"c6",
          3447 => x"ff",
          3448 => x"b4",
          3449 => x"19",
          3450 => x"76",
          3451 => x"2a",
          3452 => x"73",
          3453 => x"a1",
          3454 => x"25",
          3455 => x"02",
          3456 => x"b0",
          3457 => x"84",
          3458 => x"ff",
          3459 => x"58",
          3460 => x"05",
          3461 => x"77",
          3462 => x"a0",
          3463 => x"52",
          3464 => x"08",
          3465 => x"74",
          3466 => x"81",
          3467 => x"74",
          3468 => x"94",
          3469 => x"15",
          3470 => x"87",
          3471 => x"70",
          3472 => x"87",
          3473 => x"f9",
          3474 => x"81",
          3475 => x"84",
          3476 => x"82",
          3477 => x"82",
          3478 => x"06",
          3479 => x"33",
          3480 => x"33",
          3481 => x"55",
          3482 => x"38",
          3483 => x"f4",
          3484 => x"78",
          3485 => x"e0",
          3486 => x"82",
          3487 => x"2e",
          3488 => x"1b",
          3489 => x"ef",
          3490 => x"82",
          3491 => x"1a",
          3492 => x"08",
          3493 => x"52",
          3494 => x"98",
          3495 => x"d7",
          3496 => x"7a",
          3497 => x"8d",
          3498 => x"82",
          3499 => x"e0",
          3500 => x"df",
          3501 => x"55",
          3502 => x"38",
          3503 => x"57",
          3504 => x"17",
          3505 => x"73",
          3506 => x"17",
          3507 => x"83",
          3508 => x"1b",
          3509 => x"77",
          3510 => x"81",
          3511 => x"51",
          3512 => x"57",
          3513 => x"ff",
          3514 => x"1a",
          3515 => x"82",
          3516 => x"08",
          3517 => x"08",
          3518 => x"3f",
          3519 => x"08",
          3520 => x"ab",
          3521 => x"8c",
          3522 => x"76",
          3523 => x"3d",
          3524 => x"08",
          3525 => x"59",
          3526 => x"72",
          3527 => x"e0",
          3528 => x"80",
          3529 => x"51",
          3530 => x"54",
          3531 => x"15",
          3532 => x"83",
          3533 => x"a2",
          3534 => x"51",
          3535 => x"54",
          3536 => x"38",
          3537 => x"38",
          3538 => x"88",
          3539 => x"60",
          3540 => x"96",
          3541 => x"83",
          3542 => x"81",
          3543 => x"05",
          3544 => x"57",
          3545 => x"10",
          3546 => x"53",
          3547 => x"70",
          3548 => x"8f",
          3549 => x"df",
          3550 => x"79",
          3551 => x"7a",
          3552 => x"84",
          3553 => x"ff",
          3554 => x"38",
          3555 => x"2a",
          3556 => x"34",
          3557 => x"30",
          3558 => x"25",
          3559 => x"85",
          3560 => x"34",
          3561 => x"8c",
          3562 => x"51",
          3563 => x"30",
          3564 => x"59",
          3565 => x"80",
          3566 => x"1a",
          3567 => x"70",
          3568 => x"a0",
          3569 => x"81",
          3570 => x"89",
          3571 => x"25",
          3572 => x"38",
          3573 => x"70",
          3574 => x"74",
          3575 => x"17",
          3576 => x"77",
          3577 => x"14",
          3578 => x"87",
          3579 => x"19",
          3580 => x"73",
          3581 => x"80",
          3582 => x"19",
          3583 => x"54",
          3584 => x"1c",
          3585 => x"79",
          3586 => x"85",
          3587 => x"06",
          3588 => x"15",
          3589 => x"74",
          3590 => x"19",
          3591 => x"59",
          3592 => x"17",
          3593 => x"34",
          3594 => x"53",
          3595 => x"9c",
          3596 => x"19",
          3597 => x"53",
          3598 => x"78",
          3599 => x"82",
          3600 => x"13",
          3601 => x"08",
          3602 => x"f0",
          3603 => x"80",
          3604 => x"af",
          3605 => x"dc",
          3606 => x"38",
          3607 => x"aa",
          3608 => x"33",
          3609 => x"81",
          3610 => x"dc",
          3611 => x"07",
          3612 => x"88",
          3613 => x"73",
          3614 => x"ab",
          3615 => x"ee",
          3616 => x"e1",
          3617 => x"08",
          3618 => x"05",
          3619 => x"08",
          3620 => x"ff",
          3621 => x"38",
          3622 => x"90",
          3623 => x"19",
          3624 => x"ff",
          3625 => x"73",
          3626 => x"55",
          3627 => x"2e",
          3628 => x"38",
          3629 => x"92",
          3630 => x"38",
          3631 => x"78",
          3632 => x"19",
          3633 => x"80",
          3634 => x"af",
          3635 => x"57",
          3636 => x"80",
          3637 => x"dc",
          3638 => x"2b",
          3639 => x"8c",
          3640 => x"a5",
          3641 => x"09",
          3642 => x"22",
          3643 => x"80",
          3644 => x"2e",
          3645 => x"1a",
          3646 => x"1f",
          3647 => x"83",
          3648 => x"05",
          3649 => x"27",
          3650 => x"ab",
          3651 => x"2e",
          3652 => x"55",
          3653 => x"32",
          3654 => x"53",
          3655 => x"38",
          3656 => x"e0",
          3657 => x"80",
          3658 => x"85",
          3659 => x"99",
          3660 => x"ff",
          3661 => x"09",
          3662 => x"10",
          3663 => x"a0",
          3664 => x"83",
          3665 => x"09",
          3666 => x"57",
          3667 => x"fe",
          3668 => x"2e",
          3669 => x"55",
          3670 => x"38",
          3671 => x"ae",
          3672 => x"53",
          3673 => x"3f",
          3674 => x"10",
          3675 => x"54",
          3676 => x"a0",
          3677 => x"30",
          3678 => x"79",
          3679 => x"38",
          3680 => x"54",
          3681 => x"81",
          3682 => x"72",
          3683 => x"51",
          3684 => x"7e",
          3685 => x"2e",
          3686 => x"79",
          3687 => x"58",
          3688 => x"5d",
          3689 => x"27",
          3690 => x"b5",
          3691 => x"82",
          3692 => x"70",
          3693 => x"56",
          3694 => x"ff",
          3695 => x"54",
          3696 => x"1f",
          3697 => x"83",
          3698 => x"7d",
          3699 => x"55",
          3700 => x"c3",
          3701 => x"52",
          3702 => x"82",
          3703 => x"80",
          3704 => x"39",
          3705 => x"85",
          3706 => x"16",
          3707 => x"81",
          3708 => x"06",
          3709 => x"54",
          3710 => x"de",
          3711 => x"e5",
          3712 => x"0b",
          3713 => x"81",
          3714 => x"fc",
          3715 => x"8c",
          3716 => x"73",
          3717 => x"76",
          3718 => x"81",
          3719 => x"81",
          3720 => x"76",
          3721 => x"81",
          3722 => x"38",
          3723 => x"34",
          3724 => x"98",
          3725 => x"e0",
          3726 => x"e0",
          3727 => x"80",
          3728 => x"06",
          3729 => x"80",
          3730 => x"73",
          3731 => x"0b",
          3732 => x"39",
          3733 => x"85",
          3734 => x"81",
          3735 => x"1e",
          3736 => x"51",
          3737 => x"90",
          3738 => x"b8",
          3739 => x"82",
          3740 => x"a1",
          3741 => x"3d",
          3742 => x"ff",
          3743 => x"5c",
          3744 => x"38",
          3745 => x"9f",
          3746 => x"38",
          3747 => x"81",
          3748 => x"11",
          3749 => x"70",
          3750 => x"81",
          3751 => x"76",
          3752 => x"d2",
          3753 => x"57",
          3754 => x"70",
          3755 => x"53",
          3756 => x"e0",
          3757 => x"ff",
          3758 => x"38",
          3759 => x"51",
          3760 => x"72",
          3761 => x"70",
          3762 => x"32",
          3763 => x"73",
          3764 => x"70",
          3765 => x"19",
          3766 => x"38",
          3767 => x"74",
          3768 => x"39",
          3769 => x"e0",
          3770 => x"3d",
          3771 => x"34",
          3772 => x"75",
          3773 => x"e0",
          3774 => x"16",
          3775 => x"08",
          3776 => x"73",
          3777 => x"80",
          3778 => x"56",
          3779 => x"06",
          3780 => x"32",
          3781 => x"51",
          3782 => x"e8",
          3783 => x"53",
          3784 => x"51",
          3785 => x"55",
          3786 => x"38",
          3787 => x"8a",
          3788 => x"98",
          3789 => x"2e",
          3790 => x"98",
          3791 => x"0d",
          3792 => x"33",
          3793 => x"fc",
          3794 => x"8b",
          3795 => x"24",
          3796 => x"84",
          3797 => x"55",
          3798 => x"b1",
          3799 => x"06",
          3800 => x"ae",
          3801 => x"3f",
          3802 => x"70",
          3803 => x"76",
          3804 => x"2a",
          3805 => x"72",
          3806 => x"74",
          3807 => x"19",
          3808 => x"14",
          3809 => x"98",
          3810 => x"54",
          3811 => x"76",
          3812 => x"70",
          3813 => x"86",
          3814 => x"5b",
          3815 => x"81",
          3816 => x"38",
          3817 => x"e0",
          3818 => x"81",
          3819 => x"83",
          3820 => x"53",
          3821 => x"15",
          3822 => x"08",
          3823 => x"0c",
          3824 => x"80",
          3825 => x"8d",
          3826 => x"72",
          3827 => x"05",
          3828 => x"59",
          3829 => x"2e",
          3830 => x"9e",
          3831 => x"06",
          3832 => x"33",
          3833 => x"06",
          3834 => x"91",
          3835 => x"16",
          3836 => x"c0",
          3837 => x"f9",
          3838 => x"f1",
          3839 => x"3f",
          3840 => x"06",
          3841 => x"06",
          3842 => x"c9",
          3843 => x"ff",
          3844 => x"dc",
          3845 => x"98",
          3846 => x"c8",
          3847 => x"14",
          3848 => x"51",
          3849 => x"84",
          3850 => x"71",
          3851 => x"53",
          3852 => x"8b",
          3853 => x"80",
          3854 => x"39",
          3855 => x"82",
          3856 => x"08",
          3857 => x"8d",
          3858 => x"14",
          3859 => x"08",
          3860 => x"38",
          3861 => x"82",
          3862 => x"51",
          3863 => x"83",
          3864 => x"80",
          3865 => x"78",
          3866 => x"78",
          3867 => x"22",
          3868 => x"ec",
          3869 => x"e0",
          3870 => x"82",
          3871 => x"f5",
          3872 => x"ff",
          3873 => x"9f",
          3874 => x"39",
          3875 => x"38",
          3876 => x"a4",
          3877 => x"0c",
          3878 => x"76",
          3879 => x"80",
          3880 => x"e0",
          3881 => x"8d",
          3882 => x"91",
          3883 => x"3f",
          3884 => x"74",
          3885 => x"79",
          3886 => x"ac",
          3887 => x"2e",
          3888 => x"2a",
          3889 => x"ff",
          3890 => x"a0",
          3891 => x"0b",
          3892 => x"0c",
          3893 => x"83",
          3894 => x"80",
          3895 => x"e0",
          3896 => x"72",
          3897 => x"38",
          3898 => x"3f",
          3899 => x"82",
          3900 => x"b6",
          3901 => x"98",
          3902 => x"82",
          3903 => x"c8",
          3904 => x"82",
          3905 => x"d2",
          3906 => x"9c",
          3907 => x"98",
          3908 => x"09",
          3909 => x"51",
          3910 => x"94",
          3911 => x"dc",
          3912 => x"0c",
          3913 => x"81",
          3914 => x"72",
          3915 => x"8c",
          3916 => x"80",
          3917 => x"3d",
          3918 => x"89",
          3919 => x"08",
          3920 => x"33",
          3921 => x"13",
          3922 => x"76",
          3923 => x"13",
          3924 => x"e0",
          3925 => x"38",
          3926 => x"80",
          3927 => x"82",
          3928 => x"fa",
          3929 => x"58",
          3930 => x"9a",
          3931 => x"98",
          3932 => x"08",
          3933 => x"08",
          3934 => x"80",
          3935 => x"84",
          3936 => x"75",
          3937 => x"53",
          3938 => x"f6",
          3939 => x"73",
          3940 => x"04",
          3941 => x"80",
          3942 => x"78",
          3943 => x"06",
          3944 => x"9a",
          3945 => x"3f",
          3946 => x"98",
          3947 => x"52",
          3948 => x"3f",
          3949 => x"98",
          3950 => x"33",
          3951 => x"25",
          3952 => x"54",
          3953 => x"80",
          3954 => x"81",
          3955 => x"3f",
          3956 => x"02",
          3957 => x"81",
          3958 => x"06",
          3959 => x"88",
          3960 => x"58",
          3961 => x"70",
          3962 => x"81",
          3963 => x"ed",
          3964 => x"88",
          3965 => x"c2",
          3966 => x"15",
          3967 => x"d7",
          3968 => x"51",
          3969 => x"83",
          3970 => x"38",
          3971 => x"53",
          3972 => x"cc",
          3973 => x"82",
          3974 => x"39",
          3975 => x"33",
          3976 => x"55",
          3977 => x"55",
          3978 => x"81",
          3979 => x"38",
          3980 => x"a0",
          3981 => x"52",
          3982 => x"98",
          3983 => x"55",
          3984 => x"38",
          3985 => x"54",
          3986 => x"c0",
          3987 => x"1b",
          3988 => x"70",
          3989 => x"98",
          3990 => x"0c",
          3991 => x"3f",
          3992 => x"08",
          3993 => x"86",
          3994 => x"1a",
          3995 => x"0b",
          3996 => x"0c",
          3997 => x"54",
          3998 => x"e0",
          3999 => x"82",
          4000 => x"17",
          4001 => x"57",
          4002 => x"e7",
          4003 => x"e0",
          4004 => x"55",
          4005 => x"81",
          4006 => x"31",
          4007 => x"25",
          4008 => x"81",
          4009 => x"38",
          4010 => x"75",
          4011 => x"a2",
          4012 => x"3f",
          4013 => x"55",
          4014 => x"98",
          4015 => x"80",
          4016 => x"98",
          4017 => x"0d",
          4018 => x"59",
          4019 => x"52",
          4020 => x"98",
          4021 => x"38",
          4022 => x"86",
          4023 => x"19",
          4024 => x"80",
          4025 => x"0b",
          4026 => x"39",
          4027 => x"82",
          4028 => x"08",
          4029 => x"74",
          4030 => x"94",
          4031 => x"56",
          4032 => x"22",
          4033 => x"55",
          4034 => x"19",
          4035 => x"52",
          4036 => x"98",
          4037 => x"38",
          4038 => x"98",
          4039 => x"51",
          4040 => x"80",
          4041 => x"08",
          4042 => x"80",
          4043 => x"8a",
          4044 => x"27",
          4045 => x"54",
          4046 => x"51",
          4047 => x"08",
          4048 => x"56",
          4049 => x"16",
          4050 => x"95",
          4051 => x"b4",
          4052 => x"05",
          4053 => x"2b",
          4054 => x"94",
          4055 => x"71",
          4056 => x"38",
          4057 => x"51",
          4058 => x"fd",
          4059 => x"83",
          4060 => x"51",
          4061 => x"7e",
          4062 => x"1b",
          4063 => x"fd",
          4064 => x"98",
          4065 => x"0d",
          4066 => x"58",
          4067 => x"52",
          4068 => x"98",
          4069 => x"38",
          4070 => x"86",
          4071 => x"18",
          4072 => x"51",
          4073 => x"83",
          4074 => x"19",
          4075 => x"0b",
          4076 => x"39",
          4077 => x"74",
          4078 => x"7b",
          4079 => x"08",
          4080 => x"82",
          4081 => x"05",
          4082 => x"bf",
          4083 => x"55",
          4084 => x"98",
          4085 => x"3f",
          4086 => x"98",
          4087 => x"81",
          4088 => x"ff",
          4089 => x"18",
          4090 => x"7e",
          4091 => x"2e",
          4092 => x"ff",
          4093 => x"fe",
          4094 => x"51",
          4095 => x"08",
          4096 => x"98",
          4097 => x"78",
          4098 => x"7f",
          4099 => x"75",
          4100 => x"78",
          4101 => x"33",
          4102 => x"98",
          4103 => x"08",
          4104 => x"9c",
          4105 => x"77",
          4106 => x"16",
          4107 => x"80",
          4108 => x"56",
          4109 => x"19",
          4110 => x"bb",
          4111 => x"de",
          4112 => x"76",
          4113 => x"ff",
          4114 => x"7b",
          4115 => x"18",
          4116 => x"3f",
          4117 => x"75",
          4118 => x"ff",
          4119 => x"d4",
          4120 => x"34",
          4121 => x"0c",
          4122 => x"94",
          4123 => x"5e",
          4124 => x"55",
          4125 => x"90",
          4126 => x"90",
          4127 => x"98",
          4128 => x"0d",
          4129 => x"52",
          4130 => x"08",
          4131 => x"38",
          4132 => x"81",
          4133 => x"80",
          4134 => x"51",
          4135 => x"08",
          4136 => x"38",
          4137 => x"07",
          4138 => x"16",
          4139 => x"cc",
          4140 => x"15",
          4141 => x"b2",
          4142 => x"ed",
          4143 => x"b7",
          4144 => x"15",
          4145 => x"82",
          4146 => x"bf",
          4147 => x"76",
          4148 => x"04",
          4149 => x"fe",
          4150 => x"82",
          4151 => x"fc",
          4152 => x"82",
          4153 => x"08",
          4154 => x"0c",
          4155 => x"0d",
          4156 => x"e6",
          4157 => x"e0",
          4158 => x"98",
          4159 => x"71",
          4160 => x"04",
          4161 => x"cc",
          4162 => x"3f",
          4163 => x"98",
          4164 => x"52",
          4165 => x"3f",
          4166 => x"98",
          4167 => x"33",
          4168 => x"25",
          4169 => x"54",
          4170 => x"84",
          4171 => x"73",
          4172 => x"70",
          4173 => x"98",
          4174 => x"e0",
          4175 => x"83",
          4176 => x"0c",
          4177 => x"0d",
          4178 => x"08",
          4179 => x"80",
          4180 => x"e0",
          4181 => x"98",
          4182 => x"a1",
          4183 => x"7c",
          4184 => x"55",
          4185 => x"80",
          4186 => x"d3",
          4187 => x"82",
          4188 => x"08",
          4189 => x"52",
          4190 => x"e0",
          4191 => x"82",
          4192 => x"7b",
          4193 => x"08",
          4194 => x"51",
          4195 => x"57",
          4196 => x"80",
          4197 => x"e0",
          4198 => x"a7",
          4199 => x"51",
          4200 => x"08",
          4201 => x"c4",
          4202 => x"82",
          4203 => x"76",
          4204 => x"82",
          4205 => x"38",
          4206 => x"74",
          4207 => x"78",
          4208 => x"56",
          4209 => x"c6",
          4210 => x"33",
          4211 => x"16",
          4212 => x"75",
          4213 => x"05",
          4214 => x"11",
          4215 => x"58",
          4216 => x"ff",
          4217 => x"58",
          4218 => x"7b",
          4219 => x"18",
          4220 => x"af",
          4221 => x"33",
          4222 => x"70",
          4223 => x"56",
          4224 => x"70",
          4225 => x"f5",
          4226 => x"a7",
          4227 => x"38",
          4228 => x"81",
          4229 => x"39",
          4230 => x"74",
          4231 => x"91",
          4232 => x"18",
          4233 => x"70",
          4234 => x"eb",
          4235 => x"98",
          4236 => x"3d",
          4237 => x"54",
          4238 => x"82",
          4239 => x"08",
          4240 => x"72",
          4241 => x"73",
          4242 => x"70",
          4243 => x"57",
          4244 => x"08",
          4245 => x"75",
          4246 => x"11",
          4247 => x"73",
          4248 => x"16",
          4249 => x"98",
          4250 => x"55",
          4251 => x"98",
          4252 => x"70",
          4253 => x"71",
          4254 => x"53",
          4255 => x"a7",
          4256 => x"d3",
          4257 => x"e0",
          4258 => x"82",
          4259 => x"38",
          4260 => x"73",
          4261 => x"9f",
          4262 => x"75",
          4263 => x"17",
          4264 => x"70",
          4265 => x"80",
          4266 => x"ff",
          4267 => x"54",
          4268 => x"e0",
          4269 => x"74",
          4270 => x"98",
          4271 => x"81",
          4272 => x"9c",
          4273 => x"16",
          4274 => x"16",
          4275 => x"53",
          4276 => x"79",
          4277 => x"98",
          4278 => x"34",
          4279 => x"91",
          4280 => x"89",
          4281 => x"94",
          4282 => x"27",
          4283 => x"15",
          4284 => x"16",
          4285 => x"80",
          4286 => x"2e",
          4287 => x"53",
          4288 => x"0d",
          4289 => x"54",
          4290 => x"53",
          4291 => x"84",
          4292 => x"98",
          4293 => x"eb",
          4294 => x"51",
          4295 => x"55",
          4296 => x"ab",
          4297 => x"80",
          4298 => x"70",
          4299 => x"57",
          4300 => x"08",
          4301 => x"e0",
          4302 => x"86",
          4303 => x"75",
          4304 => x"98",
          4305 => x"06",
          4306 => x"80",
          4307 => x"54",
          4308 => x"0d",
          4309 => x"fc",
          4310 => x"3f",
          4311 => x"e0",
          4312 => x"04",
          4313 => x"fc",
          4314 => x"9a",
          4315 => x"e0",
          4316 => x"38",
          4317 => x"ff",
          4318 => x"53",
          4319 => x"52",
          4320 => x"98",
          4321 => x"2e",
          4322 => x"87",
          4323 => x"74",
          4324 => x"52",
          4325 => x"e0",
          4326 => x"72",
          4327 => x"08",
          4328 => x"e0",
          4329 => x"3d",
          4330 => x"70",
          4331 => x"3f",
          4332 => x"98",
          4333 => x"d2",
          4334 => x"82",
          4335 => x"cb",
          4336 => x"73",
          4337 => x"39",
          4338 => x"75",
          4339 => x"98",
          4340 => x"0d",
          4341 => x"3d",
          4342 => x"c5",
          4343 => x"e0",
          4344 => x"0c",
          4345 => x"94",
          4346 => x"74",
          4347 => x"e6",
          4348 => x"5b",
          4349 => x"75",
          4350 => x"81",
          4351 => x"57",
          4352 => x"ff",
          4353 => x"ff",
          4354 => x"81",
          4355 => x"30",
          4356 => x"25",
          4357 => x"5a",
          4358 => x"38",
          4359 => x"e0",
          4360 => x"77",
          4361 => x"ad",
          4362 => x"82",
          4363 => x"70",
          4364 => x"56",
          4365 => x"9e",
          4366 => x"3f",
          4367 => x"06",
          4368 => x"19",
          4369 => x"14",
          4370 => x"98",
          4371 => x"80",
          4372 => x"54",
          4373 => x"79",
          4374 => x"79",
          4375 => x"07",
          4376 => x"82",
          4377 => x"f9",
          4378 => x"53",
          4379 => x"e0",
          4380 => x"81",
          4381 => x"81",
          4382 => x"2a",
          4383 => x"55",
          4384 => x"17",
          4385 => x"81",
          4386 => x"98",
          4387 => x"51",
          4388 => x"08",
          4389 => x"39",
          4390 => x"ad",
          4391 => x"2e",
          4392 => x"82",
          4393 => x"06",
          4394 => x"a1",
          4395 => x"9c",
          4396 => x"08",
          4397 => x"51",
          4398 => x"08",
          4399 => x"90",
          4400 => x"90",
          4401 => x"75",
          4402 => x"e0",
          4403 => x"3d",
          4404 => x"05",
          4405 => x"82",
          4406 => x"08",
          4407 => x"08",
          4408 => x"cf",
          4409 => x"e0",
          4410 => x"ff",
          4411 => x"06",
          4412 => x"cb",
          4413 => x"24",
          4414 => x"33",
          4415 => x"76",
          4416 => x"ff",
          4417 => x"74",
          4418 => x"56",
          4419 => x"54",
          4420 => x"2e",
          4421 => x"98",
          4422 => x"52",
          4423 => x"98",
          4424 => x"eb",
          4425 => x"51",
          4426 => x"08",
          4427 => x"87",
          4428 => x"08",
          4429 => x"08",
          4430 => x"3f",
          4431 => x"08",
          4432 => x"80",
          4433 => x"95",
          4434 => x"53",
          4435 => x"3f",
          4436 => x"38",
          4437 => x"e0",
          4438 => x"0c",
          4439 => x"82",
          4440 => x"9b",
          4441 => x"98",
          4442 => x"b7",
          4443 => x"70",
          4444 => x"98",
          4445 => x"38",
          4446 => x"98",
          4447 => x"8f",
          4448 => x"85",
          4449 => x"74",
          4450 => x"8a",
          4451 => x"3f",
          4452 => x"82",
          4453 => x"82",
          4454 => x"06",
          4455 => x"08",
          4456 => x"81",
          4457 => x"38",
          4458 => x"ff",
          4459 => x"54",
          4460 => x"8b",
          4461 => x"a4",
          4462 => x"15",
          4463 => x"15",
          4464 => x"ce",
          4465 => x"53",
          4466 => x"ee",
          4467 => x"80",
          4468 => x"78",
          4469 => x"7f",
          4470 => x"ff",
          4471 => x"83",
          4472 => x"3f",
          4473 => x"98",
          4474 => x"52",
          4475 => x"3f",
          4476 => x"b7",
          4477 => x"15",
          4478 => x"34",
          4479 => x"e0",
          4480 => x"75",
          4481 => x"73",
          4482 => x"04",
          4483 => x"51",
          4484 => x"fe",
          4485 => x"cd",
          4486 => x"e0",
          4487 => x"ab",
          4488 => x"58",
          4489 => x"55",
          4490 => x"02",
          4491 => x"54",
          4492 => x"53",
          4493 => x"80",
          4494 => x"53",
          4495 => x"ff",
          4496 => x"73",
          4497 => x"08",
          4498 => x"63",
          4499 => x"88",
          4500 => x"38",
          4501 => x"98",
          4502 => x"bb",
          4503 => x"82",
          4504 => x"08",
          4505 => x"aa",
          4506 => x"51",
          4507 => x"33",
          4508 => x"84",
          4509 => x"73",
          4510 => x"8b",
          4511 => x"15",
          4512 => x"70",
          4513 => x"2e",
          4514 => x"e1",
          4515 => x"ad",
          4516 => x"51",
          4517 => x"e0",
          4518 => x"82",
          4519 => x"a3",
          4520 => x"80",
          4521 => x"98",
          4522 => x"54",
          4523 => x"38",
          4524 => x"b4",
          4525 => x"15",
          4526 => x"9c",
          4527 => x"e0",
          4528 => x"8c",
          4529 => x"82",
          4530 => x"98",
          4531 => x"0d",
          4532 => x"05",
          4533 => x"53",
          4534 => x"51",
          4535 => x"55",
          4536 => x"78",
          4537 => x"51",
          4538 => x"55",
          4539 => x"80",
          4540 => x"86",
          4541 => x"61",
          4542 => x"7a",
          4543 => x"74",
          4544 => x"83",
          4545 => x"3f",
          4546 => x"e0",
          4547 => x"3d",
          4548 => x"cc",
          4549 => x"3f",
          4550 => x"98",
          4551 => x"52",
          4552 => x"3f",
          4553 => x"98",
          4554 => x"33",
          4555 => x"a6",
          4556 => x"71",
          4557 => x"51",
          4558 => x"0b",
          4559 => x"a6",
          4560 => x"82",
          4561 => x"e9",
          4562 => x"53",
          4563 => x"51",
          4564 => x"82",
          4565 => x"98",
          4566 => x"79",
          4567 => x"75",
          4568 => x"fa",
          4569 => x"8d",
          4570 => x"3f",
          4571 => x"98",
          4572 => x"51",
          4573 => x"08",
          4574 => x"82",
          4575 => x"65",
          4576 => x"7b",
          4577 => x"34",
          4578 => x"38",
          4579 => x"34",
          4580 => x"70",
          4581 => x"a0",
          4582 => x"2e",
          4583 => x"34",
          4584 => x"80",
          4585 => x"c1",
          4586 => x"a4",
          4587 => x"3f",
          4588 => x"98",
          4589 => x"55",
          4590 => x"38",
          4591 => x"38",
          4592 => x"ff",
          4593 => x"7b",
          4594 => x"3d",
          4595 => x"9c",
          4596 => x"51",
          4597 => x"82",
          4598 => x"98",
          4599 => x"52",
          4600 => x"ef",
          4601 => x"56",
          4602 => x"57",
          4603 => x"82",
          4604 => x"80",
          4605 => x"96",
          4606 => x"98",
          4607 => x"98",
          4608 => x"80",
          4609 => x"b8",
          4610 => x"98",
          4611 => x"88",
          4612 => x"39",
          4613 => x"81",
          4614 => x"38",
          4615 => x"81",
          4616 => x"77",
          4617 => x"6d",
          4618 => x"26",
          4619 => x"86",
          4620 => x"38",
          4621 => x"05",
          4622 => x"73",
          4623 => x"ff",
          4624 => x"80",
          4625 => x"55",
          4626 => x"08",
          4627 => x"38",
          4628 => x"3f",
          4629 => x"98",
          4630 => x"66",
          4631 => x"82",
          4632 => x"06",
          4633 => x"2e",
          4634 => x"ff",
          4635 => x"54",
          4636 => x"53",
          4637 => x"ff",
          4638 => x"8b",
          4639 => x"51",
          4640 => x"0b",
          4641 => x"96",
          4642 => x"55",
          4643 => x"0d",
          4644 => x"88",
          4645 => x"fc",
          4646 => x"d2",
          4647 => x"82",
          4648 => x"1a",
          4649 => x"80",
          4650 => x"78",
          4651 => x"2a",
          4652 => x"90",
          4653 => x"58",
          4654 => x"39",
          4655 => x"70",
          4656 => x"a2",
          4657 => x"30",
          4658 => x"98",
          4659 => x"5a",
          4660 => x"38",
          4661 => x"82",
          4662 => x"74",
          4663 => x"81",
          4664 => x"75",
          4665 => x"98",
          4666 => x"e0",
          4667 => x"82",
          4668 => x"56",
          4669 => x"38",
          4670 => x"77",
          4671 => x"87",
          4672 => x"ba",
          4673 => x"2e",
          4674 => x"2e",
          4675 => x"75",
          4676 => x"d0",
          4677 => x"e0",
          4678 => x"16",
          4679 => x"38",
          4680 => x"90",
          4681 => x"38",
          4682 => x"0c",
          4683 => x"73",
          4684 => x"05",
          4685 => x"26",
          4686 => x"0c",
          4687 => x"84",
          4688 => x"98",
          4689 => x"0d",
          4690 => x"05",
          4691 => x"c4",
          4692 => x"e0",
          4693 => x"e0",
          4694 => x"05",
          4695 => x"84",
          4696 => x"08",
          4697 => x"8c",
          4698 => x"47",
          4699 => x"8e",
          4700 => x"ff",
          4701 => x"56",
          4702 => x"70",
          4703 => x"8c",
          4704 => x"83",
          4705 => x"82",
          4706 => x"74",
          4707 => x"80",
          4708 => x"55",
          4709 => x"78",
          4710 => x"26",
          4711 => x"8b",
          4712 => x"80",
          4713 => x"39",
          4714 => x"89",
          4715 => x"83",
          4716 => x"25",
          4717 => x"8b",
          4718 => x"38",
          4719 => x"51",
          4720 => x"e0",
          4721 => x"1b",
          4722 => x"98",
          4723 => x"56",
          4724 => x"06",
          4725 => x"83",
          4726 => x"2e",
          4727 => x"ff",
          4728 => x"83",
          4729 => x"3f",
          4730 => x"9a",
          4731 => x"51",
          4732 => x"e0",
          4733 => x"2a",
          4734 => x"41",
          4735 => x"67",
          4736 => x"c5",
          4737 => x"80",
          4738 => x"56",
          4739 => x"62",
          4740 => x"74",
          4741 => x"55",
          4742 => x"81",
          4743 => x"38",
          4744 => x"5e",
          4745 => x"5a",
          4746 => x"e1",
          4747 => x"57",
          4748 => x"5a",
          4749 => x"26",
          4750 => x"10",
          4751 => x"74",
          4752 => x"ee",
          4753 => x"c4",
          4754 => x"84",
          4755 => x"a0",
          4756 => x"fc",
          4757 => x"f0",
          4758 => x"88",
          4759 => x"57",
          4760 => x"5a",
          4761 => x"26",
          4762 => x"10",
          4763 => x"74",
          4764 => x"ee",
          4765 => x"e4",
          4766 => x"05",
          4767 => x"26",
          4768 => x"08",
          4769 => x"11",
          4770 => x"83",
          4771 => x"a0",
          4772 => x"6a",
          4773 => x"72",
          4774 => x"59",
          4775 => x"89",
          4776 => x"84",
          4777 => x"18",
          4778 => x"74",
          4779 => x"31",
          4780 => x"52",
          4781 => x"98",
          4782 => x"06",
          4783 => x"ff",
          4784 => x"b8",
          4785 => x"be",
          4786 => x"09",
          4787 => x"f5",
          4788 => x"38",
          4789 => x"80",
          4790 => x"96",
          4791 => x"2e",
          4792 => x"82",
          4793 => x"38",
          4794 => x"81",
          4795 => x"e0",
          4796 => x"81",
          4797 => x"78",
          4798 => x"8e",
          4799 => x"53",
          4800 => x"3f",
          4801 => x"51",
          4802 => x"8b",
          4803 => x"8d",
          4804 => x"52",
          4805 => x"81",
          4806 => x"70",
          4807 => x"54",
          4808 => x"ff",
          4809 => x"26",
          4810 => x"52",
          4811 => x"8a",
          4812 => x"8d",
          4813 => x"bf",
          4814 => x"3f",
          4815 => x"8d",
          4816 => x"ff",
          4817 => x"81",
          4818 => x"0a",
          4819 => x"c5",
          4820 => x"8d",
          4821 => x"ff",
          4822 => x"51",
          4823 => x"1b",
          4824 => x"0b",
          4825 => x"c2",
          4826 => x"52",
          4827 => x"88",
          4828 => x"8c",
          4829 => x"52",
          4830 => x"ff",
          4831 => x"a6",
          4832 => x"52",
          4833 => x"82",
          4834 => x"52",
          4835 => x"7e",
          4836 => x"ce",
          4837 => x"84",
          4838 => x"06",
          4839 => x"53",
          4840 => x"3f",
          4841 => x"ff",
          4842 => x"d2",
          4843 => x"86",
          4844 => x"1b",
          4845 => x"52",
          4846 => x"3f",
          4847 => x"8b",
          4848 => x"51",
          4849 => x"1f",
          4850 => x"de",
          4851 => x"52",
          4852 => x"53",
          4853 => x"3f",
          4854 => x"09",
          4855 => x"51",
          4856 => x"1b",
          4857 => x"52",
          4858 => x"ff",
          4859 => x"f8",
          4860 => x"fd",
          4861 => x"26",
          4862 => x"53",
          4863 => x"3f",
          4864 => x"84",
          4865 => x"7a",
          4866 => x"75",
          4867 => x"81",
          4868 => x"38",
          4869 => x"65",
          4870 => x"38",
          4871 => x"52",
          4872 => x"e0",
          4873 => x"75",
          4874 => x"8c",
          4875 => x"57",
          4876 => x"84",
          4877 => x"57",
          4878 => x"80",
          4879 => x"8c",
          4880 => x"81",
          4881 => x"76",
          4882 => x"e0",
          4883 => x"ff",
          4884 => x"83",
          4885 => x"38",
          4886 => x"ff",
          4887 => x"78",
          4888 => x"1b",
          4889 => x"16",
          4890 => x"83",
          4891 => x"1f",
          4892 => x"fe",
          4893 => x"34",
          4894 => x"07",
          4895 => x"98",
          4896 => x"c6",
          4897 => x"52",
          4898 => x"3f",
          4899 => x"51",
          4900 => x"e0",
          4901 => x"52",
          4902 => x"56",
          4903 => x"39",
          4904 => x"39",
          4905 => x"e0",
          4906 => x"3d",
          4907 => x"60",
          4908 => x"25",
          4909 => x"55",
          4910 => x"c8",
          4911 => x"06",
          4912 => x"8d",
          4913 => x"05",
          4914 => x"2e",
          4915 => x"34",
          4916 => x"74",
          4917 => x"04",
          4918 => x"b3",
          4919 => x"09",
          4920 => x"51",
          4921 => x"76",
          4922 => x"17",
          4923 => x"81",
          4924 => x"8b",
          4925 => x"17",
          4926 => x"79",
          4927 => x"9f",
          4928 => x"75",
          4929 => x"0c",
          4930 => x"79",
          4931 => x"24",
          4932 => x"74",
          4933 => x"c9",
          4934 => x"38",
          4935 => x"06",
          4936 => x"39",
          4937 => x"89",
          4938 => x"54",
          4939 => x"ff",
          4940 => x"3d",
          4941 => x"e3",
          4942 => x"53",
          4943 => x"51",
          4944 => x"3f",
          4945 => x"75",
          4946 => x"53",
          4947 => x"38",
          4948 => x"c3",
          4949 => x"73",
          4950 => x"38",
          4951 => x"ec",
          4952 => x"81",
          4953 => x"51",
          4954 => x"10",
          4955 => x"51",
          4956 => x"ff",
          4957 => x"0c",
          4958 => x"02",
          4959 => x"05",
          4960 => x"ff",
          4961 => x"71",
          4962 => x"38",
          4963 => x"10",
          4964 => x"51",
          4965 => x"0d",
          4966 => x"83",
          4967 => x"83",
          4968 => x"52",
          4969 => x"d9",
          4970 => x"22",
          4971 => x"26",
          4972 => x"38",
          4973 => x"88",
          4974 => x"54",
          4975 => x"d7",
          4976 => x"73",
          4977 => x"70",
          4978 => x"11",
          4979 => x"39",
          4980 => x"31",
          4981 => x"9f",
          4982 => x"12",
          4983 => x"39",
          4984 => x"12",
          4985 => x"70",
          4986 => x"73",
          4987 => x"fe",
          4988 => x"98",
          4989 => x"ff",
          4990 => x"00",
          4991 => x"31",
          4992 => x"30",
          4993 => x"30",
          4994 => x"30",
          4995 => x"30",
          4996 => x"30",
          4997 => x"30",
          4998 => x"30",
          4999 => x"30",
          5000 => x"30",
          5001 => x"47",
          5002 => x"47",
          5003 => x"47",
          5004 => x"4e",
          5005 => x"51",
          5006 => x"4c",
          5007 => x"51",
          5008 => x"51",
          5009 => x"4f",
          5010 => x"4f",
          5011 => x"50",
          5012 => x"4c",
          5013 => x"51",
          5014 => x"51",
          5015 => x"9b",
          5016 => x"9b",
          5017 => x"9b",
          5018 => x"9b",
          5019 => x"0e",
          5020 => x"17",
          5021 => x"17",
          5022 => x"17",
          5023 => x"17",
          5024 => x"17",
          5025 => x"17",
          5026 => x"0e",
          5027 => x"17",
          5028 => x"17",
          5029 => x"17",
          5030 => x"17",
          5031 => x"17",
          5032 => x"17",
          5033 => x"17",
          5034 => x"17",
          5035 => x"17",
          5036 => x"17",
          5037 => x"17",
          5038 => x"17",
          5039 => x"17",
          5040 => x"17",
          5041 => x"17",
          5042 => x"17",
          5043 => x"17",
          5044 => x"17",
          5045 => x"17",
          5046 => x"17",
          5047 => x"11",
          5048 => x"17",
          5049 => x"17",
          5050 => x"17",
          5051 => x"17",
          5052 => x"17",
          5053 => x"10",
          5054 => x"0e",
          5055 => x"17",
          5056 => x"17",
          5057 => x"0e",
          5058 => x"17",
          5059 => x"11",
          5060 => x"17",
          5061 => x"17",
          5062 => x"17",
          5063 => x"11",
          5064 => x"00",
          5065 => x"00",
          5066 => x"00",
          5067 => x"00",
          5068 => x"00",
          5069 => x"00",
          5070 => x"00",
          5071 => x"00",
          5072 => x"00",
          5073 => x"68",
          5074 => x"64",
          5075 => x"64",
          5076 => x"6c",
          5077 => x"70",
          5078 => x"74",
          5079 => x"00",
          5080 => x"00",
          5081 => x"00",
          5082 => x"00",
          5083 => x"00",
          5084 => x"73",
          5085 => x"00",
          5086 => x"61",
          5087 => x"2e",
          5088 => x"6f",
          5089 => x"2e",
          5090 => x"65",
          5091 => x"00",
          5092 => x"68",
          5093 => x"00",
          5094 => x"64",
          5095 => x"6d",
          5096 => x"63",
          5097 => x"69",
          5098 => x"6c",
          5099 => x"64",
          5100 => x"73",
          5101 => x"6c",
          5102 => x"65",
          5103 => x"64",
          5104 => x"20",
          5105 => x"65",
          5106 => x"74",
          5107 => x"69",
          5108 => x"65",
          5109 => x"76",
          5110 => x"00",
          5111 => x"6f",
          5112 => x"65",
          5113 => x"20",
          5114 => x"62",
          5115 => x"73",
          5116 => x"6f",
          5117 => x"64",
          5118 => x"72",
          5119 => x"72",
          5120 => x"6d",
          5121 => x"70",
          5122 => x"20",
          5123 => x"65",
          5124 => x"6c",
          5125 => x"63",
          5126 => x"73",
          5127 => x"6e",
          5128 => x"79",
          5129 => x"6f",
          5130 => x"70",
          5131 => x"73",
          5132 => x"72",
          5133 => x"20",
          5134 => x"63",
          5135 => x"63",
          5136 => x"00",
          5137 => x"6e",
          5138 => x"00",
          5139 => x"79",
          5140 => x"61",
          5141 => x"79",
          5142 => x"2e",
          5143 => x"61",
          5144 => x"38",
          5145 => x"20",
          5146 => x"00",
          5147 => x"20",
          5148 => x"32",
          5149 => x"00",
          5150 => x"00",
          5151 => x"20",
          5152 => x"2f",
          5153 => x"00",
          5154 => x"00",
          5155 => x"72",
          5156 => x"29",
          5157 => x"2a",
          5158 => x"55",
          5159 => x"75",
          5160 => x"6c",
          5161 => x"6d",
          5162 => x"72",
          5163 => x"32",
          5164 => x"75",
          5165 => x"43",
          5166 => x"6e",
          5167 => x"00",
          5168 => x"57",
          5169 => x"72",
          5170 => x"52",
          5171 => x"6e",
          5172 => x"00",
          5173 => x"54",
          5174 => x"72",
          5175 => x"52",
          5176 => x"6e",
          5177 => x"00",
          5178 => x"54",
          5179 => x"72",
          5180 => x"74",
          5181 => x"20",
          5182 => x"2e",
          5183 => x"6e",
          5184 => x"2e",
          5185 => x"74",
          5186 => x"61",
          5187 => x"53",
          5188 => x"74",
          5189 => x"69",
          5190 => x"69",
          5191 => x"73",
          5192 => x"72",
          5193 => x"65",
          5194 => x"74",
          5195 => x"6c",
          5196 => x"00",
          5197 => x"6e",
          5198 => x"00",
          5199 => x"67",
          5200 => x"6d",
          5201 => x"2e",
          5202 => x"38",
          5203 => x"29",
          5204 => x"28",
          5205 => x"00",
          5206 => x"65",
          5207 => x"6f",
          5208 => x"00",
          5209 => x"25",
          5210 => x"3f",
          5211 => x"25",
          5212 => x"38",
          5213 => x"58",
          5214 => x"65",
          5215 => x"63",
          5216 => x"30",
          5217 => x"0a",
          5218 => x"67",
          5219 => x"20",
          5220 => x"2e",
          5221 => x"6c",
          5222 => x"6e",
          5223 => x"20",
          5224 => x"00",
          5225 => x"74",
          5226 => x"6c",
          5227 => x"2e",
          5228 => x"6c",
          5229 => x"74",
          5230 => x"00",
          5231 => x"6e",
          5232 => x"5c",
          5233 => x"00",
          5234 => x"5c",
          5235 => x"3a",
          5236 => x"64",
          5237 => x"64",
          5238 => x"6d",
          5239 => x"61",
          5240 => x"63",
          5241 => x"72",
          5242 => x"6f",
          5243 => x"00",
          5244 => x"67",
          5245 => x"61",
          5246 => x"6e",
          5247 => x"73",
          5248 => x"2f",
          5249 => x"64",
          5250 => x"25",
          5251 => x"43",
          5252 => x"75",
          5253 => x"00",
          5254 => x"20",
          5255 => x"66",
          5256 => x"44",
          5257 => x"69",
          5258 => x"74",
          5259 => x"20",
          5260 => x"41",
          5261 => x"58",
          5262 => x"0a",
          5263 => x"52",
          5264 => x"28",
          5265 => x"38",
          5266 => x"20",
          5267 => x"52",
          5268 => x"58",
          5269 => x"0a",
          5270 => x"41",
          5271 => x"28",
          5272 => x"38",
          5273 => x"20",
          5274 => x"20",
          5275 => x"58",
          5276 => x"0a",
          5277 => x"20",
          5278 => x"28",
          5279 => x"20",
          5280 => x"0a",
          5281 => x"4d",
          5282 => x"28",
          5283 => x"20",
          5284 => x"0a",
          5285 => x"54",
          5286 => x"28",
          5287 => x"73",
          5288 => x"0a",
          5289 => x"53",
          5290 => x"55",
          5291 => x"20",
          5292 => x"00",
          5293 => x"43",
          5294 => x"20",
          5295 => x"20",
          5296 => x"64",
          5297 => x"00",
          5298 => x"55",
          5299 => x"56",
          5300 => x"64",
          5301 => x"20",
          5302 => x"00",
          5303 => x"55",
          5304 => x"20",
          5305 => x"64",
          5306 => x"20",
          5307 => x"00",
          5308 => x"61",
          5309 => x"74",
          5310 => x"73",
          5311 => x"20",
          5312 => x"00",
          5313 => x"00",
          5314 => x"55",
          5315 => x"20",
          5316 => x"20",
          5317 => x"20",
          5318 => x"00",
          5319 => x"73",
          5320 => x"63",
          5321 => x"20",
          5322 => x"20",
          5323 => x"4d",
          5324 => x"20",
          5325 => x"43",
          5326 => x"65",
          5327 => x"20",
          5328 => x"25",
          5329 => x"00",
          5330 => x"73",
          5331 => x"44",
          5332 => x"63",
          5333 => x"20",
          5334 => x"4d",
          5335 => x"61",
          5336 => x"64",
          5337 => x"65",
          5338 => x"4f",
          5339 => x"00",
          5340 => x"6e",
          5341 => x"00",
          5342 => x"a8",
          5343 => x"00",
          5344 => x"00",
          5345 => x"a8",
          5346 => x"00",
          5347 => x"00",
          5348 => x"a8",
          5349 => x"00",
          5350 => x"00",
          5351 => x"a8",
          5352 => x"00",
          5353 => x"00",
          5354 => x"a8",
          5355 => x"00",
          5356 => x"00",
          5357 => x"a8",
          5358 => x"00",
          5359 => x"00",
          5360 => x"a8",
          5361 => x"00",
          5362 => x"00",
          5363 => x"a8",
          5364 => x"00",
          5365 => x"00",
          5366 => x"a8",
          5367 => x"00",
          5368 => x"00",
          5369 => x"a7",
          5370 => x"00",
          5371 => x"00",
          5372 => x"a7",
          5373 => x"00",
          5374 => x"43",
          5375 => x"41",
          5376 => x"35",
          5377 => x"46",
          5378 => x"32",
          5379 => x"00",
          5380 => x"00",
          5381 => x"00",
          5382 => x"00",
          5383 => x"00",
          5384 => x"00",
          5385 => x"79",
          5386 => x"00",
          5387 => x"34",
          5388 => x"00",
          5389 => x"20",
          5390 => x"74",
          5391 => x"73",
          5392 => x"6c",
          5393 => x"46",
          5394 => x"6e",
          5395 => x"6e",
          5396 => x"20",
          5397 => x"20",
          5398 => x"69",
          5399 => x"2e",
          5400 => x"3a",
          5401 => x"00",
          5402 => x"00",
          5403 => x"54",
          5404 => x"90",
          5405 => x"30",
          5406 => x"45",
          5407 => x"33",
          5408 => x"20",
          5409 => x"20",
          5410 => x"20",
          5411 => x"00",
          5412 => x"00",
          5413 => x"10",
          5414 => x"00",
          5415 => x"8f",
          5416 => x"8e",
          5417 => x"55",
          5418 => x"9e",
          5419 => x"a6",
          5420 => x"ae",
          5421 => x"b6",
          5422 => x"be",
          5423 => x"c6",
          5424 => x"ce",
          5425 => x"d6",
          5426 => x"de",
          5427 => x"e6",
          5428 => x"ee",
          5429 => x"f6",
          5430 => x"fe",
          5431 => x"5d",
          5432 => x"3f",
          5433 => x"00",
          5434 => x"02",
          5435 => x"00",
          5436 => x"00",
          5437 => x"00",
          5438 => x"00",
          5439 => x"00",
          5440 => x"00",
          5441 => x"00",
          5442 => x"00",
          5443 => x"00",
          5444 => x"00",
          5445 => x"00",
          5446 => x"00",
          5447 => x"23",
          5448 => x"00",
          5449 => x"25",
          5450 => x"25",
          5451 => x"25",
          5452 => x"25",
          5453 => x"25",
          5454 => x"25",
          5455 => x"25",
          5456 => x"25",
          5457 => x"25",
          5458 => x"25",
          5459 => x"25",
          5460 => x"25",
          5461 => x"00",
          5462 => x"03",
          5463 => x"03",
          5464 => x"03",
          5465 => x"00",
          5466 => x"23",
          5467 => x"22",
          5468 => x"00",
          5469 => x"03",
          5470 => x"03",
          5471 => x"01",
          5472 => x"01",
          5473 => x"01",
          5474 => x"02",
          5475 => x"01",
          5476 => x"01",
          5477 => x"01",
          5478 => x"01",
          5479 => x"01",
          5480 => x"01",
          5481 => x"01",
          5482 => x"01",
          5483 => x"01",
          5484 => x"01",
          5485 => x"01",
          5486 => x"01",
          5487 => x"01",
          5488 => x"01",
          5489 => x"01",
          5490 => x"01",
          5491 => x"01",
          5492 => x"01",
          5493 => x"01",
          5494 => x"00",
          5495 => x"01",
          5496 => x"01",
          5497 => x"01",
          5498 => x"02",
          5499 => x"02",
          5500 => x"02",
          5501 => x"01",
          5502 => x"01",
          5503 => x"01",
          5504 => x"02",
          5505 => x"01",
          5506 => x"02",
          5507 => x"2c",
          5508 => x"01",
          5509 => x"02",
          5510 => x"02",
          5511 => x"02",
          5512 => x"02",
          5513 => x"01",
          5514 => x"02",
          5515 => x"01",
          5516 => x"02",
          5517 => x"03",
          5518 => x"03",
          5519 => x"03",
          5520 => x"03",
          5521 => x"03",
          5522 => x"00",
          5523 => x"03",
          5524 => x"03",
          5525 => x"03",
          5526 => x"03",
          5527 => x"04",
          5528 => x"04",
          5529 => x"04",
          5530 => x"01",
          5531 => x"00",
          5532 => x"1e",
          5533 => x"1f",
          5534 => x"1f",
          5535 => x"1f",
          5536 => x"1f",
          5537 => x"1f",
          5538 => x"06",
          5539 => x"1f",
          5540 => x"1f",
          5541 => x"1f",
          5542 => x"1f",
          5543 => x"06",
          5544 => x"00",
          5545 => x"1f",
          5546 => x"1f",
          5547 => x"1f",
          5548 => x"00",
          5549 => x"21",
          5550 => x"00",
          5551 => x"2c",
          5552 => x"2c",
          5553 => x"2c",
          5554 => x"ff",
          5555 => x"00",
          5556 => x"01",
          5557 => x"00",
          5558 => x"01",
          5559 => x"00",
          5560 => x"03",
          5561 => x"00",
          5562 => x"03",
          5563 => x"00",
          5564 => x"03",
          5565 => x"00",
          5566 => x"04",
          5567 => x"00",
          5568 => x"04",
          5569 => x"00",
          5570 => x"04",
          5571 => x"00",
          5572 => x"04",
          5573 => x"00",
          5574 => x"04",
          5575 => x"00",
          5576 => x"04",
          5577 => x"00",
          5578 => x"04",
          5579 => x"00",
          5580 => x"05",
          5581 => x"00",
          5582 => x"05",
          5583 => x"00",
          5584 => x"05",
          5585 => x"00",
          5586 => x"05",
          5587 => x"00",
          5588 => x"07",
          5589 => x"00",
          5590 => x"07",
          5591 => x"00",
          5592 => x"08",
          5593 => x"00",
          5594 => x"08",
          5595 => x"00",
          5596 => x"08",
          5597 => x"00",
          5598 => x"09",
          5599 => x"00",
          5600 => x"09",
          5601 => x"00",
          5602 => x"09",
          5603 => x"00",
          5604 => x"09",
          5605 => x"00",
          5606 => x"00",
          5607 => x"00",
          5608 => x"00",
          5609 => x"00",
          5610 => x"00",
          5611 => x"00",
          5612 => x"78",
          5613 => x"e1",
          5614 => x"e1",
          5615 => x"01",
          5616 => x"10",
          5617 => x"00",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"a8",
          5630 => x"a8",
          5631 => x"a8",
          5632 => x"00",
          5633 => x"00",
          5634 => x"00",
        others => X"00"
    );

    shared variable RAM6 : ramArray :=
    (
             0 => x"0d",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"08",
             5 => x"0c",
             6 => x"00",
             7 => x"00",
             8 => x"83",
             9 => x"2b",
            10 => x"00",
            11 => x"00",
            12 => x"ff",
            13 => x"82",
            14 => x"83",
            15 => x"a5",
            16 => x"05",
            17 => x"09",
            18 => x"51",
            19 => x"00",
            20 => x"2e",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"10",
            26 => x"0a",
            27 => x"00",
            28 => x"2e",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"04",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"53",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"81",
            45 => x"04",
            46 => x"00",
            47 => x"00",
            48 => x"9f",
            49 => x"06",
            50 => x"00",
            51 => x"00",
            52 => x"06",
            53 => x"05",
            54 => x"06",
            55 => x"00",
            56 => x"05",
            57 => x"81",
            58 => x"00",
            59 => x"00",
            60 => x"05",
            61 => x"09",
            62 => x"00",
            63 => x"00",
            64 => x"04",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"83",
            77 => x"10",
            78 => x"00",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"b9",
            83 => x"00",
            84 => x"08",
            85 => x"2d",
            86 => x"8c",
            87 => x"00",
            88 => x"08",
            89 => x"2d",
            90 => x"8c",
            91 => x"00",
            92 => x"09",
            93 => x"54",
            94 => x"ff",
            95 => x"00",
            96 => x"09",
            97 => x"70",
            98 => x"05",
            99 => x"04",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"71",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"04",
           133 => x"0b",
           134 => x"8c",
           135 => x"04",
           136 => x"0b",
           137 => x"8c",
           138 => x"04",
           139 => x"0b",
           140 => x"8d",
           141 => x"04",
           142 => x"0b",
           143 => x"8d",
           144 => x"04",
           145 => x"0b",
           146 => x"8e",
           147 => x"04",
           148 => x"0b",
           149 => x"8e",
           150 => x"04",
           151 => x"0b",
           152 => x"8f",
           153 => x"04",
           154 => x"0b",
           155 => x"8f",
           156 => x"04",
           157 => x"0b",
           158 => x"90",
           159 => x"04",
           160 => x"0b",
           161 => x"91",
           162 => x"04",
           163 => x"0b",
           164 => x"91",
           165 => x"04",
           166 => x"0b",
           167 => x"92",
           168 => x"04",
           169 => x"0b",
           170 => x"92",
           171 => x"04",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"82",
           193 => x"82",
           194 => x"04",
           195 => x"82",
           196 => x"04",
           197 => x"82",
           198 => x"04",
           199 => x"82",
           200 => x"04",
           201 => x"82",
           202 => x"04",
           203 => x"82",
           204 => x"04",
           205 => x"2d",
           206 => x"90",
           207 => x"ce",
           208 => x"80",
           209 => x"8c",
           210 => x"80",
           211 => x"f4",
           212 => x"80",
           213 => x"81",
           214 => x"80",
           215 => x"e0",
           216 => x"c0",
           217 => x"80",
           218 => x"80",
           219 => x"0c",
           220 => x"08",
           221 => x"a4",
           222 => x"a4",
           223 => x"e0",
           224 => x"e0",
           225 => x"82",
           226 => x"82",
           227 => x"04",
           228 => x"2d",
           229 => x"90",
           230 => x"8c",
           231 => x"80",
           232 => x"fe",
           233 => x"c0",
           234 => x"82",
           235 => x"80",
           236 => x"0c",
           237 => x"08",
           238 => x"a4",
           239 => x"a4",
           240 => x"e0",
           241 => x"e0",
           242 => x"82",
           243 => x"82",
           244 => x"04",
           245 => x"2d",
           246 => x"90",
           247 => x"bb",
           248 => x"80",
           249 => x"93",
           250 => x"c0",
           251 => x"82",
           252 => x"80",
           253 => x"0c",
           254 => x"08",
           255 => x"a4",
           256 => x"a4",
           257 => x"e0",
           258 => x"e0",
           259 => x"82",
           260 => x"82",
           261 => x"04",
           262 => x"2d",
           263 => x"90",
           264 => x"8b",
           265 => x"80",
           266 => x"8f",
           267 => x"c0",
           268 => x"82",
           269 => x"80",
           270 => x"0c",
           271 => x"08",
           272 => x"a4",
           273 => x"a4",
           274 => x"e0",
           275 => x"e0",
           276 => x"82",
           277 => x"82",
           278 => x"04",
           279 => x"2d",
           280 => x"90",
           281 => x"d5",
           282 => x"80",
           283 => x"b5",
           284 => x"c0",
           285 => x"81",
           286 => x"80",
           287 => x"0c",
           288 => x"08",
           289 => x"a4",
           290 => x"a4",
           291 => x"e0",
           292 => x"e0",
           293 => x"82",
           294 => x"82",
           295 => x"04",
           296 => x"2d",
           297 => x"90",
           298 => x"9f",
           299 => x"80",
           300 => x"af",
           301 => x"c0",
           302 => x"81",
           303 => x"80",
           304 => x"0c",
           305 => x"08",
           306 => x"10",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"51",
           311 => x"73",
           312 => x"10",
           313 => x"0c",
           314 => x"81",
           315 => x"71",
           316 => x"72",
           317 => x"82",
           318 => x"8e",
           319 => x"0c",
           320 => x"81",
           321 => x"e0",
           322 => x"fb",
           323 => x"05",
           324 => x"0c",
           325 => x"54",
           326 => x"53",
           327 => x"9a",
           328 => x"e0",
           329 => x"a4",
           330 => x"98",
           331 => x"e0",
           332 => x"02",
           333 => x"82",
           334 => x"11",
           335 => x"51",
           336 => x"0b",
           337 => x"25",
           338 => x"e0",
           339 => x"39",
           340 => x"ff",
           341 => x"0c",
           342 => x"05",
           343 => x"08",
           344 => x"82",
           345 => x"2e",
           346 => x"a4",
           347 => x"38",
           348 => x"51",
           349 => x"70",
           350 => x"52",
           351 => x"ff",
           352 => x"0b",
           353 => x"80",
           354 => x"05",
           355 => x"08",
           356 => x"a4",
           357 => x"e0",
           358 => x"a4",
           359 => x"e0",
           360 => x"39",
           361 => x"52",
           362 => x"88",
           363 => x"f4",
           364 => x"f4",
           365 => x"3d",
           366 => x"e0",
           367 => x"f4",
           368 => x"08",
           369 => x"88",
           370 => x"05",
           371 => x"08",
           372 => x"90",
           373 => x"05",
           374 => x"08",
           375 => x"08",
           376 => x"70",
           377 => x"e0",
           378 => x"dc",
           379 => x"05",
           380 => x"08",
           381 => x"e0",
           382 => x"e0",
           383 => x"e0",
           384 => x"02",
           385 => x"82",
           386 => x"e0",
           387 => x"a4",
           388 => x"a4",
           389 => x"a4",
           390 => x"3f",
           391 => x"a4",
           392 => x"08",
           393 => x"0c",
           394 => x"a4",
           395 => x"82",
           396 => x"0b",
           397 => x"82",
           398 => x"80",
           399 => x"08",
           400 => x"81",
           401 => x"51",
           402 => x"8d",
           403 => x"e0",
           404 => x"a4",
           405 => x"53",
           406 => x"34",
           407 => x"2e",
           408 => x"8c",
           409 => x"08",
           410 => x"e4",
           411 => x"72",
           412 => x"a4",
           413 => x"27",
           414 => x"f8",
           415 => x"ee",
           416 => x"33",
           417 => x"80",
           418 => x"05",
           419 => x"51",
           420 => x"a4",
           421 => x"70",
           422 => x"51",
           423 => x"e0",
           424 => x"80",
           425 => x"08",
           426 => x"e0",
           427 => x"2b",
           428 => x"72",
           429 => x"51",
           430 => x"e8",
           431 => x"05",
           432 => x"05",
           433 => x"53",
           434 => x"34",
           435 => x"70",
           436 => x"53",
           437 => x"0b",
           438 => x"82",
           439 => x"83",
           440 => x"72",
           441 => x"e8",
           442 => x"2b",
           443 => x"51",
           444 => x"08",
           445 => x"e0",
           446 => x"2a",
           447 => x"80",
           448 => x"e8",
           449 => x"2c",
           450 => x"0b",
           451 => x"82",
           452 => x"11",
           453 => x"53",
           454 => x"80",
           455 => x"a4",
           456 => x"82",
           457 => x"51",
           458 => x"e4",
           459 => x"72",
           460 => x"82",
           461 => x"a0",
           462 => x"08",
           463 => x"e0",
           464 => x"80",
           465 => x"08",
           466 => x"e0",
           467 => x"c0",
           468 => x"08",
           469 => x"e0",
           470 => x"07",
           471 => x"e4",
           472 => x"08",
           473 => x"e0",
           474 => x"07",
           475 => x"e4",
           476 => x"82",
           477 => x"e0",
           478 => x"51",
           479 => x"05",
           480 => x"08",
           481 => x"e0",
           482 => x"a4",
           483 => x"e0",
           484 => x"51",
           485 => x"05",
           486 => x"22",
           487 => x"a4",
           488 => x"82",
           489 => x"e0",
           490 => x"82",
           491 => x"08",
           492 => x"82",
           493 => x"83",
           494 => x"53",
           495 => x"a4",
           496 => x"53",
           497 => x"08",
           498 => x"3f",
           499 => x"e0",
           500 => x"82",
           501 => x"9d",
           502 => x"72",
           503 => x"82",
           504 => x"82",
           505 => x"71",
           506 => x"08",
           507 => x"e0",
           508 => x"a4",
           509 => x"e0",
           510 => x"82",
           511 => x"e0",
           512 => x"2a",
           513 => x"72",
           514 => x"08",
           515 => x"72",
           516 => x"fc",
           517 => x"82",
           518 => x"a4",
           519 => x"e0",
           520 => x"f3",
           521 => x"82",
           522 => x"e0",
           523 => x"e0",
           524 => x"31",
           525 => x"ec",
           526 => x"a4",
           527 => x"70",
           528 => x"2e",
           529 => x"05",
           530 => x"08",
           531 => x"05",
           532 => x"dc",
           533 => x"a4",
           534 => x"08",
           535 => x"a4",
           536 => x"e0",
           537 => x"e0",
           538 => x"a4",
           539 => x"08",
           540 => x"82",
           541 => x"82",
           542 => x"08",
           543 => x"fc",
           544 => x"fc",
           545 => x"05",
           546 => x"72",
           547 => x"81",
           548 => x"08",
           549 => x"a4",
           550 => x"07",
           551 => x"e4",
           552 => x"a4",
           553 => x"e0",
           554 => x"a4",
           555 => x"70",
           556 => x"2e",
           557 => x"05",
           558 => x"08",
           559 => x"05",
           560 => x"d8",
           561 => x"a4",
           562 => x"08",
           563 => x"a4",
           564 => x"e0",
           565 => x"e0",
           566 => x"a4",
           567 => x"08",
           568 => x"53",
           569 => x"23",
           570 => x"08",
           571 => x"f0",
           572 => x"05",
           573 => x"08",
           574 => x"aa",
           575 => x"72",
           576 => x"05",
           577 => x"0c",
           578 => x"70",
           579 => x"38",
           580 => x"53",
           581 => x"f8",
           582 => x"51",
           583 => x"05",
           584 => x"f0",
           585 => x"51",
           586 => x"05",
           587 => x"08",
           588 => x"33",
           589 => x"05",
           590 => x"f0",
           591 => x"05",
           592 => x"fc",
           593 => x"82",
           594 => x"08",
           595 => x"08",
           596 => x"fe",
           597 => x"05",
           598 => x"54",
           599 => x"82",
           600 => x"e0",
           601 => x"06",
           602 => x"82",
           603 => x"11",
           604 => x"ec",
           605 => x"05",
           606 => x"51",
           607 => x"38",
           608 => x"70",
           609 => x"05",
           610 => x"08",
           611 => x"05",
           612 => x"22",
           613 => x"06",
           614 => x"05",
           615 => x"a4",
           616 => x"e0",
           617 => x"53",
           618 => x"23",
           619 => x"82",
           620 => x"e0",
           621 => x"2a",
           622 => x"80",
           623 => x"08",
           624 => x"98",
           625 => x"33",
           626 => x"97",
           627 => x"22",
           628 => x"e0",
           629 => x"82",
           630 => x"82",
           631 => x"71",
           632 => x"08",
           633 => x"e4",
           634 => x"06",
           635 => x"38",
           636 => x"70",
           637 => x"2c",
           638 => x"53",
           639 => x"05",
           640 => x"82",
           641 => x"39",
           642 => x"70",
           643 => x"2c",
           644 => x"53",
           645 => x"05",
           646 => x"82",
           647 => x"e0",
           648 => x"80",
           649 => x"e0",
           650 => x"54",
           651 => x"05",
           652 => x"51",
           653 => x"e0",
           654 => x"51",
           655 => x"a4",
           656 => x"70",
           657 => x"2e",
           658 => x"05",
           659 => x"80",
           660 => x"05",
           661 => x"51",
           662 => x"82",
           663 => x"ab",
           664 => x"e0",
           665 => x"2a",
           666 => x"80",
           667 => x"88",
           668 => x"3f",
           669 => x"70",
           670 => x"53",
           671 => x"a4",
           672 => x"89",
           673 => x"05",
           674 => x"06",
           675 => x"05",
           676 => x"05",
           677 => x"a4",
           678 => x"70",
           679 => x"2e",
           680 => x"05",
           681 => x"e0",
           682 => x"2b",
           683 => x"25",
           684 => x"05",
           685 => x"d2",
           686 => x"22",
           687 => x"51",
           688 => x"e0",
           689 => x"54",
           690 => x"05",
           691 => x"51",
           692 => x"e0",
           693 => x"51",
           694 => x"a4",
           695 => x"70",
           696 => x"38",
           697 => x"ff",
           698 => x"08",
           699 => x"90",
           700 => x"38",
           701 => x"52",
           702 => x"82",
           703 => x"72",
           704 => x"38",
           705 => x"52",
           706 => x"51",
           707 => x"e0",
           708 => x"80",
           709 => x"38",
           710 => x"ff",
           711 => x"08",
           712 => x"06",
           713 => x"bb",
           714 => x"08",
           715 => x"08",
           716 => x"fc",
           717 => x"08",
           718 => x"ff",
           719 => x"05",
           720 => x"81",
           721 => x"08",
           722 => x"72",
           723 => x"72",
           724 => x"ff",
           725 => x"a4",
           726 => x"a4",
           727 => x"53",
           728 => x"fc",
           729 => x"08",
           730 => x"e0",
           731 => x"a8",
           732 => x"88",
           733 => x"f0",
           734 => x"08",
           735 => x"f0",
           736 => x"e0",
           737 => x"e4",
           738 => x"06",
           739 => x"c3",
           740 => x"22",
           741 => x"a4",
           742 => x"70",
           743 => x"a3",
           744 => x"08",
           745 => x"39",
           746 => x"52",
           747 => x"51",
           748 => x"a4",
           749 => x"82",
           750 => x"72",
           751 => x"81",
           752 => x"23",
           753 => x"05",
           754 => x"e8",
           755 => x"08",
           756 => x"e0",
           757 => x"e0",
           758 => x"b0",
           759 => x"08",
           760 => x"82",
           761 => x"53",
           762 => x"82",
           763 => x"e0",
           764 => x"02",
           765 => x"82",
           766 => x"08",
           767 => x"08",
           768 => x"82",
           769 => x"0c",
           770 => x"0c",
           771 => x"e0",
           772 => x"82",
           773 => x"fb",
           774 => x"2a",
           775 => x"51",
           776 => x"38",
           777 => x"05",
           778 => x"08",
           779 => x"e0",
           780 => x"82",
           781 => x"72",
           782 => x"72",
           783 => x"b0",
           784 => x"fc",
           785 => x"05",
           786 => x"72",
           787 => x"80",
           788 => x"e0",
           789 => x"39",
           790 => x"08",
           791 => x"53",
           792 => x"72",
           793 => x"e0",
           794 => x"a4",
           795 => x"a4",
           796 => x"a4",
           797 => x"0c",
           798 => x"04",
           799 => x"a4",
           800 => x"e0",
           801 => x"a4",
           802 => x"70",
           803 => x"06",
           804 => x"2e",
           805 => x"08",
           806 => x"e0",
           807 => x"33",
           808 => x"81",
           809 => x"0c",
           810 => x"05",
           811 => x"80",
           812 => x"8c",
           813 => x"05",
           814 => x"05",
           815 => x"72",
           816 => x"80",
           817 => x"e0",
           818 => x"39",
           819 => x"70",
           820 => x"53",
           821 => x"82",
           822 => x"e0",
           823 => x"02",
           824 => x"82",
           825 => x"08",
           826 => x"e0",
           827 => x"53",
           828 => x"04",
           829 => x"a4",
           830 => x"08",
           831 => x"81",
           832 => x"51",
           833 => x"8d",
           834 => x"fc",
           835 => x"a4",
           836 => x"70",
           837 => x"51",
           838 => x"82",
           839 => x"e0",
           840 => x"8c",
           841 => x"38",
           842 => x"70",
           843 => x"05",
           844 => x"34",
           845 => x"e0",
           846 => x"08",
           847 => x"a4",
           848 => x"a4",
           849 => x"d7",
           850 => x"08",
           851 => x"53",
           852 => x"70",
           853 => x"51",
           854 => x"08",
           855 => x"08",
           856 => x"05",
           857 => x"88",
           858 => x"fc",
           859 => x"0b",
           860 => x"82",
           861 => x"e0",
           862 => x"a4",
           863 => x"82",
           864 => x"e0",
           865 => x"33",
           866 => x"51",
           867 => x"ff",
           868 => x"0c",
           869 => x"88",
           870 => x"2a",
           871 => x"71",
           872 => x"a4",
           873 => x"08",
           874 => x"33",
           875 => x"85",
           876 => x"05",
           877 => x"12",
           878 => x"08",
           879 => x"08",
           880 => x"b6",
           881 => x"08",
           882 => x"81",
           883 => x"2e",
           884 => x"88",
           885 => x"e0",
           886 => x"82",
           887 => x"38",
           888 => x"82",
           889 => x"53",
           890 => x"52",
           891 => x"e0",
           892 => x"39",
           893 => x"70",
           894 => x"a1",
           895 => x"08",
           896 => x"52",
           897 => x"82",
           898 => x"08",
           899 => x"08",
           900 => x"38",
           901 => x"82",
           902 => x"e0",
           903 => x"33",
           904 => x"52",
           905 => x"ff",
           906 => x"e0",
           907 => x"52",
           908 => x"34",
           909 => x"05",
           910 => x"a4",
           911 => x"08",
           912 => x"08",
           913 => x"0b",
           914 => x"a6",
           915 => x"08",
           916 => x"0c",
           917 => x"70",
           918 => x"08",
           919 => x"e0",
           920 => x"98",
           921 => x"0c",
           922 => x"e0",
           923 => x"a4",
           924 => x"08",
           925 => x"8c",
           926 => x"05",
           927 => x"08",
           928 => x"a4",
           929 => x"08",
           930 => x"82",
           931 => x"e0",
           932 => x"82",
           933 => x"27",
           934 => x"fc",
           935 => x"05",
           936 => x"05",
           937 => x"08",
           938 => x"05",
           939 => x"82",
           940 => x"05",
           941 => x"82",
           942 => x"05",
           943 => x"82",
           944 => x"2e",
           945 => x"fc",
           946 => x"08",
           947 => x"f8",
           948 => x"08",
           949 => x"fc",
           950 => x"05",
           951 => x"ff",
           952 => x"05",
           953 => x"90",
           954 => x"05",
           955 => x"90",
           956 => x"05",
           957 => x"a4",
           958 => x"82",
           959 => x"05",
           960 => x"82",
           961 => x"52",
           962 => x"fc",
           963 => x"08",
           964 => x"e0",
           965 => x"e0",
           966 => x"e0",
           967 => x"02",
           968 => x"82",
           969 => x"e0",
           970 => x"a4",
           971 => x"82",
           972 => x"05",
           973 => x"70",
           974 => x"2e",
           975 => x"08",
           976 => x"a4",
           977 => x"08",
           978 => x"88",
           979 => x"0c",
           980 => x"0c",
           981 => x"e0",
           982 => x"a4",
           983 => x"08",
           984 => x"8c",
           985 => x"a4",
           986 => x"e0",
           987 => x"a4",
           988 => x"72",
           989 => x"08",
           990 => x"05",
           991 => x"80",
           992 => x"e0",
           993 => x"e0",
           994 => x"e0",
           995 => x"02",
           996 => x"82",
           997 => x"e0",
           998 => x"a4",
           999 => x"08",
          1000 => x"90",
          1001 => x"82",
          1002 => x"05",
          1003 => x"82",
          1004 => x"05",
          1005 => x"82",
          1006 => x"2e",
          1007 => x"05",
          1008 => x"08",
          1009 => x"a4",
          1010 => x"08",
          1011 => x"34",
          1012 => x"81",
          1013 => x"0c",
          1014 => x"88",
          1015 => x"51",
          1016 => x"04",
          1017 => x"a4",
          1018 => x"08",
          1019 => x"38",
          1020 => x"52",
          1021 => x"05",
          1022 => x"8c",
          1023 => x"05",
          1024 => x"53",
          1025 => x"38",
          1026 => x"88",
          1027 => x"a4",
          1028 => x"e0",
          1029 => x"ff",
          1030 => x"0b",
          1031 => x"81",
          1032 => x"05",
          1033 => x"90",
          1034 => x"05",
          1035 => x"39",
          1036 => x"80",
          1037 => x"08",
          1038 => x"70",
          1039 => x"08",
          1040 => x"e0",
          1041 => x"82",
          1042 => x"e0",
          1043 => x"52",
          1044 => x"e0",
          1045 => x"82",
          1046 => x"33",
          1047 => x"70",
          1048 => x"a4",
          1049 => x"52",
          1050 => x"a4",
          1051 => x"08",
          1052 => x"85",
          1053 => x"82",
          1054 => x"0c",
          1055 => x"8c",
          1056 => x"88",
          1057 => x"e0",
          1058 => x"f8",
          1059 => x"05",
          1060 => x"80",
          1061 => x"70",
          1062 => x"54",
          1063 => x"8c",
          1064 => x"f4",
          1065 => x"08",
          1066 => x"f8",
          1067 => x"82",
          1068 => x"82",
          1069 => x"82",
          1070 => x"fb",
          1071 => x"82",
          1072 => x"82",
          1073 => x"e0",
          1074 => x"a4",
          1075 => x"82",
          1076 => x"e0",
          1077 => x"a4",
          1078 => x"08",
          1079 => x"82",
          1080 => x"ec",
          1081 => x"08",
          1082 => x"f8",
          1083 => x"08",
          1084 => x"51",
          1085 => x"e0",
          1086 => x"82",
          1087 => x"e0",
          1088 => x"84",
          1089 => x"08",
          1090 => x"a4",
          1091 => x"08",
          1092 => x"88",
          1093 => x"08",
          1094 => x"08",
          1095 => x"85",
          1096 => x"82",
          1097 => x"0c",
          1098 => x"88",
          1099 => x"05",
          1100 => x"08",
          1101 => x"a4",
          1102 => x"e0",
          1103 => x"a4",
          1104 => x"e0",
          1105 => x"a4",
          1106 => x"38",
          1107 => x"51",
          1108 => x"08",
          1109 => x"a4",
          1110 => x"e0",
          1111 => x"39",
          1112 => x"70",
          1113 => x"0d",
          1114 => x"a4",
          1115 => x"3d",
          1116 => x"08",
          1117 => x"08",
          1118 => x"70",
          1119 => x"0d",
          1120 => x"a4",
          1121 => x"3d",
          1122 => x"fc",
          1123 => x"05",
          1124 => x"a4",
          1125 => x"3f",
          1126 => x"a4",
          1127 => x"82",
          1128 => x"e0",
          1129 => x"a4",
          1130 => x"38",
          1131 => x"51",
          1132 => x"82",
          1133 => x"31",
          1134 => x"52",
          1135 => x"05",
          1136 => x"08",
          1137 => x"0c",
          1138 => x"82",
          1139 => x"e0",
          1140 => x"52",
          1141 => x"08",
          1142 => x"a4",
          1143 => x"82",
          1144 => x"05",
          1145 => x"05",
          1146 => x"82",
          1147 => x"82",
          1148 => x"82",
          1149 => x"05",
          1150 => x"f8",
          1151 => x"05",
          1152 => x"08",
          1153 => x"0c",
          1154 => x"82",
          1155 => x"82",
          1156 => x"2b",
          1157 => x"52",
          1158 => x"05",
          1159 => x"08",
          1160 => x"a4",
          1161 => x"a4",
          1162 => x"e0",
          1163 => x"70",
          1164 => x"05",
          1165 => x"08",
          1166 => x"05",
          1167 => x"05",
          1168 => x"08",
          1169 => x"31",
          1170 => x"05",
          1171 => x"e0",
          1172 => x"a4",
          1173 => x"e0",
          1174 => x"a4",
          1175 => x"08",
          1176 => x"08",
          1177 => x"a4",
          1178 => x"08",
          1179 => x"a4",
          1180 => x"51",
          1181 => x"82",
          1182 => x"70",
          1183 => x"07",
          1184 => x"82",
          1185 => x"82",
          1186 => x"52",
          1187 => x"82",
          1188 => x"e0",
          1189 => x"02",
          1190 => x"82",
          1191 => x"e0",
          1192 => x"a4",
          1193 => x"06",
          1194 => x"e0",
          1195 => x"80",
          1196 => x"0c",
          1197 => x"82",
          1198 => x"0b",
          1199 => x"31",
          1200 => x"71",
          1201 => x"0c",
          1202 => x"82",
          1203 => x"e0",
          1204 => x"80",
          1205 => x"0b",
          1206 => x"8a",
          1207 => x"ec",
          1208 => x"05",
          1209 => x"0c",
          1210 => x"05",
          1211 => x"05",
          1212 => x"fc",
          1213 => x"05",
          1214 => x"08",
          1215 => x"0c",
          1216 => x"81",
          1217 => x"84",
          1218 => x"0c",
          1219 => x"08",
          1220 => x"e8",
          1221 => x"05",
          1222 => x"f8",
          1223 => x"fc",
          1224 => x"08",
          1225 => x"f4",
          1226 => x"05",
          1227 => x"05",
          1228 => x"08",
          1229 => x"82",
          1230 => x"0c",
          1231 => x"08",
          1232 => x"e4",
          1233 => x"05",
          1234 => x"f8",
          1235 => x"fc",
          1236 => x"08",
          1237 => x"f4",
          1238 => x"05",
          1239 => x"05",
          1240 => x"fc",
          1241 => x"fc",
          1242 => x"70",
          1243 => x"82",
          1244 => x"70",
          1245 => x"55",
          1246 => x"3d",
          1247 => x"e0",
          1248 => x"fe",
          1249 => x"05",
          1250 => x"05",
          1251 => x"98",
          1252 => x"05",
          1253 => x"05",
          1254 => x"0c",
          1255 => x"e0",
          1256 => x"02",
          1257 => x"82",
          1258 => x"82",
          1259 => x"93",
          1260 => x"e0",
          1261 => x"e0",
          1262 => x"02",
          1263 => x"a0",
          1264 => x"0c",
          1265 => x"80",
          1266 => x"8c",
          1267 => x"e0",
          1268 => x"e4",
          1269 => x"a4",
          1270 => x"08",
          1271 => x"88",
          1272 => x"e0",
          1273 => x"db",
          1274 => x"a4",
          1275 => x"e0",
          1276 => x"39",
          1277 => x"82",
          1278 => x"82",
          1279 => x"e0",
          1280 => x"a4",
          1281 => x"08",
          1282 => x"82",
          1283 => x"94",
          1284 => x"08",
          1285 => x"0c",
          1286 => x"08",
          1287 => x"82",
          1288 => x"09",
          1289 => x"e0",
          1290 => x"39",
          1291 => x"81",
          1292 => x"0c",
          1293 => x"82",
          1294 => x"82",
          1295 => x"e0",
          1296 => x"a4",
          1297 => x"a4",
          1298 => x"e0",
          1299 => x"0b",
          1300 => x"82",
          1301 => x"2e",
          1302 => x"f4",
          1303 => x"fc",
          1304 => x"08",
          1305 => x"07",
          1306 => x"82",
          1307 => x"70",
          1308 => x"07",
          1309 => x"82",
          1310 => x"e0",
          1311 => x"11",
          1312 => x"ff",
          1313 => x"08",
          1314 => x"ec",
          1315 => x"08",
          1316 => x"8c",
          1317 => x"05",
          1318 => x"05",
          1319 => x"f4",
          1320 => x"05",
          1321 => x"f8",
          1322 => x"51",
          1323 => x"a4",
          1324 => x"a4",
          1325 => x"a4",
          1326 => x"0c",
          1327 => x"04",
          1328 => x"a4",
          1329 => x"e0",
          1330 => x"a4",
          1331 => x"08",
          1332 => x"08",
          1333 => x"8c",
          1334 => x"05",
          1335 => x"05",
          1336 => x"08",
          1337 => x"32",
          1338 => x"08",
          1339 => x"0c",
          1340 => x"82",
          1341 => x"70",
          1342 => x"31",
          1343 => x"82",
          1344 => x"e0",
          1345 => x"e0",
          1346 => x"a4",
          1347 => x"a4",
          1348 => x"f1",
          1349 => x"82",
          1350 => x"70",
          1351 => x"31",
          1352 => x"53",
          1353 => x"04",
          1354 => x"a4",
          1355 => x"e0",
          1356 => x"a4",
          1357 => x"0c",
          1358 => x"70",
          1359 => x"82",
          1360 => x"81",
          1361 => x"81",
          1362 => x"88",
          1363 => x"0c",
          1364 => x"f8",
          1365 => x"81",
          1366 => x"a4",
          1367 => x"08",
          1368 => x"71",
          1369 => x"82",
          1370 => x"e0",
          1371 => x"b0",
          1372 => x"82",
          1373 => x"08",
          1374 => x"53",
          1375 => x"05",
          1376 => x"33",
          1377 => x"82",
          1378 => x"e2",
          1379 => x"e8",
          1380 => x"80",
          1381 => x"08",
          1382 => x"88",
          1383 => x"0c",
          1384 => x"e0",
          1385 => x"39",
          1386 => x"05",
          1387 => x"08",
          1388 => x"08",
          1389 => x"08",
          1390 => x"e0",
          1391 => x"a0",
          1392 => x"a4",
          1393 => x"82",
          1394 => x"af",
          1395 => x"08",
          1396 => x"83",
          1397 => x"a4",
          1398 => x"88",
          1399 => x"34",
          1400 => x"05",
          1401 => x"82",
          1402 => x"72",
          1403 => x"0b",
          1404 => x"82",
          1405 => x"08",
          1406 => x"a4",
          1407 => x"08",
          1408 => x"81",
          1409 => x"05",
          1410 => x"38",
          1411 => x"e0",
          1412 => x"08",
          1413 => x"f8",
          1414 => x"82",
          1415 => x"e0",
          1416 => x"73",
          1417 => x"f8",
          1418 => x"82",
          1419 => x"e0",
          1420 => x"89",
          1421 => x"a4",
          1422 => x"82",
          1423 => x"e0",
          1424 => x"72",
          1425 => x"e0",
          1426 => x"39",
          1427 => x"70",
          1428 => x"29",
          1429 => x"70",
          1430 => x"0c",
          1431 => x"70",
          1432 => x"51",
          1433 => x"e0",
          1434 => x"39",
          1435 => x"53",
          1436 => x"a4",
          1437 => x"a4",
          1438 => x"08",
          1439 => x"fc",
          1440 => x"82",
          1441 => x"e0",
          1442 => x"98",
          1443 => x"0c",
          1444 => x"e0",
          1445 => x"82",
          1446 => x"e0",
          1447 => x"73",
          1448 => x"08",
          1449 => x"72",
          1450 => x"72",
          1451 => x"09",
          1452 => x"08",
          1453 => x"71",
          1454 => x"08",
          1455 => x"09",
          1456 => x"e0",
          1457 => x"a4",
          1458 => x"05",
          1459 => x"33",
          1460 => x"82",
          1461 => x"72",
          1462 => x"38",
          1463 => x"70",
          1464 => x"51",
          1465 => x"f8",
          1466 => x"05",
          1467 => x"0c",
          1468 => x"80",
          1469 => x"08",
          1470 => x"38",
          1471 => x"a4",
          1472 => x"08",
          1473 => x"71",
          1474 => x"82",
          1475 => x"a4",
          1476 => x"f4",
          1477 => x"05",
          1478 => x"70",
          1479 => x"a4",
          1480 => x"82",
          1481 => x"72",
          1482 => x"e0",
          1483 => x"39",
          1484 => x"53",
          1485 => x"a4",
          1486 => x"26",
          1487 => x"e0",
          1488 => x"39",
          1489 => x"05",
          1490 => x"f8",
          1491 => x"38",
          1492 => x"53",
          1493 => x"80",
          1494 => x"0c",
          1495 => x"a4",
          1496 => x"e0",
          1497 => x"a4",
          1498 => x"27",
          1499 => x"f8",
          1500 => x"94",
          1501 => x"33",
          1502 => x"a4",
          1503 => x"08",
          1504 => x"72",
          1505 => x"82",
          1506 => x"90",
          1507 => x"08",
          1508 => x"72",
          1509 => x"82",
          1510 => x"72",
          1511 => x"e0",
          1512 => x"39",
          1513 => x"82",
          1514 => x"54",
          1515 => x"82",
          1516 => x"f7",
          1517 => x"33",
          1518 => x"08",
          1519 => x"33",
          1520 => x"05",
          1521 => x"08",
          1522 => x"08",
          1523 => x"82",
          1524 => x"a5",
          1525 => x"33",
          1526 => x"e0",
          1527 => x"e0",
          1528 => x"a4",
          1529 => x"08",
          1530 => x"0b",
          1531 => x"82",
          1532 => x"e0",
          1533 => x"a4",
          1534 => x"08",
          1535 => x"80",
          1536 => x"0c",
          1537 => x"74",
          1538 => x"06",
          1539 => x"80",
          1540 => x"05",
          1541 => x"82",
          1542 => x"54",
          1543 => x"88",
          1544 => x"84",
          1545 => x"b4",
          1546 => x"58",
          1547 => x"54",
          1548 => x"0d",
          1549 => x"0c",
          1550 => x"93",
          1551 => x"82",
          1552 => x"82",
          1553 => x"bd",
          1554 => x"80",
          1555 => x"51",
          1556 => x"80",
          1557 => x"dd",
          1558 => x"39",
          1559 => x"82",
          1560 => x"bf",
          1561 => x"9c",
          1562 => x"b5",
          1563 => x"82",
          1564 => x"84",
          1565 => x"9d",
          1566 => x"82",
          1567 => x"e4",
          1568 => x"85",
          1569 => x"3f",
          1570 => x"77",
          1571 => x"8a",
          1572 => x"51",
          1573 => x"e3",
          1574 => x"75",
          1575 => x"08",
          1576 => x"98",
          1577 => x"0d",
          1578 => x"05",
          1579 => x"68",
          1580 => x"51",
          1581 => x"ff",
          1582 => x"07",
          1583 => x"56",
          1584 => x"52",
          1585 => x"99",
          1586 => x"e0",
          1587 => x"08",
          1588 => x"98",
          1589 => x"84",
          1590 => x"97",
          1591 => x"82",
          1592 => x"74",
          1593 => x"19",
          1594 => x"05",
          1595 => x"70",
          1596 => x"9f",
          1597 => x"74",
          1598 => x"53",
          1599 => x"51",
          1600 => x"e0",
          1601 => x"3d",
          1602 => x"33",
          1603 => x"52",
          1604 => x"98",
          1605 => x"38",
          1606 => x"82",
          1607 => x"82",
          1608 => x"78",
          1609 => x"39",
          1610 => x"8a",
          1611 => x"61",
          1612 => x"33",
          1613 => x"5b",
          1614 => x"f1",
          1615 => x"06",
          1616 => x"38",
          1617 => x"38",
          1618 => x"a0",
          1619 => x"ff",
          1620 => x"ff",
          1621 => x"27",
          1622 => x"38",
          1623 => x"39",
          1624 => x"38",
          1625 => x"ff",
          1626 => x"dc",
          1627 => x"55",
          1628 => x"7a",
          1629 => x"c1",
          1630 => x"39",
          1631 => x"3f",
          1632 => x"53",
          1633 => x"52",
          1634 => x"3f",
          1635 => x"ad",
          1636 => x"fc",
          1637 => x"fe",
          1638 => x"ad",
          1639 => x"80",
          1640 => x"53",
          1641 => x"81",
          1642 => x"38",
          1643 => x"ff",
          1644 => x"38",
          1645 => x"fb",
          1646 => x"82",
          1647 => x"e8",
          1648 => x"82",
          1649 => x"19",
          1650 => x"e0",
          1651 => x"70",
          1652 => x"09",
          1653 => x"c8",
          1654 => x"70",
          1655 => x"72",
          1656 => x"73",
          1657 => x"57",
          1658 => x"76",
          1659 => x"53",
          1660 => x"53",
          1661 => x"0d",
          1662 => x"33",
          1663 => x"c1",
          1664 => x"ac",
          1665 => x"a6",
          1666 => x"c2",
          1667 => x"82",
          1668 => x"74",
          1669 => x"86",
          1670 => x"c0",
          1671 => x"81",
          1672 => x"51",
          1673 => x"3f",
          1674 => x"52",
          1675 => x"99",
          1676 => x"b6",
          1677 => x"82",
          1678 => x"80",
          1679 => x"3f",
          1680 => x"80",
          1681 => x"70",
          1682 => x"92",
          1683 => x"c2",
          1684 => x"98",
          1685 => x"06",
          1686 => x"81",
          1687 => x"51",
          1688 => x"3f",
          1689 => x"52",
          1690 => x"98",
          1691 => x"be",
          1692 => x"86",
          1693 => x"80",
          1694 => x"3f",
          1695 => x"80",
          1696 => x"70",
          1697 => x"92",
          1698 => x"c3",
          1699 => x"97",
          1700 => x"06",
          1701 => x"81",
          1702 => x"51",
          1703 => x"3f",
          1704 => x"fb",
          1705 => x"05",
          1706 => x"75",
          1707 => x"db",
          1708 => x"53",
          1709 => x"51",
          1710 => x"08",
          1711 => x"80",
          1712 => x"73",
          1713 => x"0b",
          1714 => x"2e",
          1715 => x"a8",
          1716 => x"af",
          1717 => x"8b",
          1718 => x"e1",
          1719 => x"81",
          1720 => x"82",
          1721 => x"9c",
          1722 => x"06",
          1723 => x"52",
          1724 => x"82",
          1725 => x"cd",
          1726 => x"7e",
          1727 => x"7d",
          1728 => x"98",
          1729 => x"2e",
          1730 => x"59",
          1731 => x"51",
          1732 => x"82",
          1733 => x"82",
          1734 => x"82",
          1735 => x"70",
          1736 => x"a7",
          1737 => x"80",
          1738 => x"b5",
          1739 => x"3f",
          1740 => x"90",
          1741 => x"87",
          1742 => x"38",
          1743 => x"bd",
          1744 => x"ba",
          1745 => x"8a",
          1746 => x"99",
          1747 => x"38",
          1748 => x"c5",
          1749 => x"38",
          1750 => x"80",
          1751 => x"f8",
          1752 => x"78",
          1753 => x"81",
          1754 => x"2e",
          1755 => x"81",
          1756 => x"39",
          1757 => x"84",
          1758 => x"98",
          1759 => x"3d",
          1760 => x"51",
          1761 => x"80",
          1762 => x"f8",
          1763 => x"81",
          1764 => x"82",
          1765 => x"51",
          1766 => x"5a",
          1767 => x"59",
          1768 => x"7a",
          1769 => x"b5",
          1770 => x"05",
          1771 => x"08",
          1772 => x"fe",
          1773 => x"eb",
          1774 => x"2e",
          1775 => x"11",
          1776 => x"3f",
          1777 => x"b2",
          1778 => x"f6",
          1779 => x"89",
          1780 => x"5b",
          1781 => x"eb",
          1782 => x"ff",
          1783 => x"e0",
          1784 => x"b5",
          1785 => x"05",
          1786 => x"08",
          1787 => x"fe",
          1788 => x"ea",
          1789 => x"2e",
          1790 => x"ff",
          1791 => x"27",
          1792 => x"5e",
          1793 => x"78",
          1794 => x"52",
          1795 => x"3f",
          1796 => x"d5",
          1797 => x"92",
          1798 => x"ff",
          1799 => x"e0",
          1800 => x"fc",
          1801 => x"82",
          1802 => x"82",
          1803 => x"88",
          1804 => x"39",
          1805 => x"2e",
          1806 => x"ab",
          1807 => x"80",
          1808 => x"45",
          1809 => x"78",
          1810 => x"08",
          1811 => x"fc",
          1812 => x"11",
          1813 => x"3f",
          1814 => x"82",
          1815 => x"89",
          1816 => x"cc",
          1817 => x"80",
          1818 => x"44",
          1819 => x"78",
          1820 => x"08",
          1821 => x"59",
          1822 => x"d0",
          1823 => x"33",
          1824 => x"de",
          1825 => x"e4",
          1826 => x"f8",
          1827 => x"81",
          1828 => x"a7",
          1829 => x"2e",
          1830 => x"70",
          1831 => x"7f",
          1832 => x"2e",
          1833 => x"88",
          1834 => x"c1",
          1835 => x"63",
          1836 => x"c5",
          1837 => x"ff",
          1838 => x"e7",
          1839 => x"2e",
          1840 => x"11",
          1841 => x"3f",
          1842 => x"38",
          1843 => x"79",
          1844 => x"fe",
          1845 => x"e6",
          1846 => x"38",
          1847 => x"52",
          1848 => x"3f",
          1849 => x"52",
          1850 => x"46",
          1851 => x"e2",
          1852 => x"3d",
          1853 => x"51",
          1854 => x"80",
          1855 => x"cf",
          1856 => x"45",
          1857 => x"ff",
          1858 => x"3d",
          1859 => x"51",
          1860 => x"80",
          1861 => x"f0",
          1862 => x"98",
          1863 => x"a6",
          1864 => x"22",
          1865 => x"42",
          1866 => x"84",
          1867 => x"98",
          1868 => x"70",
          1869 => x"ff",
          1870 => x"53",
          1871 => x"e3",
          1872 => x"ae",
          1873 => x"87",
          1874 => x"b5",
          1875 => x"05",
          1876 => x"08",
          1877 => x"80",
          1878 => x"5b",
          1879 => x"c5",
          1880 => x"9e",
          1881 => x"ff",
          1882 => x"e0",
          1883 => x"b5",
          1884 => x"05",
          1885 => x"08",
          1886 => x"0c",
          1887 => x"fe",
          1888 => x"de",
          1889 => x"38",
          1890 => x"52",
          1891 => x"3f",
          1892 => x"52",
          1893 => x"46",
          1894 => x"8a",
          1895 => x"3d",
          1896 => x"51",
          1897 => x"80",
          1898 => x"59",
          1899 => x"82",
          1900 => x"ff",
          1901 => x"53",
          1902 => x"82",
          1903 => x"38",
          1904 => x"9d",
          1905 => x"3d",
          1906 => x"51",
          1907 => x"80",
          1908 => x"c6",
          1909 => x"59",
          1910 => x"2e",
          1911 => x"52",
          1912 => x"3f",
          1913 => x"ff",
          1914 => x"f4",
          1915 => x"b8",
          1916 => x"92",
          1917 => x"33",
          1918 => x"80",
          1919 => x"82",
          1920 => x"08",
          1921 => x"98",
          1922 => x"51",
          1923 => x"60",
          1924 => x"81",
          1925 => x"c4",
          1926 => x"26",
          1927 => x"2e",
          1928 => x"7a",
          1929 => x"7a",
          1930 => x"82",
          1931 => x"fc",
          1932 => x"b5",
          1933 => x"86",
          1934 => x"ff",
          1935 => x"39",
          1936 => x"53",
          1937 => x"b0",
          1938 => x"39",
          1939 => x"52",
          1940 => x"9d",
          1941 => x"e0",
          1942 => x"54",
          1943 => x"52",
          1944 => x"c6",
          1945 => x"98",
          1946 => x"80",
          1947 => x"7a",
          1948 => x"7a",
          1949 => x"81",
          1950 => x"7a",
          1951 => x"81",
          1952 => x"ff",
          1953 => x"c7",
          1954 => x"51",
          1955 => x"c7",
          1956 => x"9a",
          1957 => x"e0",
          1958 => x"08",
          1959 => x"51",
          1960 => x"90",
          1961 => x"80",
          1962 => x"82",
          1963 => x"c0",
          1964 => x"84",
          1965 => x"82",
          1966 => x"55",
          1967 => x"ca",
          1968 => x"07",
          1969 => x"c0",
          1970 => x"87",
          1971 => x"5a",
          1972 => x"05",
          1973 => x"f8",
          1974 => x"70",
          1975 => x"8a",
          1976 => x"e0",
          1977 => x"ec",
          1978 => x"b1",
          1979 => x"91",
          1980 => x"3d",
          1981 => x"73",
          1982 => x"38",
          1983 => x"81",
          1984 => x"39",
          1985 => x"81",
          1986 => x"54",
          1987 => x"06",
          1988 => x"80",
          1989 => x"83",
          1990 => x"38",
          1991 => x"52",
          1992 => x"2e",
          1993 => x"84",
          1994 => x"52",
          1995 => x"83",
          1996 => x"30",
          1997 => x"51",
          1998 => x"70",
          1999 => x"72",
          2000 => x"3d",
          2001 => x"72",
          2002 => x"fc",
          2003 => x"82",
          2004 => x"83",
          2005 => x"0c",
          2006 => x"76",
          2007 => x"81",
          2008 => x"83",
          2009 => x"70",
          2010 => x"33",
          2011 => x"fe",
          2012 => x"70",
          2013 => x"33",
          2014 => x"e6",
          2015 => x"74",
          2016 => x"13",
          2017 => x"26",
          2018 => x"98",
          2019 => x"bc",
          2020 => x"b8",
          2021 => x"b4",
          2022 => x"b0",
          2023 => x"ac",
          2024 => x"a8",
          2025 => x"73",
          2026 => x"87",
          2027 => x"82",
          2028 => x"f3",
          2029 => x"9c",
          2030 => x"bc",
          2031 => x"98",
          2032 => x"87",
          2033 => x"1c",
          2034 => x"79",
          2035 => x"08",
          2036 => x"98",
          2037 => x"87",
          2038 => x"1c",
          2039 => x"79",
          2040 => x"83",
          2041 => x"ff",
          2042 => x"1b",
          2043 => x"1b",
          2044 => x"83",
          2045 => x"51",
          2046 => x"04",
          2047 => x"53",
          2048 => x"06",
          2049 => x"70",
          2050 => x"51",
          2051 => x"97",
          2052 => x"e0",
          2053 => x"51",
          2054 => x"9e",
          2055 => x"81",
          2056 => x"32",
          2057 => x"51",
          2058 => x"82",
          2059 => x"fd",
          2060 => x"88",
          2061 => x"82",
          2062 => x"2c",
          2063 => x"73",
          2064 => x"98",
          2065 => x"0d",
          2066 => x"33",
          2067 => x"87",
          2068 => x"86",
          2069 => x"08",
          2070 => x"54",
          2071 => x"91",
          2072 => x"d7",
          2073 => x"51",
          2074 => x"93",
          2075 => x"ff",
          2076 => x"87",
          2077 => x"86",
          2078 => x"72",
          2079 => x"3d",
          2080 => x"05",
          2081 => x"52",
          2082 => x"3d",
          2083 => x"05",
          2084 => x"06",
          2085 => x"3f",
          2086 => x"06",
          2087 => x"76",
          2088 => x"94",
          2089 => x"81",
          2090 => x"8c",
          2091 => x"51",
          2092 => x"70",
          2093 => x"8d",
          2094 => x"51",
          2095 => x"ff",
          2096 => x"72",
          2097 => x"90",
          2098 => x"e0",
          2099 => x"3d",
          2100 => x"81",
          2101 => x"2e",
          2102 => x"81",
          2103 => x"ff",
          2104 => x"94",
          2105 => x"87",
          2106 => x"96",
          2107 => x"70",
          2108 => x"70",
          2109 => x"72",
          2110 => x"70",
          2111 => x"70",
          2112 => x"38",
          2113 => x"94",
          2114 => x"87",
          2115 => x"81",
          2116 => x"53",
          2117 => x"82",
          2118 => x"fe",
          2119 => x"81",
          2120 => x"84",
          2121 => x"c0",
          2122 => x"2a",
          2123 => x"80",
          2124 => x"51",
          2125 => x"2e",
          2126 => x"71",
          2127 => x"98",
          2128 => x"af",
          2129 => x"06",
          2130 => x"0d",
          2131 => x"06",
          2132 => x"70",
          2133 => x"94",
          2134 => x"81",
          2135 => x"80",
          2136 => x"51",
          2137 => x"2e",
          2138 => x"71",
          2139 => x"51",
          2140 => x"84",
          2141 => x"c0",
          2142 => x"06",
          2143 => x"38",
          2144 => x"b4",
          2145 => x"de",
          2146 => x"82",
          2147 => x"08",
          2148 => x"9c",
          2149 => x"9e",
          2150 => x"c0",
          2151 => x"87",
          2152 => x"0c",
          2153 => x"d4",
          2154 => x"de",
          2155 => x"82",
          2156 => x"08",
          2157 => x"c4",
          2158 => x"9e",
          2159 => x"23",
          2160 => x"ec",
          2161 => x"de",
          2162 => x"82",
          2163 => x"f8",
          2164 => x"08",
          2165 => x"52",
          2166 => x"71",
          2167 => x"c0",
          2168 => x"06",
          2169 => x"38",
          2170 => x"80",
          2171 => x"90",
          2172 => x"80",
          2173 => x"de",
          2174 => x"90",
          2175 => x"52",
          2176 => x"52",
          2177 => x"87",
          2178 => x"80",
          2179 => x"83",
          2180 => x"34",
          2181 => x"70",
          2182 => x"70",
          2183 => x"82",
          2184 => x"9e",
          2185 => x"51",
          2186 => x"81",
          2187 => x"0b",
          2188 => x"80",
          2189 => x"2e",
          2190 => x"80",
          2191 => x"08",
          2192 => x"52",
          2193 => x"71",
          2194 => x"c0",
          2195 => x"06",
          2196 => x"38",
          2197 => x"80",
          2198 => x"a0",
          2199 => x"2e",
          2200 => x"83",
          2201 => x"98",
          2202 => x"51",
          2203 => x"87",
          2204 => x"06",
          2205 => x"38",
          2206 => x"87",
          2207 => x"06",
          2208 => x"82",
          2209 => x"9e",
          2210 => x"52",
          2211 => x"71",
          2212 => x"90",
          2213 => x"82",
          2214 => x"fb",
          2215 => x"89",
          2216 => x"73",
          2217 => x"51",
          2218 => x"51",
          2219 => x"33",
          2220 => x"de",
          2221 => x"54",
          2222 => x"96",
          2223 => x"80",
          2224 => x"82",
          2225 => x"c8",
          2226 => x"de",
          2227 => x"38",
          2228 => x"08",
          2229 => x"ff",
          2230 => x"54",
          2231 => x"bc",
          2232 => x"52",
          2233 => x"3f",
          2234 => x"2e",
          2235 => x"de",
          2236 => x"cc",
          2237 => x"83",
          2238 => x"82",
          2239 => x"51",
          2240 => x"33",
          2241 => x"df",
          2242 => x"ff",
          2243 => x"54",
          2244 => x"86",
          2245 => x"87",
          2246 => x"73",
          2247 => x"51",
          2248 => x"33",
          2249 => x"ca",
          2250 => x"df",
          2251 => x"38",
          2252 => x"3f",
          2253 => x"2e",
          2254 => x"a3",
          2255 => x"73",
          2256 => x"51",
          2257 => x"51",
          2258 => x"08",
          2259 => x"ee",
          2260 => x"cb",
          2261 => x"de",
          2262 => x"ff",
          2263 => x"ff",
          2264 => x"52",
          2265 => x"3f",
          2266 => x"c0",
          2267 => x"82",
          2268 => x"76",
          2269 => x"08",
          2270 => x"96",
          2271 => x"80",
          2272 => x"56",
          2273 => x"b7",
          2274 => x"84",
          2275 => x"82",
          2276 => x"51",
          2277 => x"33",
          2278 => x"de",
          2279 => x"75",
          2280 => x"98",
          2281 => x"31",
          2282 => x"82",
          2283 => x"8a",
          2284 => x"0d",
          2285 => x"33",
          2286 => x"38",
          2287 => x"52",
          2288 => x"9d",
          2289 => x"82",
          2290 => x"d4",
          2291 => x"85",
          2292 => x"e6",
          2293 => x"80",
          2294 => x"84",
          2295 => x"c0",
          2296 => x"76",
          2297 => x"2b",
          2298 => x"82",
          2299 => x"80",
          2300 => x"53",
          2301 => x"e8",
          2302 => x"05",
          2303 => x"72",
          2304 => x"53",
          2305 => x"0d",
          2306 => x"05",
          2307 => x"54",
          2308 => x"fc",
          2309 => x"3f",
          2310 => x"ff",
          2311 => x"52",
          2312 => x"33",
          2313 => x"81",
          2314 => x"ff",
          2315 => x"3d",
          2316 => x"84",
          2317 => x"bb",
          2318 => x"84",
          2319 => x"51",
          2320 => x"2e",
          2321 => x"82",
          2322 => x"df",
          2323 => x"56",
          2324 => x"08",
          2325 => x"84",
          2326 => x"51",
          2327 => x"75",
          2328 => x"d3",
          2329 => x"55",
          2330 => x"ff",
          2331 => x"80",
          2332 => x"2e",
          2333 => x"75",
          2334 => x"33",
          2335 => x"05",
          2336 => x"80",
          2337 => x"52",
          2338 => x"df",
          2339 => x"8c",
          2340 => x"df",
          2341 => x"71",
          2342 => x"d3",
          2343 => x"14",
          2344 => x"80",
          2345 => x"e4",
          2346 => x"71",
          2347 => x"e4",
          2348 => x"82",
          2349 => x"dc",
          2350 => x"df",
          2351 => x"82",
          2352 => x"df",
          2353 => x"3d",
          2354 => x"82",
          2355 => x"75",
          2356 => x"98",
          2357 => x"08",
          2358 => x"ff",
          2359 => x"34",
          2360 => x"d0",
          2361 => x"74",
          2362 => x"38",
          2363 => x"aa",
          2364 => x"81",
          2365 => x"e4",
          2366 => x"e0",
          2367 => x"82",
          2368 => x"52",
          2369 => x"c7",
          2370 => x"a5",
          2371 => x"82",
          2372 => x"80",
          2373 => x"38",
          2374 => x"17",
          2375 => x"70",
          2376 => x"55",
          2377 => x"ff",
          2378 => x"11",
          2379 => x"82",
          2380 => x"82",
          2381 => x"78",
          2382 => x"75",
          2383 => x"79",
          2384 => x"08",
          2385 => x"80",
          2386 => x"3d",
          2387 => x"71",
          2388 => x"58",
          2389 => x"38",
          2390 => x"27",
          2391 => x"71",
          2392 => x"09",
          2393 => x"ea",
          2394 => x"df",
          2395 => x"a6",
          2396 => x"79",
          2397 => x"3f",
          2398 => x"84",
          2399 => x"38",
          2400 => x"fc",
          2401 => x"8c",
          2402 => x"c4",
          2403 => x"2e",
          2404 => x"77",
          2405 => x"08",
          2406 => x"74",
          2407 => x"ff",
          2408 => x"8b",
          2409 => x"0c",
          2410 => x"b0",
          2411 => x"08",
          2412 => x"34",
          2413 => x"08",
          2414 => x"82",
          2415 => x"38",
          2416 => x"38",
          2417 => x"80",
          2418 => x"89",
          2419 => x"e4",
          2420 => x"81",
          2421 => x"e0",
          2422 => x"82",
          2423 => x"82",
          2424 => x"80",
          2425 => x"82",
          2426 => x"90",
          2427 => x"3f",
          2428 => x"98",
          2429 => x"d0",
          2430 => x"a4",
          2431 => x"80",
          2432 => x"38",
          2433 => x"17",
          2434 => x"74",
          2435 => x"c2",
          2436 => x"5c",
          2437 => x"5b",
          2438 => x"97",
          2439 => x"34",
          2440 => x"80",
          2441 => x"3d",
          2442 => x"e0",
          2443 => x"51",
          2444 => x"81",
          2445 => x"98",
          2446 => x"33",
          2447 => x"98",
          2448 => x"e8",
          2449 => x"51",
          2450 => x"58",
          2451 => x"38",
          2452 => x"80",
          2453 => x"98",
          2454 => x"ce",
          2455 => x"f6",
          2456 => x"ff",
          2457 => x"74",
          2458 => x"39",
          2459 => x"0a",
          2460 => x"06",
          2461 => x"38",
          2462 => x"cc",
          2463 => x"06",
          2464 => x"56",
          2465 => x"1c",
          2466 => x"98",
          2467 => x"33",
          2468 => x"10",
          2469 => x"11",
          2470 => x"51",
          2471 => x"fe",
          2472 => x"7d",
          2473 => x"80",
          2474 => x"75",
          2475 => x"d0",
          2476 => x"0c",
          2477 => x"38",
          2478 => x"54",
          2479 => x"54",
          2480 => x"f7",
          2481 => x"38",
          2482 => x"55",
          2483 => x"54",
          2484 => x"80",
          2485 => x"98",
          2486 => x"55",
          2487 => x"11",
          2488 => x"73",
          2489 => x"82",
          2490 => x"89",
          2491 => x"d8",
          2492 => x"80",
          2493 => x"98",
          2494 => x"56",
          2495 => x"fb",
          2496 => x"52",
          2497 => x"80",
          2498 => x"98",
          2499 => x"55",
          2500 => x"dc",
          2501 => x"82",
          2502 => x"74",
          2503 => x"fc",
          2504 => x"3f",
          2505 => x"0a",
          2506 => x"33",
          2507 => x"38",
          2508 => x"0b",
          2509 => x"80",
          2510 => x"3f",
          2511 => x"70",
          2512 => x"2e",
          2513 => x"ff",
          2514 => x"ff",
          2515 => x"82",
          2516 => x"96",
          2517 => x"98",
          2518 => x"33",
          2519 => x"ad",
          2520 => x"74",
          2521 => x"33",
          2522 => x"80",
          2523 => x"98",
          2524 => x"55",
          2525 => x"fc",
          2526 => x"3f",
          2527 => x"70",
          2528 => x"51",
          2529 => x"38",
          2530 => x"ff",
          2531 => x"29",
          2532 => x"82",
          2533 => x"75",
          2534 => x"f7",
          2535 => x"34",
          2536 => x"ff",
          2537 => x"79",
          2538 => x"08",
          2539 => x"82",
          2540 => x"8f",
          2541 => x"f1",
          2542 => x"80",
          2543 => x"82",
          2544 => x"0c",
          2545 => x"33",
          2546 => x"82",
          2547 => x"94",
          2548 => x"05",
          2549 => x"81",
          2550 => x"dc",
          2551 => x"73",
          2552 => x"54",
          2553 => x"2b",
          2554 => x"56",
          2555 => x"74",
          2556 => x"82",
          2557 => x"ff",
          2558 => x"29",
          2559 => x"82",
          2560 => x"75",
          2561 => x"52",
          2562 => x"f7",
          2563 => x"2c",
          2564 => x"57",
          2565 => x"fb",
          2566 => x"b0",
          2567 => x"80",
          2568 => x"d8",
          2569 => x"de",
          2570 => x"33",
          2571 => x"33",
          2572 => x"e6",
          2573 => x"14",
          2574 => x"1a",
          2575 => x"3f",
          2576 => x"06",
          2577 => x"75",
          2578 => x"82",
          2579 => x"b8",
          2580 => x"f7",
          2581 => x"34",
          2582 => x"df",
          2583 => x"38",
          2584 => x"e0",
          2585 => x"e0",
          2586 => x"53",
          2587 => x"3f",
          2588 => x"29",
          2589 => x"56",
          2590 => x"51",
          2591 => x"08",
          2592 => x"08",
          2593 => x"52",
          2594 => x"1b",
          2595 => x"74",
          2596 => x"ff",
          2597 => x"2e",
          2598 => x"90",
          2599 => x"74",
          2600 => x"98",
          2601 => x"98",
          2602 => x"74",
          2603 => x"80",
          2604 => x"94",
          2605 => x"2e",
          2606 => x"3f",
          2607 => x"34",
          2608 => x"81",
          2609 => x"9b",
          2610 => x"ff",
          2611 => x"d8",
          2612 => x"53",
          2613 => x"ec",
          2614 => x"dc",
          2615 => x"d8",
          2616 => x"f5",
          2617 => x"81",
          2618 => x"74",
          2619 => x"88",
          2620 => x"33",
          2621 => x"82",
          2622 => x"8f",
          2623 => x"05",
          2624 => x"c6",
          2625 => x"0b",
          2626 => x"82",
          2627 => x"80",
          2628 => x"9f",
          2629 => x"58",
          2630 => x"15",
          2631 => x"84",
          2632 => x"e0",
          2633 => x"76",
          2634 => x"82",
          2635 => x"80",
          2636 => x"88",
          2637 => x"17",
          2638 => x"84",
          2639 => x"08",
          2640 => x"82",
          2641 => x"3d",
          2642 => x"81",
          2643 => x"12",
          2644 => x"ff",
          2645 => x"98",
          2646 => x"0d",
          2647 => x"aa",
          2648 => x"08",
          2649 => x"2b",
          2650 => x"71",
          2651 => x"05",
          2652 => x"70",
          2653 => x"5b",
          2654 => x"34",
          2655 => x"08",
          2656 => x"82",
          2657 => x"e0",
          2658 => x"12",
          2659 => x"2b",
          2660 => x"52",
          2661 => x"70",
          2662 => x"12",
          2663 => x"83",
          2664 => x"56",
          2665 => x"89",
          2666 => x"e0",
          2667 => x"22",
          2668 => x"33",
          2669 => x"83",
          2670 => x"52",
          2671 => x"33",
          2672 => x"54",
          2673 => x"73",
          2674 => x"70",
          2675 => x"71",
          2676 => x"59",
          2677 => x"87",
          2678 => x"88",
          2679 => x"13",
          2680 => x"88",
          2681 => x"71",
          2682 => x"06",
          2683 => x"53",
          2684 => x"87",
          2685 => x"a2",
          2686 => x"83",
          2687 => x"33",
          2688 => x"15",
          2689 => x"2b",
          2690 => x"55",
          2691 => x"80",
          2692 => x"ab",
          2693 => x"70",
          2694 => x"71",
          2695 => x"81",
          2696 => x"83",
          2697 => x"54",
          2698 => x"74",
          2699 => x"34",
          2700 => x"08",
          2701 => x"71",
          2702 => x"59",
          2703 => x"12",
          2704 => x"ff",
          2705 => x"52",
          2706 => x"15",
          2707 => x"0d",
          2708 => x"9e",
          2709 => x"82",
          2710 => x"2b",
          2711 => x"52",
          2712 => x"13",
          2713 => x"05",
          2714 => x"2a",
          2715 => x"34",
          2716 => x"08",
          2717 => x"71",
          2718 => x"59",
          2719 => x"83",
          2720 => x"88",
          2721 => x"13",
          2722 => x"88",
          2723 => x"33",
          2724 => x"0c",
          2725 => x"3d",
          2726 => x"83",
          2727 => x"53",
          2728 => x"88",
          2729 => x"11",
          2730 => x"71",
          2731 => x"81",
          2732 => x"2b",
          2733 => x"58",
          2734 => x"38",
          2735 => x"9d",
          2736 => x"85",
          2737 => x"2b",
          2738 => x"51",
          2739 => x"75",
          2740 => x"34",
          2741 => x"12",
          2742 => x"07",
          2743 => x"53",
          2744 => x"34",
          2745 => x"0b",
          2746 => x"34",
          2747 => x"14",
          2748 => x"88",
          2749 => x"71",
          2750 => x"07",
          2751 => x"54",
          2752 => x"8b",
          2753 => x"52",
          2754 => x"f1",
          2755 => x"51",
          2756 => x"f5",
          2757 => x"e2",
          2758 => x"ff",
          2759 => x"33",
          2760 => x"70",
          2761 => x"ff",
          2762 => x"75",
          2763 => x"33",
          2764 => x"ff",
          2765 => x"06",
          2766 => x"59",
          2767 => x"80",
          2768 => x"84",
          2769 => x"2b",
          2770 => x"81",
          2771 => x"59",
          2772 => x"88",
          2773 => x"71",
          2774 => x"06",
          2775 => x"75",
          2776 => x"79",
          2777 => x"74",
          2778 => x"2e",
          2779 => x"f8",
          2780 => x"80",
          2781 => x"3f",
          2782 => x"11",
          2783 => x"71",
          2784 => x"74",
          2785 => x"06",
          2786 => x"78",
          2787 => x"57",
          2788 => x"08",
          2789 => x"86",
          2790 => x"2b",
          2791 => x"53",
          2792 => x"75",
          2793 => x"70",
          2794 => x"71",
          2795 => x"5d",
          2796 => x"15",
          2797 => x"88",
          2798 => x"33",
          2799 => x"70",
          2800 => x"54",
          2801 => x"34",
          2802 => x"54",
          2803 => x"0d",
          2804 => x"e0",
          2805 => x"71",
          2806 => x"51",
          2807 => x"53",
          2808 => x"0d",
          2809 => x"5c",
          2810 => x"08",
          2811 => x"f4",
          2812 => x"ff",
          2813 => x"83",
          2814 => x"fc",
          2815 => x"7e",
          2816 => x"08",
          2817 => x"08",
          2818 => x"ff",
          2819 => x"70",
          2820 => x"07",
          2821 => x"06",
          2822 => x"29",
          2823 => x"88",
          2824 => x"4e",
          2825 => x"41",
          2826 => x"8f",
          2827 => x"31",
          2828 => x"82",
          2829 => x"2b",
          2830 => x"81",
          2831 => x"2b",
          2832 => x"73",
          2833 => x"70",
          2834 => x"7b",
          2835 => x"73",
          2836 => x"78",
          2837 => x"ff",
          2838 => x"38",
          2839 => x"f6",
          2840 => x"55",
          2841 => x"1d",
          2842 => x"88",
          2843 => x"3f",
          2844 => x"82",
          2845 => x"7e",
          2846 => x"e0",
          2847 => x"59",
          2848 => x"08",
          2849 => x"06",
          2850 => x"54",
          2851 => x"51",
          2852 => x"1d",
          2853 => x"88",
          2854 => x"3f",
          2855 => x"82",
          2856 => x"7e",
          2857 => x"e0",
          2858 => x"59",
          2859 => x"08",
          2860 => x"55",
          2861 => x"a9",
          2862 => x"3f",
          2863 => x"98",
          2864 => x"73",
          2865 => x"8b",
          2866 => x"7a",
          2867 => x"53",
          2868 => x"7a",
          2869 => x"05",
          2870 => x"54",
          2871 => x"0d",
          2872 => x"70",
          2873 => x"98",
          2874 => x"2e",
          2875 => x"e0",
          2876 => x"74",
          2877 => x"04",
          2878 => x"51",
          2879 => x"82",
          2880 => x"e0",
          2881 => x"3d",
          2882 => x"05",
          2883 => x"72",
          2884 => x"2b",
          2885 => x"88",
          2886 => x"88",
          2887 => x"8c",
          2888 => x"87",
          2889 => x"08",
          2890 => x"2e",
          2891 => x"51",
          2892 => x"80",
          2893 => x"98",
          2894 => x"38",
          2895 => x"e0",
          2896 => x"98",
          2897 => x"0d",
          2898 => x"05",
          2899 => x"52",
          2900 => x"08",
          2901 => x"be",
          2902 => x"c0",
          2903 => x"12",
          2904 => x"40",
          2905 => x"98",
          2906 => x"0c",
          2907 => x"06",
          2908 => x"38",
          2909 => x"05",
          2910 => x"a2",
          2911 => x"38",
          2912 => x"38",
          2913 => x"98",
          2914 => x"c0",
          2915 => x"87",
          2916 => x"81",
          2917 => x"53",
          2918 => x"71",
          2919 => x"84",
          2920 => x"06",
          2921 => x"38",
          2922 => x"87",
          2923 => x"73",
          2924 => x"2e",
          2925 => x"82",
          2926 => x"f3",
          2927 => x"05",
          2928 => x"83",
          2929 => x"3f",
          2930 => x"54",
          2931 => x"81",
          2932 => x"c0",
          2933 => x"12",
          2934 => x"5f",
          2935 => x"8c",
          2936 => x"80",
          2937 => x"81",
          2938 => x"8c",
          2939 => x"7c",
          2940 => x"70",
          2941 => x"8a",
          2942 => x"71",
          2943 => x"52",
          2944 => x"80",
          2945 => x"c0",
          2946 => x"82",
          2947 => x"19",
          2948 => x"ff",
          2949 => x"78",
          2950 => x"80",
          2951 => x"26",
          2952 => x"06",
          2953 => x"52",
          2954 => x"8f",
          2955 => x"02",
          2956 => x"05",
          2957 => x"57",
          2958 => x"81",
          2959 => x"38",
          2960 => x"81",
          2961 => x"71",
          2962 => x"87",
          2963 => x"80",
          2964 => x"83",
          2965 => x"72",
          2966 => x"51",
          2967 => x"87",
          2968 => x"38",
          2969 => x"96",
          2970 => x"8c",
          2971 => x"51",
          2972 => x"56",
          2973 => x"85",
          2974 => x"83",
          2975 => x"e0",
          2976 => x"3d",
          2977 => x"71",
          2978 => x"53",
          2979 => x"0d",
          2980 => x"71",
          2981 => x"14",
          2982 => x"33",
          2983 => x"53",
          2984 => x"04",
          2985 => x"92",
          2986 => x"81",
          2987 => x"70",
          2988 => x"3d",
          2989 => x"70",
          2990 => x"51",
          2991 => x"70",
          2992 => x"05",
          2993 => x"72",
          2994 => x"0d",
          2995 => x"80",
          2996 => x"53",
          2997 => x"ff",
          2998 => x"04",
          2999 => x"52",
          3000 => x"34",
          3001 => x"3d",
          3002 => x"79",
          3003 => x"56",
          3004 => x"71",
          3005 => x"52",
          3006 => x"2e",
          3007 => x"86",
          3008 => x"76",
          3009 => x"8a",
          3010 => x"71",
          3011 => x"0c",
          3012 => x"e0",
          3013 => x"70",
          3014 => x"70",
          3015 => x"55",
          3016 => x"80",
          3017 => x"51",
          3018 => x"08",
          3019 => x"2e",
          3020 => x"74",
          3021 => x"04",
          3022 => x"83",
          3023 => x"80",
          3024 => x"53",
          3025 => x"52",
          3026 => x"08",
          3027 => x"82",
          3028 => x"16",
          3029 => x"18",
          3030 => x"9f",
          3031 => x"2e",
          3032 => x"76",
          3033 => x"51",
          3034 => x"79",
          3035 => x"04",
          3036 => x"80",
          3037 => x"38",
          3038 => x"98",
          3039 => x"38",
          3040 => x"81",
          3041 => x"e0",
          3042 => x"55",
          3043 => x"82",
          3044 => x"f8",
          3045 => x"c0",
          3046 => x"e0",
          3047 => x"55",
          3048 => x"f0",
          3049 => x"2e",
          3050 => x"80",
          3051 => x"17",
          3052 => x"d4",
          3053 => x"d8",
          3054 => x"75",
          3055 => x"e4",
          3056 => x"de",
          3057 => x"17",
          3058 => x"52",
          3059 => x"a4",
          3060 => x"0c",
          3061 => x"33",
          3062 => x"34",
          3063 => x"51",
          3064 => x"80",
          3065 => x"e0",
          3066 => x"3d",
          3067 => x"fe",
          3068 => x"73",
          3069 => x"71",
          3070 => x"75",
          3071 => x"04",
          3072 => x"56",
          3073 => x"38",
          3074 => x"38",
          3075 => x"2e",
          3076 => x"38",
          3077 => x"39",
          3078 => x"b6",
          3079 => x"2a",
          3080 => x"55",
          3081 => x"81",
          3082 => x"b8",
          3083 => x"a8",
          3084 => x"57",
          3085 => x"08",
          3086 => x"14",
          3087 => x"07",
          3088 => x"52",
          3089 => x"75",
          3090 => x"76",
          3091 => x"73",
          3092 => x"08",
          3093 => x"06",
          3094 => x"3f",
          3095 => x"06",
          3096 => x"15",
          3097 => x"3f",
          3098 => x"82",
          3099 => x"05",
          3100 => x"08",
          3101 => x"58",
          3102 => x"0d",
          3103 => x"5a",
          3104 => x"82",
          3105 => x"82",
          3106 => x"2e",
          3107 => x"38",
          3108 => x"39",
          3109 => x"f7",
          3110 => x"2a",
          3111 => x"55",
          3112 => x"59",
          3113 => x"74",
          3114 => x"16",
          3115 => x"53",
          3116 => x"2b",
          3117 => x"71",
          3118 => x"0b",
          3119 => x"17",
          3120 => x"3f",
          3121 => x"98",
          3122 => x"06",
          3123 => x"54",
          3124 => x"33",
          3125 => x"51",
          3126 => x"76",
          3127 => x"75",
          3128 => x"08",
          3129 => x"38",
          3130 => x"10",
          3131 => x"51",
          3132 => x"2a",
          3133 => x"f9",
          3134 => x"82",
          3135 => x"0a",
          3136 => x"70",
          3137 => x"54",
          3138 => x"8f",
          3139 => x"f6",
          3140 => x"78",
          3141 => x"04",
          3142 => x"08",
          3143 => x"a4",
          3144 => x"38",
          3145 => x"73",
          3146 => x"e0",
          3147 => x"80",
          3148 => x"eb",
          3149 => x"e0",
          3150 => x"52",
          3151 => x"98",
          3152 => x"2e",
          3153 => x"81",
          3154 => x"ff",
          3155 => x"75",
          3156 => x"08",
          3157 => x"94",
          3158 => x"27",
          3159 => x"84",
          3160 => x"17",
          3161 => x"a6",
          3162 => x"0c",
          3163 => x"7c",
          3164 => x"95",
          3165 => x"2e",
          3166 => x"b2",
          3167 => x"7a",
          3168 => x"82",
          3169 => x"82",
          3170 => x"08",
          3171 => x"08",
          3172 => x"38",
          3173 => x"54",
          3174 => x"7a",
          3175 => x"81",
          3176 => x"83",
          3177 => x"f9",
          3178 => x"08",
          3179 => x"82",
          3180 => x"08",
          3181 => x"25",
          3182 => x"54",
          3183 => x"38",
          3184 => x"38",
          3185 => x"90",
          3186 => x"38",
          3187 => x"38",
          3188 => x"08",
          3189 => x"78",
          3190 => x"51",
          3191 => x"80",
          3192 => x"98",
          3193 => x"38",
          3194 => x"98",
          3195 => x"80",
          3196 => x"55",
          3197 => x"09",
          3198 => x"80",
          3199 => x"51",
          3200 => x"82",
          3201 => x"98",
          3202 => x"79",
          3203 => x"8f",
          3204 => x"f9",
          3205 => x"74",
          3206 => x"17",
          3207 => x"54",
          3208 => x"94",
          3209 => x"54",
          3210 => x"56",
          3211 => x"80",
          3212 => x"55",
          3213 => x"82",
          3214 => x"f8",
          3215 => x"f0",
          3216 => x"56",
          3217 => x"7b",
          3218 => x"e0",
          3219 => x"17",
          3220 => x"b8",
          3221 => x"77",
          3222 => x"15",
          3223 => x"81",
          3224 => x"15",
          3225 => x"98",
          3226 => x"22",
          3227 => x"70",
          3228 => x"82",
          3229 => x"f8",
          3230 => x"56",
          3231 => x"f1",
          3232 => x"e9",
          3233 => x"08",
          3234 => x"82",
          3235 => x"54",
          3236 => x"82",
          3237 => x"79",
          3238 => x"98",
          3239 => x"22",
          3240 => x"26",
          3241 => x"b0",
          3242 => x"e0",
          3243 => x"0b",
          3244 => x"9c",
          3245 => x"85",
          3246 => x"31",
          3247 => x"f4",
          3248 => x"18",
          3249 => x"08",
          3250 => x"38",
          3251 => x"89",
          3252 => x"ff",
          3253 => x"80",
          3254 => x"3d",
          3255 => x"08",
          3256 => x"54",
          3257 => x"80",
          3258 => x"53",
          3259 => x"38",
          3260 => x"b5",
          3261 => x"14",
          3262 => x"2a",
          3263 => x"26",
          3264 => x"16",
          3265 => x"53",
          3266 => x"51",
          3267 => x"53",
          3268 => x"08",
          3269 => x"e0",
          3270 => x"9c",
          3271 => x"80",
          3272 => x"15",
          3273 => x"14",
          3274 => x"82",
          3275 => x"e0",
          3276 => x"82",
          3277 => x"ba",
          3278 => x"ff",
          3279 => x"52",
          3280 => x"98",
          3281 => x"72",
          3282 => x"e0",
          3283 => x"15",
          3284 => x"0c",
          3285 => x"8a",
          3286 => x"7d",
          3287 => x"76",
          3288 => x"08",
          3289 => x"38",
          3290 => x"08",
          3291 => x"e0",
          3292 => x"80",
          3293 => x"18",
          3294 => x"81",
          3295 => x"81",
          3296 => x"83",
          3297 => x"72",
          3298 => x"75",
          3299 => x"a5",
          3300 => x"52",
          3301 => x"98",
          3302 => x"2e",
          3303 => x"81",
          3304 => x"e0",
          3305 => x"3d",
          3306 => x"ae",
          3307 => x"ff",
          3308 => x"71",
          3309 => x"94",
          3310 => x"98",
          3311 => x"82",
          3312 => x"fc",
          3313 => x"ff",
          3314 => x"eb",
          3315 => x"72",
          3316 => x"73",
          3317 => x"98",
          3318 => x"0d",
          3319 => x"81",
          3320 => x"70",
          3321 => x"81",
          3322 => x"51",
          3323 => x"0c",
          3324 => x"60",
          3325 => x"5b",
          3326 => x"08",
          3327 => x"08",
          3328 => x"e0",
          3329 => x"82",
          3330 => x"55",
          3331 => x"dc",
          3332 => x"81",
          3333 => x"34",
          3334 => x"e5",
          3335 => x"56",
          3336 => x"2e",
          3337 => x"75",
          3338 => x"e0",
          3339 => x"72",
          3340 => x"81",
          3341 => x"ff",
          3342 => x"09",
          3343 => x"2a",
          3344 => x"2e",
          3345 => x"bf",
          3346 => x"0c",
          3347 => x"81",
          3348 => x"53",
          3349 => x"8f",
          3350 => x"5a",
          3351 => x"83",
          3352 => x"38",
          3353 => x"29",
          3354 => x"58",
          3355 => x"51",
          3356 => x"83",
          3357 => x"96",
          3358 => x"38",
          3359 => x"73",
          3360 => x"83",
          3361 => x"38",
          3362 => x"38",
          3363 => x"06",
          3364 => x"38",
          3365 => x"10",
          3366 => x"70",
          3367 => x"81",
          3368 => x"93",
          3369 => x"e0",
          3370 => x"7d",
          3371 => x"0c",
          3372 => x"d2",
          3373 => x"e0",
          3374 => x"fd",
          3375 => x"1a",
          3376 => x"3d",
          3377 => x"08",
          3378 => x"d7",
          3379 => x"e0",
          3380 => x"70",
          3381 => x"98",
          3382 => x"3f",
          3383 => x"98",
          3384 => x"70",
          3385 => x"58",
          3386 => x"06",
          3387 => x"86",
          3388 => x"c3",
          3389 => x"51",
          3390 => x"82",
          3391 => x"06",
          3392 => x"86",
          3393 => x"73",
          3394 => x"81",
          3395 => x"38",
          3396 => x"70",
          3397 => x"5d",
          3398 => x"81",
          3399 => x"76",
          3400 => x"8c",
          3401 => x"b6",
          3402 => x"ff",
          3403 => x"33",
          3404 => x"59",
          3405 => x"a8",
          3406 => x"3f",
          3407 => x"06",
          3408 => x"81",
          3409 => x"80",
          3410 => x"78",
          3411 => x"19",
          3412 => x"82",
          3413 => x"80",
          3414 => x"83",
          3415 => x"38",
          3416 => x"a5",
          3417 => x"81",
          3418 => x"90",
          3419 => x"10",
          3420 => x"38",
          3421 => x"54",
          3422 => x"bb",
          3423 => x"b5",
          3424 => x"06",
          3425 => x"19",
          3426 => x"8b",
          3427 => x"51",
          3428 => x"80",
          3429 => x"0b",
          3430 => x"f5",
          3431 => x"82",
          3432 => x"38",
          3433 => x"0d",
          3434 => x"ab",
          3435 => x"5a",
          3436 => x"8c",
          3437 => x"73",
          3438 => x"10",
          3439 => x"39",
          3440 => x"3d",
          3441 => x"02",
          3442 => x"73",
          3443 => x"0b",
          3444 => x"08",
          3445 => x"78",
          3446 => x"80",
          3447 => x"83",
          3448 => x"2e",
          3449 => x"82",
          3450 => x"06",
          3451 => x"90",
          3452 => x"56",
          3453 => x"a0",
          3454 => x"80",
          3455 => x"87",
          3456 => x"74",
          3457 => x"27",
          3458 => x"34",
          3459 => x"57",
          3460 => x"ec",
          3461 => x"80",
          3462 => x"73",
          3463 => x"33",
          3464 => x"98",
          3465 => x"54",
          3466 => x"55",
          3467 => x"38",
          3468 => x"39",
          3469 => x"78",
          3470 => x"76",
          3471 => x"15",
          3472 => x"34",
          3473 => x"f9",
          3474 => x"38",
          3475 => x"fe",
          3476 => x"2e",
          3477 => x"55",
          3478 => x"81",
          3479 => x"05",
          3480 => x"05",
          3481 => x"51",
          3482 => x"90",
          3483 => x"eb",
          3484 => x"59",
          3485 => x"82",
          3486 => x"08",
          3487 => x"80",
          3488 => x"90",
          3489 => x"51",
          3490 => x"57",
          3491 => x"a0",
          3492 => x"98",
          3493 => x"08",
          3494 => x"e0",
          3495 => x"81",
          3496 => x"08",
          3497 => x"7c",
          3498 => x"34",
          3499 => x"82",
          3500 => x"df",
          3501 => x"77",
          3502 => x"8b",
          3503 => x"17",
          3504 => x"a8",
          3505 => x"3f",
          3506 => x"81",
          3507 => x"73",
          3508 => x"10",
          3509 => x"38",
          3510 => x"34",
          3511 => x"79",
          3512 => x"08",
          3513 => x"38",
          3514 => x"98",
          3515 => x"3f",
          3516 => x"98",
          3517 => x"98",
          3518 => x"c0",
          3519 => x"1a",
          3520 => x"08",
          3521 => x"73",
          3522 => x"34",
          3523 => x"94",
          3524 => x"70",
          3525 => x"56",
          3526 => x"38",
          3527 => x"82",
          3528 => x"08",
          3529 => x"75",
          3530 => x"08",
          3531 => x"9c",
          3532 => x"0b",
          3533 => x"27",
          3534 => x"74",
          3535 => x"08",
          3536 => x"c3",
          3537 => x"83",
          3538 => x"0c",
          3539 => x"7e",
          3540 => x"0b",
          3541 => x"2e",
          3542 => x"2e",
          3543 => x"8c",
          3544 => x"5c",
          3545 => x"78",
          3546 => x"56",
          3547 => x"15",
          3548 => x"72",
          3549 => x"80",
          3550 => x"ff",
          3551 => x"52",
          3552 => x"d7",
          3553 => x"ff",
          3554 => x"95",
          3555 => x"88",
          3556 => x"15",
          3557 => x"76",
          3558 => x"80",
          3559 => x"2e",
          3560 => x"7a",
          3561 => x"5b",
          3562 => x"22",
          3563 => x"7a",
          3564 => x"06",
          3565 => x"53",
          3566 => x"89",
          3567 => x"19",
          3568 => x"74",
          3569 => x"09",
          3570 => x"78",
          3571 => x"80",
          3572 => x"90",
          3573 => x"76",
          3574 => x"57",
          3575 => x"81",
          3576 => x"38",
          3577 => x"81",
          3578 => x"81",
          3579 => x"96",
          3580 => x"72",
          3581 => x"72",
          3582 => x"89",
          3583 => x"11",
          3584 => x"9c",
          3585 => x"88",
          3586 => x"53",
          3587 => x"81",
          3588 => x"a0",
          3589 => x"53",
          3590 => x"81",
          3591 => x"56",
          3592 => x"77",
          3593 => x"14",
          3594 => x"51",
          3595 => x"34",
          3596 => x"88",
          3597 => x"52",
          3598 => x"08",
          3599 => x"3f",
          3600 => x"98",
          3601 => x"98",
          3602 => x"04",
          3603 => x"5e",
          3604 => x"73",
          3605 => x"80",
          3606 => x"8d",
          3607 => x"0c",
          3608 => x"70",
          3609 => x"09",
          3610 => x"80",
          3611 => x"78",
          3612 => x"73",
          3613 => x"54",
          3614 => x"0b",
          3615 => x"e7",
          3616 => x"87",
          3617 => x"11",
          3618 => x"fc",
          3619 => x"98",
          3620 => x"ff",
          3621 => x"92",
          3622 => x"08",
          3623 => x"81",
          3624 => x"ff",
          3625 => x"9f",
          3626 => x"51",
          3627 => x"dc",
          3628 => x"91",
          3629 => x"d9",
          3630 => x"de",
          3631 => x"38",
          3632 => x"81",
          3633 => x"41",
          3634 => x"73",
          3635 => x"81",
          3636 => x"70",
          3637 => x"73",
          3638 => x"82",
          3639 => x"06",
          3640 => x"2e",
          3641 => x"2e",
          3642 => x"1a",
          3643 => x"06",
          3644 => x"ae",
          3645 => x"10",
          3646 => x"a0",
          3647 => x"26",
          3648 => x"81",
          3649 => x"78",
          3650 => x"73",
          3651 => x"80",
          3652 => x"05",
          3653 => x"a0",
          3654 => x"51",
          3655 => x"84",
          3656 => x"78",
          3657 => x"56",
          3658 => x"56",
          3659 => x"83",
          3660 => x"ff",
          3661 => x"2e",
          3662 => x"70",
          3663 => x"73",
          3664 => x"74",
          3665 => x"2e",
          3666 => x"07",
          3667 => x"16",
          3668 => x"ae",
          3669 => x"05",
          3670 => x"8f",
          3671 => x"73",
          3672 => x"8b",
          3673 => x"e8",
          3674 => x"7c",
          3675 => x"57",
          3676 => x"75",
          3677 => x"70",
          3678 => x"7c",
          3679 => x"89",
          3680 => x"80",
          3681 => x"38",
          3682 => x"70",
          3683 => x"51",
          3684 => x"38",
          3685 => x"79",
          3686 => x"7c",
          3687 => x"88",
          3688 => x"06",
          3689 => x"76",
          3690 => x"83",
          3691 => x"3f",
          3692 => x"06",
          3693 => x"55",
          3694 => x"80",
          3695 => x"57",
          3696 => x"ff",
          3697 => x"76",
          3698 => x"39",
          3699 => x"55",
          3700 => x"80",
          3701 => x"75",
          3702 => x"3f",
          3703 => x"38",
          3704 => x"a4",
          3705 => x"26",
          3706 => x"9f",
          3707 => x"7b",
          3708 => x"ff",
          3709 => x"05",
          3710 => x"fd",
          3711 => x"81",
          3712 => x"85",
          3713 => x"09",
          3714 => x"81",
          3715 => x"73",
          3716 => x"54",
          3717 => x"38",
          3718 => x"70",
          3719 => x"7b",
          3720 => x"38",
          3721 => x"70",
          3722 => x"85",
          3723 => x"1f",
          3724 => x"e0",
          3725 => x"82",
          3726 => x"82",
          3727 => x"06",
          3728 => x"81",
          3729 => x"73",
          3730 => x"54",
          3731 => x"80",
          3732 => x"c2",
          3733 => x"38",
          3734 => x"70",
          3735 => x"86",
          3736 => x"06",
          3737 => x"38",
          3738 => x"05",
          3739 => x"3f",
          3740 => x"f8",
          3741 => x"92",
          3742 => x"5b",
          3743 => x"59",
          3744 => x"c6",
          3745 => x"70",
          3746 => x"8d",
          3747 => x"09",
          3748 => x"d0",
          3749 => x"53",
          3750 => x"73",
          3751 => x"71",
          3752 => x"82",
          3753 => x"55",
          3754 => x"74",
          3755 => x"12",
          3756 => x"38",
          3757 => x"51",
          3758 => x"89",
          3759 => x"53",
          3760 => x"51",
          3761 => x"38",
          3762 => x"77",
          3763 => x"2a",
          3764 => x"51",
          3765 => x"84",
          3766 => x"94",
          3767 => x"38",
          3768 => x"86",
          3769 => x"82",
          3770 => x"fa",
          3771 => x"17",
          3772 => x"52",
          3773 => x"82",
          3774 => x"b6",
          3775 => x"98",
          3776 => x"55",
          3777 => x"06",
          3778 => x"33",
          3779 => x"81",
          3780 => x"eb",
          3781 => x"07",
          3782 => x"81",
          3783 => x"83",
          3784 => x"16",
          3785 => x"08",
          3786 => x"9d",
          3787 => x"81",
          3788 => x"e0",
          3789 => x"80",
          3790 => x"e0",
          3791 => x"3d",
          3792 => x"05",
          3793 => x"51",
          3794 => x"58",
          3795 => x"08",
          3796 => x"08",
          3797 => x"08",
          3798 => x"87",
          3799 => x"fe",
          3800 => x"2e",
          3801 => x"a0",
          3802 => x"06",
          3803 => x"38",
          3804 => x"82",
          3805 => x"56",
          3806 => x"80",
          3807 => x"8c",
          3808 => x"81",
          3809 => x"e0",
          3810 => x"06",
          3811 => x"38",
          3812 => x"2a",
          3813 => x"72",
          3814 => x"52",
          3815 => x"08",
          3816 => x"93",
          3817 => x"82",
          3818 => x"2e",
          3819 => x"59",
          3820 => x"58",
          3821 => x"fe",
          3822 => x"98",
          3823 => x"5b",
          3824 => x"75",
          3825 => x"e0",
          3826 => x"2a",
          3827 => x"29",
          3828 => x"57",
          3829 => x"80",
          3830 => x"fc",
          3831 => x"ff",
          3832 => x"1a",
          3833 => x"81",
          3834 => x"27",
          3835 => x"81",
          3836 => x"27",
          3837 => x"84",
          3838 => x"84",
          3839 => x"86",
          3840 => x"ff",
          3841 => x"81",
          3842 => x"51",
          3843 => x"83",
          3844 => x"80",
          3845 => x"e0",
          3846 => x"80",
          3847 => x"c8",
          3848 => x"06",
          3849 => x"26",
          3850 => x"78",
          3851 => x"59",
          3852 => x"2e",
          3853 => x"72",
          3854 => x"f2",
          3855 => x"3f",
          3856 => x"98",
          3857 => x"57",
          3858 => x"cb",
          3859 => x"98",
          3860 => x"8d",
          3861 => x"3f",
          3862 => x"14",
          3863 => x"08",
          3864 => x"72",
          3865 => x"22",
          3866 => x"5a",
          3867 => x"14",
          3868 => x"d3",
          3869 => x"82",
          3870 => x"38",
          3871 => x"ff",
          3872 => x"83",
          3873 => x"74",
          3874 => x"89",
          3875 => x"ca",
          3876 => x"7b",
          3877 => x"17",
          3878 => x"55",
          3879 => x"38",
          3880 => x"82",
          3881 => x"53",
          3882 => x"82",
          3883 => x"bd",
          3884 => x"0c",
          3885 => x"56",
          3886 => x"13",
          3887 => x"82",
          3888 => x"81",
          3889 => x"83",
          3890 => x"72",
          3891 => x"ff",
          3892 => x"15",
          3893 => x"76",
          3894 => x"38",
          3895 => x"82",
          3896 => x"53",
          3897 => x"f9",
          3898 => x"88",
          3899 => x"38",
          3900 => x"84",
          3901 => x"e0",
          3902 => x"72",
          3903 => x"80",
          3904 => x"3f",
          3905 => x"a4",
          3906 => x"84",
          3907 => x"e0",
          3908 => x"2e",
          3909 => x"14",
          3910 => x"08",
          3911 => x"c5",
          3912 => x"15",
          3913 => x"22",
          3914 => x"23",
          3915 => x"0b",
          3916 => x"0c",
          3917 => x"90",
          3918 => x"54",
          3919 => x"73",
          3920 => x"72",
          3921 => x"86",
          3922 => x"71",
          3923 => x"81",
          3924 => x"82",
          3925 => x"88",
          3926 => x"39",
          3927 => x"74",
          3928 => x"04",
          3929 => x"7a",
          3930 => x"f4",
          3931 => x"e0",
          3932 => x"98",
          3933 => x"70",
          3934 => x"38",
          3935 => x"2e",
          3936 => x"0c",
          3937 => x"80",
          3938 => x"51",
          3939 => x"54",
          3940 => x"0d",
          3941 => x"05",
          3942 => x"54",
          3943 => x"bf",
          3944 => x"53",
          3945 => x"ae",
          3946 => x"e0",
          3947 => x"69",
          3948 => x"b0",
          3949 => x"e0",
          3950 => x"05",
          3951 => x"80",
          3952 => x"06",
          3953 => x"74",
          3954 => x"09",
          3955 => x"b1",
          3956 => x"39",
          3957 => x"73",
          3958 => x"81",
          3959 => x"38",
          3960 => x"07",
          3961 => x"2a",
          3962 => x"2e",
          3963 => x"d6",
          3964 => x"82",
          3965 => x"51",
          3966 => x"8b",
          3967 => x"51",
          3968 => x"05",
          3969 => x"0b",
          3970 => x"f1",
          3971 => x"80",
          3972 => x"51",
          3973 => x"55",
          3974 => x"b7",
          3975 => x"05",
          3976 => x"51",
          3977 => x"84",
          3978 => x"70",
          3979 => x"a9",
          3980 => x"2e",
          3981 => x"73",
          3982 => x"e0",
          3983 => x"0c",
          3984 => x"f8",
          3985 => x"51",
          3986 => x"80",
          3987 => x"a0",
          3988 => x"53",
          3989 => x"e0",
          3990 => x"1b",
          3991 => x"dd",
          3992 => x"98",
          3993 => x"56",
          3994 => x"90",
          3995 => x"80",
          3996 => x"1a",
          3997 => x"51",
          3998 => x"82",
          3999 => x"38",
          4000 => x"8a",
          4001 => x"59",
          4002 => x"c5",
          4003 => x"82",
          4004 => x"82",
          4005 => x"09",
          4006 => x"78",
          4007 => x"80",
          4008 => x"38",
          4009 => x"c3",
          4010 => x"38",
          4011 => x"2e",
          4012 => x"ee",
          4013 => x"82",
          4014 => x"e0",
          4015 => x"39",
          4016 => x"e0",
          4017 => x"3d",
          4018 => x"5d",
          4019 => x"05",
          4020 => x"e0",
          4021 => x"8a",
          4022 => x"2e",
          4023 => x"90",
          4024 => x"74",
          4025 => x"82",
          4026 => x"ad",
          4027 => x"56",
          4028 => x"1a",
          4029 => x"38",
          4030 => x"38",
          4031 => x"56",
          4032 => x"11",
          4033 => x"5b",
          4034 => x"88",
          4035 => x"08",
          4036 => x"e0",
          4037 => x"9f",
          4038 => x"74",
          4039 => x"7e",
          4040 => x"08",
          4041 => x"98",
          4042 => x"77",
          4043 => x"7f",
          4044 => x"75",
          4045 => x"77",
          4046 => x"33",
          4047 => x"98",
          4048 => x"33",
          4049 => x"b4",
          4050 => x"27",
          4051 => x"52",
          4052 => x"7d",
          4053 => x"89",
          4054 => x"0c",
          4055 => x"80",
          4056 => x"83",
          4057 => x"7e",
          4058 => x"08",
          4059 => x"08",
          4060 => x"7c",
          4061 => x"31",
          4062 => x"94",
          4063 => x"5c",
          4064 => x"e0",
          4065 => x"3d",
          4066 => x"5d",
          4067 => x"05",
          4068 => x"e0",
          4069 => x"8a",
          4070 => x"2e",
          4071 => x"90",
          4072 => x"06",
          4073 => x"2e",
          4074 => x"91",
          4075 => x"81",
          4076 => x"95",
          4077 => x"56",
          4078 => x"5c",
          4079 => x"18",
          4080 => x"74",
          4081 => x"ff",
          4082 => x"7a",
          4083 => x"08",
          4084 => x"39",
          4085 => x"ac",
          4086 => x"e0",
          4087 => x"74",
          4088 => x"2e",
          4089 => x"88",
          4090 => x"0c",
          4091 => x"08",
          4092 => x"51",
          4093 => x"08",
          4094 => x"7e",
          4095 => x"98",
          4096 => x"e0",
          4097 => x"57",
          4098 => x"1b",
          4099 => x"75",
          4100 => x"59",
          4101 => x"1a",
          4102 => x"e0",
          4103 => x"11",
          4104 => x"27",
          4105 => x"08",
          4106 => x"b8",
          4107 => x"55",
          4108 => x"2b",
          4109 => x"94",
          4110 => x"ff",
          4111 => x"fd",
          4112 => x"55",
          4113 => x"83",
          4114 => x"55",
          4115 => x"9c",
          4116 => x"b8",
          4117 => x"38",
          4118 => x"83",
          4119 => x"b9",
          4120 => x"16",
          4121 => x"7f",
          4122 => x"70",
          4123 => x"58",
          4124 => x"75",
          4125 => x"39",
          4126 => x"74",
          4127 => x"e0",
          4128 => x"3d",
          4129 => x"70",
          4130 => x"98",
          4131 => x"80",
          4132 => x"70",
          4133 => x"2e",
          4134 => x"78",
          4135 => x"98",
          4136 => x"d8",
          4137 => x"a0",
          4138 => x"88",
          4139 => x"51",
          4140 => x"9c",
          4141 => x"88",
          4142 => x"b7",
          4143 => x"ff",
          4144 => x"83",
          4145 => x"3f",
          4146 => x"81",
          4147 => x"34",
          4148 => x"0d",
          4149 => x"54",
          4150 => x"53",
          4151 => x"3d",
          4152 => x"3f",
          4153 => x"98",
          4154 => x"74",
          4155 => x"3d",
          4156 => x"51",
          4157 => x"82",
          4158 => x"e0",
          4159 => x"52",
          4160 => x"0d",
          4161 => x"3d",
          4162 => x"e6",
          4163 => x"e0",
          4164 => x"64",
          4165 => x"e8",
          4166 => x"e0",
          4167 => x"05",
          4168 => x"80",
          4169 => x"0c",
          4170 => x"70",
          4171 => x"56",
          4172 => x"53",
          4173 => x"e0",
          4174 => x"82",
          4175 => x"06",
          4176 => x"98",
          4177 => x"3d",
          4178 => x"3d",
          4179 => x"53",
          4180 => x"80",
          4181 => x"e0",
          4182 => x"83",
          4183 => x"7a",
          4184 => x"0c",
          4185 => x"73",
          4186 => x"80",
          4187 => x"3f",
          4188 => x"98",
          4189 => x"08",
          4190 => x"82",
          4191 => x"08",
          4192 => x"52",
          4193 => x"98",
          4194 => x"74",
          4195 => x"08",
          4196 => x"38",
          4197 => x"82",
          4198 => x"08",
          4199 => x"7b",
          4200 => x"98",
          4201 => x"51",
          4202 => x"57",
          4203 => x"38",
          4204 => x"38",
          4205 => x"ea",
          4206 => x"52",
          4207 => x"3d",
          4208 => x"5a",
          4209 => x"80",
          4210 => x"70",
          4211 => x"81",
          4212 => x"38",
          4213 => x"82",
          4214 => x"08",
          4215 => x"55",
          4216 => x"38",
          4217 => x"55",
          4218 => x"77",
          4219 => x"ff",
          4220 => x"58",
          4221 => x"f4",
          4222 => x"05",
          4223 => x"56",
          4224 => x"16",
          4225 => x"73",
          4226 => x"26",
          4227 => x"91",
          4228 => x"70",
          4229 => x"ec",
          4230 => x"34",
          4231 => x"38",
          4232 => x"08",
          4233 => x"7a",
          4234 => x"26",
          4235 => x"e0",
          4236 => x"f7",
          4237 => x"05",
          4238 => x"3f",
          4239 => x"98",
          4240 => x"53",
          4241 => x"54",
          4242 => x"33",
          4243 => x"54",
          4244 => x"15",
          4245 => x"58",
          4246 => x"8a",
          4247 => x"53",
          4248 => x"ff",
          4249 => x"e0",
          4250 => x"53",
          4251 => x"e0",
          4252 => x"30",
          4253 => x"77",
          4254 => x"51",
          4255 => x"73",
          4256 => x"bb",
          4257 => x"82",
          4258 => x"38",
          4259 => x"9e",
          4260 => x"0c",
          4261 => x"81",
          4262 => x"38",
          4263 => x"94",
          4264 => x"2a",
          4265 => x"72",
          4266 => x"51",
          4267 => x"08",
          4268 => x"82",
          4269 => x"52",
          4270 => x"e0",
          4271 => x"38",
          4272 => x"73",
          4273 => x"98",
          4274 => x"08",
          4275 => x"06",
          4276 => x"52",
          4277 => x"e0",
          4278 => x"16",
          4279 => x"0b",
          4280 => x"75",
          4281 => x"58",
          4282 => x"74",
          4283 => x"90",
          4284 => x"90",
          4285 => x"72",
          4286 => x"08",
          4287 => x"80",
          4288 => x"3d",
          4289 => x"89",
          4290 => x"80",
          4291 => x"3d",
          4292 => x"e0",
          4293 => x"80",
          4294 => x"75",
          4295 => x"08",
          4296 => x"38",
          4297 => x"57",
          4298 => x"33",
          4299 => x"55",
          4300 => x"16",
          4301 => x"82",
          4302 => x"54",
          4303 => x"52",
          4304 => x"e0",
          4305 => x"81",
          4306 => x"74",
          4307 => x"74",
          4308 => x"3d",
          4309 => x"3d",
          4310 => x"bb",
          4311 => x"82",
          4312 => x"0d",
          4313 => x"3d",
          4314 => x"e7",
          4315 => x"82",
          4316 => x"94",
          4317 => x"51",
          4318 => x"08",
          4319 => x"08",
          4320 => x"e0",
          4321 => x"84",
          4322 => x"53",
          4323 => x"38",
          4324 => x"72",
          4325 => x"82",
          4326 => x"70",
          4327 => x"98",
          4328 => x"82",
          4329 => x"ed",
          4330 => x"3d",
          4331 => x"9e",
          4332 => x"e0",
          4333 => x"51",
          4334 => x"55",
          4335 => x"80",
          4336 => x"58",
          4337 => x"8d",
          4338 => x"52",
          4339 => x"e0",
          4340 => x"3d",
          4341 => x"92",
          4342 => x"dd",
          4343 => x"82",
          4344 => x"74",
          4345 => x"11",
          4346 => x"75",
          4347 => x"81",
          4348 => x"82",
          4349 => x"08",
          4350 => x"09",
          4351 => x"5f",
          4352 => x"51",
          4353 => x"08",
          4354 => x"08",
          4355 => x"08",
          4356 => x"80",
          4357 => x"59",
          4358 => x"c9",
          4359 => x"82",
          4360 => x"38",
          4361 => x"ff",
          4362 => x"5b",
          4363 => x"7c",
          4364 => x"52",
          4365 => x"06",
          4366 => x"8e",
          4367 => x"ff",
          4368 => x"82",
          4369 => x"b8",
          4370 => x"e0",
          4371 => x"70",
          4372 => x"51",
          4373 => x"56",
          4374 => x"7c",
          4375 => x"81",
          4376 => x"7a",
          4377 => x"04",
          4378 => x"05",
          4379 => x"82",
          4380 => x"08",
          4381 => x"75",
          4382 => x"81",
          4383 => x"87",
          4384 => x"94",
          4385 => x"27",
          4386 => x"e0",
          4387 => x"76",
          4388 => x"98",
          4389 => x"ca",
          4390 => x"ff",
          4391 => x"ff",
          4392 => x"56",
          4393 => x"81",
          4394 => x"75",
          4395 => x"08",
          4396 => x"17",
          4397 => x"76",
          4398 => x"98",
          4399 => x"0c",
          4400 => x"73",
          4401 => x"38",
          4402 => x"82",
          4403 => x"e0",
          4404 => x"9c",
          4405 => x"3f",
          4406 => x"98",
          4407 => x"3d",
          4408 => x"cd",
          4409 => x"82",
          4410 => x"80",
          4411 => x"81",
          4412 => x"81",
          4413 => x"74",
          4414 => x"05",
          4415 => x"55",
          4416 => x"51",
          4417 => x"08",
          4418 => x"55",
          4419 => x"78",
          4420 => x"08",
          4421 => x"e0",
          4422 => x"70",
          4423 => x"e0",
          4424 => x"80",
          4425 => x"73",
          4426 => x"98",
          4427 => x"38",
          4428 => x"98",
          4429 => x"98",
          4430 => x"ab",
          4431 => x"98",
          4432 => x"07",
          4433 => x"2e",
          4434 => x"80",
          4435 => x"90",
          4436 => x"8c",
          4437 => x"82",
          4438 => x"98",
          4439 => x"0d",
          4440 => x"52",
          4441 => x"e0",
          4442 => x"82",
          4443 => x"3d",
          4444 => x"e0",
          4445 => x"86",
          4446 => x"e0",
          4447 => x"82",
          4448 => x"70",
          4449 => x"54",
          4450 => x"52",
          4451 => x"bc",
          4452 => x"56",
          4453 => x"54",
          4454 => x"81",
          4455 => x"98",
          4456 => x"38",
          4457 => x"b6",
          4458 => x"51",
          4459 => x"08",
          4460 => x"38",
          4461 => x"ff",
          4462 => x"b8",
          4463 => x"c3",
          4464 => x"80",
          4465 => x"75",
          4466 => x"b7",
          4467 => x"53",
          4468 => x"3f",
          4469 => x"34",
          4470 => x"51",
          4471 => x"0b",
          4472 => x"89",
          4473 => x"e0",
          4474 => x"0a",
          4475 => x"86",
          4476 => x"ff",
          4477 => x"8b",
          4478 => x"15",
          4479 => x"82",
          4480 => x"53",
          4481 => x"3f",
          4482 => x"0d",
          4483 => x"05",
          4484 => x"3d",
          4485 => x"d4",
          4486 => x"82",
          4487 => x"4e",
          4488 => x"52",
          4489 => x"08",
          4490 => x"38",
          4491 => x"06",
          4492 => x"a0",
          4493 => x"ff",
          4494 => x"b0",
          4495 => x"54",
          4496 => x"52",
          4497 => x"98",
          4498 => x"38",
          4499 => x"06",
          4500 => x"92",
          4501 => x"e0",
          4502 => x"81",
          4503 => x"3f",
          4504 => x"98",
          4505 => x"53",
          4506 => x"16",
          4507 => x"05",
          4508 => x"70",
          4509 => x"55",
          4510 => x"73",
          4511 => x"83",
          4512 => x"2a",
          4513 => x"80",
          4514 => x"80",
          4515 => x"b4",
          4516 => x"78",
          4517 => x"82",
          4518 => x"38",
          4519 => x"ff",
          4520 => x"79",
          4521 => x"e0",
          4522 => x"33",
          4523 => x"9a",
          4524 => x"ff",
          4525 => x"83",
          4526 => x"08",
          4527 => x"82",
          4528 => x"08",
          4529 => x"3f",
          4530 => x"e0",
          4531 => x"3d",
          4532 => x"84",
          4533 => x"82",
          4534 => x"3d",
          4535 => x"08",
          4536 => x"38",
          4537 => x"05",
          4538 => x"08",
          4539 => x"02",
          4540 => x"54",
          4541 => x"06",
          4542 => x"06",
          4543 => x"56",
          4544 => x"0b",
          4545 => x"97",
          4546 => x"82",
          4547 => x"ee",
          4548 => x"3d",
          4549 => x"ce",
          4550 => x"e0",
          4551 => x"64",
          4552 => x"d0",
          4553 => x"e0",
          4554 => x"05",
          4555 => x"73",
          4556 => x"22",
          4557 => x"1f",
          4558 => x"81",
          4559 => x"a1",
          4560 => x"74",
          4561 => x"04",
          4562 => x"80",
          4563 => x"3d",
          4564 => x"08",
          4565 => x"e0",
          4566 => x"57",
          4567 => x"70",
          4568 => x"80",
          4569 => x"52",
          4570 => x"97",
          4571 => x"e0",
          4572 => x"73",
          4573 => x"98",
          4574 => x"38",
          4575 => x"08",
          4576 => x"19",
          4577 => x"74",
          4578 => x"ec",
          4579 => x"74",
          4580 => x"16",
          4581 => x"73",
          4582 => x"84",
          4583 => x"7a",
          4584 => x"07",
          4585 => x"80",
          4586 => x"7b",
          4587 => x"80",
          4588 => x"e0",
          4589 => x"55",
          4590 => x"8b",
          4591 => x"83",
          4592 => x"51",
          4593 => x"08",
          4594 => x"99",
          4595 => x"53",
          4596 => x"3d",
          4597 => x"08",
          4598 => x"e0",
          4599 => x"a0",
          4600 => x"9b",
          4601 => x"55",
          4602 => x"77",
          4603 => x"3f",
          4604 => x"26",
          4605 => x"51",
          4606 => x"e0",
          4607 => x"e0",
          4608 => x"74",
          4609 => x"d3",
          4610 => x"e0",
          4611 => x"27",
          4612 => x"8b",
          4613 => x"55",
          4614 => x"8f",
          4615 => x"70",
          4616 => x"74",
          4617 => x"16",
          4618 => x"9f",
          4619 => x"54",
          4620 => x"b1",
          4621 => x"a3",
          4622 => x"54",
          4623 => x"38",
          4624 => x"40",
          4625 => x"52",
          4626 => x"98",
          4627 => x"f7",
          4628 => x"bc",
          4629 => x"e0",
          4630 => x"38",
          4631 => x"39",
          4632 => x"81",
          4633 => x"74",
          4634 => x"51",
          4635 => x"08",
          4636 => x"a0",
          4637 => x"51",
          4638 => x"0b",
          4639 => x"66",
          4640 => x"81",
          4641 => x"9c",
          4642 => x"73",
          4643 => x"3d",
          4644 => x"02",
          4645 => x"3d",
          4646 => x"5a",
          4647 => x"58",
          4648 => x"91",
          4649 => x"7c",
          4650 => x"59",
          4651 => x"81",
          4652 => x"73",
          4653 => x"82",
          4654 => x"8b",
          4655 => x"2b",
          4656 => x"fe",
          4657 => x"70",
          4658 => x"e0",
          4659 => x"40",
          4660 => x"88",
          4661 => x"38",
          4662 => x"56",
          4663 => x"3f",
          4664 => x"08",
          4665 => x"e0",
          4666 => x"82",
          4667 => x"38",
          4668 => x"16",
          4669 => x"87",
          4670 => x"74",
          4671 => x"38",
          4672 => x"2e",
          4673 => x"80",
          4674 => x"81",
          4675 => x"56",
          4676 => x"9d",
          4677 => x"82",
          4678 => x"81",
          4679 => x"d3",
          4680 => x"7c",
          4681 => x"b3",
          4682 => x"1b",
          4683 => x"54",
          4684 => x"fe",
          4685 => x"74",
          4686 => x"16",
          4687 => x"73",
          4688 => x"e0",
          4689 => x"3d",
          4690 => x"ef",
          4691 => x"59",
          4692 => x"82",
          4693 => x"82",
          4694 => x"e0",
          4695 => x"2e",
          4696 => x"98",
          4697 => x"e0",
          4698 => x"33",
          4699 => x"ff",
          4700 => x"81",
          4701 => x"83",
          4702 => x"2a",
          4703 => x"74",
          4704 => x"53",
          4705 => x"3f",
          4706 => x"55",
          4707 => x"80",
          4708 => x"06",
          4709 => x"49",
          4710 => x"79",
          4711 => x"26",
          4712 => x"74",
          4713 => x"fe",
          4714 => x"70",
          4715 => x"7a",
          4716 => x"80",
          4717 => x"74",
          4718 => x"e0",
          4719 => x"7f",
          4720 => x"82",
          4721 => x"fe",
          4722 => x"e0",
          4723 => x"8e",
          4724 => x"81",
          4725 => x"1b",
          4726 => x"80",
          4727 => x"51",
          4728 => x"08",
          4729 => x"cd",
          4730 => x"39",
          4731 => x"7f",
          4732 => x"82",
          4733 => x"83",
          4734 => x"08",
          4735 => x"5f",
          4736 => x"8a",
          4737 => x"56",
          4738 => x"93",
          4739 => x"38",
          4740 => x"44",
          4741 => x"06",
          4742 => x"62",
          4743 => x"83",
          4744 => x"82",
          4745 => x"78",
          4746 => x"80",
          4747 => x"2a",
          4748 => x"56",
          4749 => x"77",
          4750 => x"79",
          4751 => x"5a",
          4752 => x"27",
          4753 => x"9c",
          4754 => x"29",
          4755 => x"55",
          4756 => x"08",
          4757 => x"ff",
          4758 => x"89",
          4759 => x"2a",
          4760 => x"56",
          4761 => x"77",
          4762 => x"79",
          4763 => x"5a",
          4764 => x"27",
          4765 => x"9b",
          4766 => x"84",
          4767 => x"f5",
          4768 => x"98",
          4769 => x"71",
          4770 => x"5e",
          4771 => x"5c",
          4772 => x"05",
          4773 => x"70",
          4774 => x"57",
          4775 => x"06",
          4776 => x"5c",
          4777 => x"29",
          4778 => x"55",
          4779 => x"7c",
          4780 => x"31",
          4781 => x"e0",
          4782 => x"81",
          4783 => x"83",
          4784 => x"87",
          4785 => x"fd",
          4786 => x"2e",
          4787 => x"ff",
          4788 => x"a0",
          4789 => x"74",
          4790 => x"fd",
          4791 => x"80",
          4792 => x"39",
          4793 => x"92",
          4794 => x"59",
          4795 => x"86",
          4796 => x"09",
          4797 => x"f5",
          4798 => x"55",
          4799 => x"80",
          4800 => x"b0",
          4801 => x"7a",
          4802 => x"52",
          4803 => x"79",
          4804 => x"06",
          4805 => x"3f",
          4806 => x"32",
          4807 => x"06",
          4808 => x"8d",
          4809 => x"ff",
          4810 => x"06",
          4811 => x"3f",
          4812 => x"ff",
          4813 => x"34",
          4814 => x"d0",
          4815 => x"ff",
          4816 => x"51",
          4817 => x"09",
          4818 => x"b2",
          4819 => x"8d",
          4820 => x"ff",
          4821 => x"51",
          4822 => x"1b",
          4823 => x"b2",
          4824 => x"80",
          4825 => x"80",
          4826 => x"f0",
          4827 => x"82",
          4828 => x"ff",
          4829 => x"06",
          4830 => x"3f",
          4831 => x"0b",
          4832 => x"84",
          4833 => x"3f",
          4834 => x"70",
          4835 => x"54",
          4836 => x"88",
          4837 => x"08",
          4838 => x"81",
          4839 => x"1f",
          4840 => x"af",
          4841 => x"51",
          4842 => x"a4",
          4843 => x"3f",
          4844 => x"e4",
          4845 => x"18",
          4846 => x"ee",
          4847 => x"ff",
          4848 => x"78",
          4849 => x"87",
          4850 => x"87",
          4851 => x"7a",
          4852 => x"66",
          4853 => x"88",
          4854 => x"2e",
          4855 => x"7a",
          4856 => x"84",
          4857 => x"0a",
          4858 => x"ff",
          4859 => x"38",
          4860 => x"8a",
          4861 => x"62",
          4862 => x"75",
          4863 => x"f7",
          4864 => x"38",
          4865 => x"52",
          4866 => x"16",
          4867 => x"38",
          4868 => x"8d",
          4869 => x"38",
          4870 => x"83",
          4871 => x"7a",
          4872 => x"82",
          4873 => x"16",
          4874 => x"38",
          4875 => x"86",
          4876 => x"38",
          4877 => x"81",
          4878 => x"54",
          4879 => x"84",
          4880 => x"08",
          4881 => x"55",
          4882 => x"82",
          4883 => x"51",
          4884 => x"62",
          4885 => x"fd",
          4886 => x"51",
          4887 => x"52",
          4888 => x"be",
          4889 => x"81",
          4890 => x"77",
          4891 => x"67",
          4892 => x"51",
          4893 => x"16",
          4894 => x"bf",
          4895 => x"e0",
          4896 => x"83",
          4897 => x"67",
          4898 => x"ce",
          4899 => x"7f",
          4900 => x"82",
          4901 => x"80",
          4902 => x"81",
          4903 => x"89",
          4904 => x"86",
          4905 => x"82",
          4906 => x"f5",
          4907 => x"79",
          4908 => x"78",
          4909 => x"55",
          4910 => x"51",
          4911 => x"81",
          4912 => x"74",
          4913 => x"81",
          4914 => x"8a",
          4915 => x"76",
          4916 => x"55",
          4917 => x"0d",
          4918 => x"05",
          4919 => x"2e",
          4920 => x"76",
          4921 => x"80",
          4922 => x"77",
          4923 => x"34",
          4924 => x"38",
          4925 => x"8c",
          4926 => x"3f",
          4927 => x"07",
          4928 => x"56",
          4929 => x"18",
          4930 => x"0d",
          4931 => x"75",
          4932 => x"54",
          4933 => x"51",
          4934 => x"91",
          4935 => x"81",
          4936 => x"83",
          4937 => x"0c",
          4938 => x"75",
          4939 => x"51",
          4940 => x"85",
          4941 => x"80",
          4942 => x"70",
          4943 => x"72",
          4944 => x"8d",
          4945 => x"0d",
          4946 => x"55",
          4947 => x"8a",
          4948 => x"80",
          4949 => x"51",
          4950 => x"b4",
          4951 => x"d3",
          4952 => x"38",
          4953 => x"53",
          4954 => x"71",
          4955 => x"51",
          4956 => x"81",
          4957 => x"98",
          4958 => x"0d",
          4959 => x"96",
          4960 => x"80",
          4961 => x"39",
          4962 => x"91",
          4963 => x"70",
          4964 => x"54",
          4965 => x"3d",
          4966 => x"70",
          4967 => x"70",
          4968 => x"57",
          4969 => x"82",
          4970 => x"57",
          4971 => x"75",
          4972 => x"fb",
          4973 => x"70",
          4974 => x"18",
          4975 => x"80",
          4976 => x"38",
          4977 => x"51",
          4978 => x"76",
          4979 => x"c3",
          4980 => x"71",
          4981 => x"51",
          4982 => x"d0",
          4983 => x"90",
          4984 => x"b0",
          4985 => x"51",
          4986 => x"39",
          4987 => x"56",
          4988 => x"e0",
          4989 => x"ff",
          4990 => x"ff",
          4991 => x"00",
          4992 => x"00",
          4993 => x"00",
          4994 => x"00",
          4995 => x"00",
          4996 => x"00",
          4997 => x"00",
          4998 => x"00",
          4999 => x"00",
          5000 => x"00",
          5001 => x"00",
          5002 => x"00",
          5003 => x"00",
          5004 => x"00",
          5005 => x"00",
          5006 => x"00",
          5007 => x"00",
          5008 => x"00",
          5009 => x"00",
          5010 => x"00",
          5011 => x"00",
          5012 => x"00",
          5013 => x"00",
          5014 => x"00",
          5015 => x"00",
          5016 => x"00",
          5017 => x"00",
          5018 => x"00",
          5019 => x"00",
          5020 => x"00",
          5021 => x"00",
          5022 => x"00",
          5023 => x"00",
          5024 => x"00",
          5025 => x"00",
          5026 => x"00",
          5027 => x"00",
          5028 => x"00",
          5029 => x"00",
          5030 => x"00",
          5031 => x"00",
          5032 => x"00",
          5033 => x"00",
          5034 => x"00",
          5035 => x"00",
          5036 => x"00",
          5037 => x"00",
          5038 => x"00",
          5039 => x"00",
          5040 => x"00",
          5041 => x"00",
          5042 => x"00",
          5043 => x"00",
          5044 => x"00",
          5045 => x"00",
          5046 => x"00",
          5047 => x"00",
          5048 => x"00",
          5049 => x"00",
          5050 => x"00",
          5051 => x"00",
          5052 => x"00",
          5053 => x"00",
          5054 => x"00",
          5055 => x"00",
          5056 => x"00",
          5057 => x"00",
          5058 => x"00",
          5059 => x"00",
          5060 => x"00",
          5061 => x"00",
          5062 => x"00",
          5063 => x"00",
          5064 => x"00",
          5065 => x"6c",
          5066 => x"00",
          5067 => x"00",
          5068 => x"00",
          5069 => x"72",
          5070 => x"00",
          5071 => x"00",
          5072 => x"00",
          5073 => x"65",
          5074 => x"69",
          5075 => x"66",
          5076 => x"61",
          5077 => x"6d",
          5078 => x"72",
          5079 => x"00",
          5080 => x"00",
          5081 => x"63",
          5082 => x"63",
          5083 => x"00",
          5084 => x"69",
          5085 => x"72",
          5086 => x"6e",
          5087 => x"72",
          5088 => x"6e",
          5089 => x"79",
          5090 => x"6c",
          5091 => x"2e",
          5092 => x"74",
          5093 => x"2e",
          5094 => x"69",
          5095 => x"61",
          5096 => x"63",
          5097 => x"6e",
          5098 => x"69",
          5099 => x"61",
          5100 => x"74",
          5101 => x"69",
          5102 => x"6c",
          5103 => x"69",
          5104 => x"44",
          5105 => x"74",
          5106 => x"63",
          5107 => x"72",
          5108 => x"62",
          5109 => x"6e",
          5110 => x"00",
          5111 => x"6e",
          5112 => x"6c",
          5113 => x"6f",
          5114 => x"69",
          5115 => x"65",
          5116 => x"66",
          5117 => x"20",
          5118 => x"6f",
          5119 => x"6f",
          5120 => x"69",
          5121 => x"6f",
          5122 => x"6e",
          5123 => x"6c",
          5124 => x"69",
          5125 => x"6f",
          5126 => x"6e",
          5127 => x"65",
          5128 => x"72",
          5129 => x"6f",
          5130 => x"6f",
          5131 => x"65",
          5132 => x"61",
          5133 => x"73",
          5134 => x"65",
          5135 => x"75",
          5136 => x"00",
          5137 => x"77",
          5138 => x"2e",
          5139 => x"62",
          5140 => x"20",
          5141 => x"62",
          5142 => x"63",
          5143 => x"65",
          5144 => x"30",
          5145 => x"20",
          5146 => x"00",
          5147 => x"20",
          5148 => x"30",
          5149 => x"20",
          5150 => x"00",
          5151 => x"2a",
          5152 => x"31",
          5153 => x"30",
          5154 => x"00",
          5155 => x"20",
          5156 => x"78",
          5157 => x"20",
          5158 => x"50",
          5159 => x"72",
          5160 => x"64",
          5161 => x"69",
          5162 => x"65",
          5163 => x"53",
          5164 => x"72",
          5165 => x"4f",
          5166 => x"69",
          5167 => x"74",
          5168 => x"20",
          5169 => x"72",
          5170 => x"41",
          5171 => x"69",
          5172 => x"74",
          5173 => x"20",
          5174 => x"72",
          5175 => x"41",
          5176 => x"69",
          5177 => x"74",
          5178 => x"20",
          5179 => x"72",
          5180 => x"65",
          5181 => x"70",
          5182 => x"2e",
          5183 => x"69",
          5184 => x"72",
          5185 => x"75",
          5186 => x"62",
          5187 => x"4f",
          5188 => x"73",
          5189 => x"61",
          5190 => x"20",
          5191 => x"69",
          5192 => x"61",
          5193 => x"6c",
          5194 => x"69",
          5195 => x"6c",
          5196 => x"20",
          5197 => x"69",
          5198 => x"00",
          5199 => x"6e",
          5200 => x"6f",
          5201 => x"2e",
          5202 => x"30",
          5203 => x"78",
          5204 => x"78",
          5205 => x"00",
          5206 => x"4d",
          5207 => x"43",
          5208 => x"2e",
          5209 => x"20",
          5210 => x"3f",
          5211 => x"20",
          5212 => x"30",
          5213 => x"6c",
          5214 => x"78",
          5215 => x"20",
          5216 => x"25",
          5217 => x"2e",
          5218 => x"6e",
          5219 => x"40",
          5220 => x"2e",
          5221 => x"61",
          5222 => x"72",
          5223 => x"65",
          5224 => x"00",
          5225 => x"72",
          5226 => x"70",
          5227 => x"6e",
          5228 => x"6f",
          5229 => x"6f",
          5230 => x"00",
          5231 => x"69",
          5232 => x"73",
          5233 => x"00",
          5234 => x"73",
          5235 => x"64",
          5236 => x"61",
          5237 => x"6e",
          5238 => x"65",
          5239 => x"68",
          5240 => x"20",
          5241 => x"70",
          5242 => x"63",
          5243 => x"00",
          5244 => x"6e",
          5245 => x"6e",
          5246 => x"69",
          5247 => x"74",
          5248 => x"64",
          5249 => x"25",
          5250 => x"2e",
          5251 => x"6f",
          5252 => x"67",
          5253 => x"00",
          5254 => x"6d",
          5255 => x"6e",
          5256 => x"0a",
          5257 => x"20",
          5258 => x"6e",
          5259 => x"20",
          5260 => x"52",
          5261 => x"38",
          5262 => x"2e",
          5263 => x"44",
          5264 => x"20",
          5265 => x"30",
          5266 => x"20",
          5267 => x"42",
          5268 => x"38",
          5269 => x"2e",
          5270 => x"52",
          5271 => x"20",
          5272 => x"30",
          5273 => x"20",
          5274 => x"20",
          5275 => x"38",
          5276 => x"2e",
          5277 => x"44",
          5278 => x"20",
          5279 => x"73",
          5280 => x"2e",
          5281 => x"49",
          5282 => x"20",
          5283 => x"20",
          5284 => x"2e",
          5285 => x"4e",
          5286 => x"20",
          5287 => x"6c",
          5288 => x"2e",
          5289 => x"49",
          5290 => x"42",
          5291 => x"20",
          5292 => x"43",
          5293 => x"4f",
          5294 => x"20",
          5295 => x"20",
          5296 => x"64",
          5297 => x"3a",
          5298 => x"50",
          5299 => x"20",
          5300 => x"41",
          5301 => x"3d",
          5302 => x"00",
          5303 => x"50",
          5304 => x"79",
          5305 => x"41",
          5306 => x"3d",
          5307 => x"00",
          5308 => x"74",
          5309 => x"72",
          5310 => x"73",
          5311 => x"3d",
          5312 => x"00",
          5313 => x"00",
          5314 => x"50",
          5315 => x"20",
          5316 => x"20",
          5317 => x"3d",
          5318 => x"00",
          5319 => x"79",
          5320 => x"6f",
          5321 => x"20",
          5322 => x"3d",
          5323 => x"64",
          5324 => x"20",
          5325 => x"20",
          5326 => x"72",
          5327 => x"20",
          5328 => x"2e",
          5329 => x"0a",
          5330 => x"69",
          5331 => x"53",
          5332 => x"6f",
          5333 => x"3d",
          5334 => x"64",
          5335 => x"6d",
          5336 => x"65",
          5337 => x"6c",
          5338 => x"56",
          5339 => x"00",
          5340 => x"77",
          5341 => x"00",
          5342 => x"00",
          5343 => x"00",
          5344 => x"00",
          5345 => x"00",
          5346 => x"00",
          5347 => x"00",
          5348 => x"00",
          5349 => x"00",
          5350 => x"00",
          5351 => x"00",
          5352 => x"00",
          5353 => x"00",
          5354 => x"00",
          5355 => x"00",
          5356 => x"00",
          5357 => x"00",
          5358 => x"00",
          5359 => x"00",
          5360 => x"00",
          5361 => x"00",
          5362 => x"00",
          5363 => x"00",
          5364 => x"00",
          5365 => x"00",
          5366 => x"00",
          5367 => x"00",
          5368 => x"00",
          5369 => x"00",
          5370 => x"00",
          5371 => x"00",
          5372 => x"00",
          5373 => x"00",
          5374 => x"5b",
          5375 => x"5b",
          5376 => x"5b",
          5377 => x"30",
          5378 => x"5b",
          5379 => x"00",
          5380 => x"00",
          5381 => x"00",
          5382 => x"00",
          5383 => x"00",
          5384 => x"00",
          5385 => x"72",
          5386 => x"00",
          5387 => x"30",
          5388 => x"0a",
          5389 => x"64",
          5390 => x"65",
          5391 => x"69",
          5392 => x"69",
          5393 => x"4f",
          5394 => x"61",
          5395 => x"65",
          5396 => x"65",
          5397 => x"79",
          5398 => x"64",
          5399 => x"67",
          5400 => x"2a",
          5401 => x"00",
          5402 => x"5d",
          5403 => x"41",
          5404 => x"fe",
          5405 => x"2e",
          5406 => x"4d",
          5407 => x"54",
          5408 => x"4f",
          5409 => x"20",
          5410 => x"20",
          5411 => x"00",
          5412 => x"00",
          5413 => x"0e",
          5414 => x"00",
          5415 => x"41",
          5416 => x"49",
          5417 => x"4f",
          5418 => x"9d",
          5419 => x"a5",
          5420 => x"ad",
          5421 => x"b5",
          5422 => x"bd",
          5423 => x"c5",
          5424 => x"cd",
          5425 => x"d5",
          5426 => x"dd",
          5427 => x"e5",
          5428 => x"ed",
          5429 => x"f5",
          5430 => x"fd",
          5431 => x"5b",
          5432 => x"3e",
          5433 => x"01",
          5434 => x"00",
          5435 => x"01",
          5436 => x"10",
          5437 => x"c7",
          5438 => x"e4",
          5439 => x"ea",
          5440 => x"ee",
          5441 => x"c9",
          5442 => x"f6",
          5443 => x"ff",
          5444 => x"a3",
          5445 => x"e1",
          5446 => x"f1",
          5447 => x"bf",
          5448 => x"bc",
          5449 => x"91",
          5450 => x"24",
          5451 => x"55",
          5452 => x"5d",
          5453 => x"14",
          5454 => x"00",
          5455 => x"5a",
          5456 => x"60",
          5457 => x"68",
          5458 => x"58",
          5459 => x"6a",
          5460 => x"84",
          5461 => x"b1",
          5462 => x"a3",
          5463 => x"a6",
          5464 => x"1e",
          5465 => x"61",
          5466 => x"20",
          5467 => x"b0",
          5468 => x"7f",
          5469 => x"61",
          5470 => x"f8",
          5471 => x"78",
          5472 => x"06",
          5473 => x"2e",
          5474 => x"4d",
          5475 => x"82",
          5476 => x"87",
          5477 => x"8b",
          5478 => x"8f",
          5479 => x"93",
          5480 => x"97",
          5481 => x"9b",
          5482 => x"9f",
          5483 => x"a2",
          5484 => x"a7",
          5485 => x"ab",
          5486 => x"af",
          5487 => x"b3",
          5488 => x"b7",
          5489 => x"bb",
          5490 => x"f7",
          5491 => x"c3",
          5492 => x"c7",
          5493 => x"cb",
          5494 => x"dd",
          5495 => x"12",
          5496 => x"f4",
          5497 => x"22",
          5498 => x"65",
          5499 => x"66",
          5500 => x"41",
          5501 => x"40",
          5502 => x"89",
          5503 => x"5a",
          5504 => x"5e",
          5505 => x"62",
          5506 => x"66",
          5507 => x"6a",
          5508 => x"6e",
          5509 => x"9d",
          5510 => x"76",
          5511 => x"7a",
          5512 => x"7e",
          5513 => x"82",
          5514 => x"86",
          5515 => x"b1",
          5516 => x"8e",
          5517 => x"b7",
          5518 => x"fe",
          5519 => x"86",
          5520 => x"b1",
          5521 => x"a3",
          5522 => x"cc",
          5523 => x"8f",
          5524 => x"0a",
          5525 => x"f5",
          5526 => x"f9",
          5527 => x"20",
          5528 => x"22",
          5529 => x"0e",
          5530 => x"d0",
          5531 => x"00",
          5532 => x"63",
          5533 => x"5a",
          5534 => x"06",
          5535 => x"08",
          5536 => x"07",
          5537 => x"54",
          5538 => x"60",
          5539 => x"ba",
          5540 => x"ca",
          5541 => x"f8",
          5542 => x"fa",
          5543 => x"90",
          5544 => x"b0",
          5545 => x"b2",
          5546 => x"c3",
          5547 => x"02",
          5548 => x"f3",
          5549 => x"01",
          5550 => x"84",
          5551 => x"1a",
          5552 => x"02",
          5553 => x"02",
          5554 => x"26",
          5555 => x"00",
          5556 => x"02",
          5557 => x"00",
          5558 => x"04",
          5559 => x"00",
          5560 => x"14",
          5561 => x"00",
          5562 => x"2b",
          5563 => x"00",
          5564 => x"30",
          5565 => x"00",
          5566 => x"3c",
          5567 => x"00",
          5568 => x"3d",
          5569 => x"00",
          5570 => x"3f",
          5571 => x"00",
          5572 => x"40",
          5573 => x"00",
          5574 => x"41",
          5575 => x"00",
          5576 => x"42",
          5577 => x"00",
          5578 => x"43",
          5579 => x"00",
          5580 => x"50",
          5581 => x"00",
          5582 => x"51",
          5583 => x"00",
          5584 => x"54",
          5585 => x"00",
          5586 => x"55",
          5587 => x"00",
          5588 => x"79",
          5589 => x"00",
          5590 => x"78",
          5591 => x"00",
          5592 => x"82",
          5593 => x"00",
          5594 => x"83",
          5595 => x"00",
          5596 => x"85",
          5597 => x"00",
          5598 => x"8c",
          5599 => x"00",
          5600 => x"8d",
          5601 => x"00",
          5602 => x"8e",
          5603 => x"00",
          5604 => x"8f",
          5605 => x"00",
          5606 => x"00",
          5607 => x"00",
          5608 => x"01",
          5609 => x"01",
          5610 => x"00",
          5611 => x"00",
          5612 => x"00",
          5613 => x"f5",
          5614 => x"f5",
          5615 => x"01",
          5616 => x"01",
          5617 => x"00",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"00",
          5630 => x"00",
          5631 => x"00",
          5632 => x"00",
          5633 => x"01",
          5634 => x"00",
        others => X"00"
    );

    shared variable RAM7 : ramArray :=
    (
             0 => x"f8",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"90",
             5 => x"8c",
             6 => x"00",
             7 => x"00",
             8 => x"72",
             9 => x"83",
            10 => x"04",
            11 => x"00",
            12 => x"83",
            13 => x"05",
            14 => x"73",
            15 => x"83",
            16 => x"72",
            17 => x"73",
            18 => x"53",
            19 => x"00",
            20 => x"73",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"0a",
            26 => x"05",
            27 => x"04",
            28 => x"73",
            29 => x"00",
            30 => x"00",
            31 => x"00",
            32 => x"00",
            33 => x"00",
            34 => x"00",
            35 => x"00",
            36 => x"d1",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"0a",
            41 => x"00",
            42 => x"00",
            43 => x"00",
            44 => x"09",
            45 => x"05",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"81",
            50 => x"04",
            51 => x"00",
            52 => x"04",
            53 => x"82",
            54 => x"fc",
            55 => x"00",
            56 => x"72",
            57 => x"0a",
            58 => x"00",
            59 => x"00",
            60 => x"72",
            61 => x"0a",
            62 => x"00",
            63 => x"00",
            64 => x"52",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"05",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"73",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"72",
            77 => x"10",
            78 => x"04",
            79 => x"00",
            80 => x"0b",
            81 => x"10",
            82 => x"93",
            83 => x"00",
            84 => x"90",
            85 => x"fe",
            86 => x"0c",
            87 => x"00",
            88 => x"90",
            89 => x"fc",
            90 => x"0c",
            91 => x"00",
            92 => x"05",
            93 => x"70",
            94 => x"05",
            95 => x"04",
            96 => x"05",
            97 => x"05",
            98 => x"74",
            99 => x"51",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"04",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"10",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"05",
           125 => x"ff",
           126 => x"ff",
           127 => x"ff",
           128 => x"ff",
           129 => x"ff",
           130 => x"ff",
           131 => x"ff",
           132 => x"81",
           133 => x"0b",
           134 => x"0b",
           135 => x"b6",
           136 => x"0b",
           137 => x"0b",
           138 => x"f7",
           139 => x"0b",
           140 => x"0b",
           141 => x"b8",
           142 => x"0b",
           143 => x"0b",
           144 => x"fc",
           145 => x"0b",
           146 => x"0b",
           147 => x"c0",
           148 => x"0b",
           149 => x"0b",
           150 => x"84",
           151 => x"0b",
           152 => x"0b",
           153 => x"c8",
           154 => x"0b",
           155 => x"0b",
           156 => x"8c",
           157 => x"0b",
           158 => x"0b",
           159 => x"d0",
           160 => x"0b",
           161 => x"0b",
           162 => x"94",
           163 => x"0b",
           164 => x"0b",
           165 => x"d8",
           166 => x"0b",
           167 => x"0b",
           168 => x"9c",
           169 => x"0b",
           170 => x"0b",
           171 => x"e0",
           172 => x"0b",
           173 => x"ff",
           174 => x"ff",
           175 => x"ff",
           176 => x"ff",
           177 => x"ff",
           178 => x"ff",
           179 => x"ff",
           180 => x"ff",
           181 => x"ff",
           182 => x"ff",
           183 => x"ff",
           184 => x"ff",
           185 => x"ff",
           186 => x"ff",
           187 => x"ff",
           188 => x"ff",
           189 => x"ff",
           190 => x"ff",
           191 => x"ff",
           192 => x"04",
           193 => x"2d",
           194 => x"90",
           195 => x"2d",
           196 => x"90",
           197 => x"2d",
           198 => x"90",
           199 => x"2d",
           200 => x"90",
           201 => x"2d",
           202 => x"90",
           203 => x"2d",
           204 => x"90",
           205 => x"9f",
           206 => x"80",
           207 => x"d4",
           208 => x"c0",
           209 => x"94",
           210 => x"c0",
           211 => x"96",
           212 => x"c0",
           213 => x"98",
           214 => x"c0",
           215 => x"80",
           216 => x"80",
           217 => x"0c",
           218 => x"08",
           219 => x"a4",
           220 => x"a4",
           221 => x"e0",
           222 => x"e0",
           223 => x"82",
           224 => x"82",
           225 => x"04",
           226 => x"2d",
           227 => x"90",
           228 => x"a7",
           229 => x"80",
           230 => x"fb",
           231 => x"c0",
           232 => x"81",
           233 => x"80",
           234 => x"0c",
           235 => x"08",
           236 => x"a4",
           237 => x"a4",
           238 => x"e0",
           239 => x"e0",
           240 => x"82",
           241 => x"82",
           242 => x"04",
           243 => x"2d",
           244 => x"90",
           245 => x"c7",
           246 => x"80",
           247 => x"95",
           248 => x"c0",
           249 => x"82",
           250 => x"80",
           251 => x"0c",
           252 => x"08",
           253 => x"a4",
           254 => x"a4",
           255 => x"e0",
           256 => x"e0",
           257 => x"82",
           258 => x"82",
           259 => x"04",
           260 => x"2d",
           261 => x"90",
           262 => x"e0",
           263 => x"80",
           264 => x"85",
           265 => x"c0",
           266 => x"82",
           267 => x"80",
           268 => x"0c",
           269 => x"08",
           270 => x"a4",
           271 => x"a4",
           272 => x"e0",
           273 => x"e0",
           274 => x"82",
           275 => x"82",
           276 => x"04",
           277 => x"2d",
           278 => x"90",
           279 => x"e9",
           280 => x"80",
           281 => x"b2",
           282 => x"c0",
           283 => x"81",
           284 => x"80",
           285 => x"0c",
           286 => x"08",
           287 => x"a4",
           288 => x"a4",
           289 => x"e0",
           290 => x"e0",
           291 => x"82",
           292 => x"82",
           293 => x"04",
           294 => x"2d",
           295 => x"90",
           296 => x"ef",
           297 => x"80",
           298 => x"af",
           299 => x"c0",
           300 => x"81",
           301 => x"80",
           302 => x"0c",
           303 => x"08",
           304 => x"a4",
           305 => x"a4",
           306 => x"04",
           307 => x"10",
           308 => x"10",
           309 => x"10",
           310 => x"53",
           311 => x"06",
           312 => x"05",
           313 => x"06",
           314 => x"72",
           315 => x"05",
           316 => x"53",
           317 => x"04",
           318 => x"27",
           319 => x"53",
           320 => x"8c",
           321 => x"82",
           322 => x"0c",
           323 => x"8c",
           324 => x"05",
           325 => x"08",
           326 => x"08",
           327 => x"84",
           328 => x"82",
           329 => x"e0",
           330 => x"e0",
           331 => x"82",
           332 => x"08",
           333 => x"0d",
           334 => x"85",
           335 => x"06",
           336 => x"80",
           337 => x"08",
           338 => x"82",
           339 => x"c4",
           340 => x"08",
           341 => x"05",
           342 => x"f8",
           343 => x"05",
           344 => x"0c",
           345 => x"8a",
           346 => x"e0",
           347 => x"e9",
           348 => x"08",
           349 => x"08",
           350 => x"0c",
           351 => x"08",
           352 => x"80",
           353 => x"0c",
           354 => x"fc",
           355 => x"05",
           356 => x"e0",
           357 => x"82",
           358 => x"e0",
           359 => x"82",
           360 => x"80",
           361 => x"08",
           362 => x"08",
           363 => x"08",
           364 => x"08",
           365 => x"87",
           366 => x"82",
           367 => x"0c",
           368 => x"a4",
           369 => x"08",
           370 => x"e0",
           371 => x"a4",
           372 => x"08",
           373 => x"fc",
           374 => x"05",
           375 => x"05",
           376 => x"05",
           377 => x"82",
           378 => x"08",
           379 => x"ec",
           380 => x"05",
           381 => x"82",
           382 => x"82",
           383 => x"82",
           384 => x"08",
           385 => x"0d",
           386 => x"82",
           387 => x"e0",
           388 => x"e0",
           389 => x"e0",
           390 => x"a3",
           391 => x"e0",
           392 => x"a4",
           393 => x"98",
           394 => x"e0",
           395 => x"02",
           396 => x"80",
           397 => x"23",
           398 => x"53",
           399 => x"a4",
           400 => x"70",
           401 => x"06",
           402 => x"2e",
           403 => x"08",
           404 => x"e0",
           405 => x"33",
           406 => x"05",
           407 => x"80",
           408 => x"08",
           409 => x"a4",
           410 => x"08",
           411 => x"53",
           412 => x"e0",
           413 => x"73",
           414 => x"08",
           415 => x"81",
           416 => x"05",
           417 => x"06",
           418 => x"e8",
           419 => x"2c",
           420 => x"e0",
           421 => x"2a",
           422 => x"51",
           423 => x"82",
           424 => x"82",
           425 => x"a4",
           426 => x"82",
           427 => x"98",
           428 => x"2b",
           429 => x"53",
           430 => x"08",
           431 => x"e8",
           432 => x"f8",
           433 => x"51",
           434 => x"05",
           435 => x"33",
           436 => x"51",
           437 => x"ff",
           438 => x"34",
           439 => x"70",
           440 => x"53",
           441 => x"08",
           442 => x"90",
           443 => x"51",
           444 => x"a4",
           445 => x"82",
           446 => x"83",
           447 => x"72",
           448 => x"08",
           449 => x"98",
           450 => x"81",
           451 => x"34",
           452 => x"e0",
           453 => x"0c",
           454 => x"08",
           455 => x"e0",
           456 => x"2b",
           457 => x"51",
           458 => x"08",
           459 => x"53",
           460 => x"23",
           461 => x"70",
           462 => x"a4",
           463 => x"82",
           464 => x"81",
           465 => x"a4",
           466 => x"82",
           467 => x"80",
           468 => x"a4",
           469 => x"82",
           470 => x"88",
           471 => x"08",
           472 => x"a4",
           473 => x"82",
           474 => x"84",
           475 => x"08",
           476 => x"0b",
           477 => x"82",
           478 => x"11",
           479 => x"ec",
           480 => x"a4",
           481 => x"82",
           482 => x"e0",
           483 => x"82",
           484 => x"08",
           485 => x"fc",
           486 => x"05",
           487 => x"e0",
           488 => x"39",
           489 => x"82",
           490 => x"05",
           491 => x"70",
           492 => x"0c",
           493 => x"70",
           494 => x"51",
           495 => x"e0",
           496 => x"2b",
           497 => x"a4",
           498 => x"83",
           499 => x"82",
           500 => x"39",
           501 => x"51",
           502 => x"53",
           503 => x"23",
           504 => x"53",
           505 => x"73",
           506 => x"a4",
           507 => x"82",
           508 => x"e0",
           509 => x"82",
           510 => x"08",
           511 => x"82",
           512 => x"83",
           513 => x"53",
           514 => x"a4",
           515 => x"53",
           516 => x"08",
           517 => x"3f",
           518 => x"e0",
           519 => x"82",
           520 => x"9b",
           521 => x"72",
           522 => x"82",
           523 => x"82",
           524 => x"71",
           525 => x"08",
           526 => x"e0",
           527 => x"2a",
           528 => x"80",
           529 => x"90",
           530 => x"05",
           531 => x"90",
           532 => x"08",
           533 => x"e0",
           534 => x"a4",
           535 => x"e0",
           536 => x"82",
           537 => x"82",
           538 => x"e0",
           539 => x"a4",
           540 => x"38",
           541 => x"70",
           542 => x"a4",
           543 => x"08",
           544 => x"08",
           545 => x"e4",
           546 => x"53",
           547 => x"23",
           548 => x"a4",
           549 => x"e0",
           550 => x"c0",
           551 => x"08",
           552 => x"e0",
           553 => x"82",
           554 => x"e0",
           555 => x"2a",
           556 => x"80",
           557 => x"90",
           558 => x"05",
           559 => x"90",
           560 => x"08",
           561 => x"e0",
           562 => x"a4",
           563 => x"e0",
           564 => x"82",
           565 => x"82",
           566 => x"e0",
           567 => x"a4",
           568 => x"51",
           569 => x"05",
           570 => x"a4",
           571 => x"08",
           572 => x"f4",
           573 => x"05",
           574 => x"55",
           575 => x"53",
           576 => x"f0",
           577 => x"05",
           578 => x"08",
           579 => x"a4",
           580 => x"08",
           581 => x"08",
           582 => x"51",
           583 => x"d0",
           584 => x"08",
           585 => x"11",
           586 => x"d0",
           587 => x"05",
           588 => x"05",
           589 => x"f0",
           590 => x"08",
           591 => x"f4",
           592 => x"08",
           593 => x"3f",
           594 => x"a4",
           595 => x"a4",
           596 => x"38",
           597 => x"f0",
           598 => x"72",
           599 => x"72",
           600 => x"82",
           601 => x"b2",
           602 => x"38",
           603 => x"ff",
           604 => x"08",
           605 => x"e4",
           606 => x"06",
           607 => x"e7",
           608 => x"22",
           609 => x"cc",
           610 => x"05",
           611 => x"cc",
           612 => x"05",
           613 => x"81",
           614 => x"cc",
           615 => x"e0",
           616 => x"82",
           617 => x"05",
           618 => x"05",
           619 => x"22",
           620 => x"82",
           621 => x"83",
           622 => x"72",
           623 => x"a4",
           624 => x"70",
           625 => x"05",
           626 => x"24",
           627 => x"05",
           628 => x"82",
           629 => x"39",
           630 => x"53",
           631 => x"73",
           632 => x"a4",
           633 => x"08",
           634 => x"81",
           635 => x"b1",
           636 => x"33",
           637 => x"90",
           638 => x"51",
           639 => x"ec",
           640 => x"72",
           641 => x"af",
           642 => x"33",
           643 => x"90",
           644 => x"51",
           645 => x"ec",
           646 => x"72",
           647 => x"82",
           648 => x"83",
           649 => x"82",
           650 => x"11",
           651 => x"ec",
           652 => x"2c",
           653 => x"82",
           654 => x"a0",
           655 => x"e0",
           656 => x"2a",
           657 => x"80",
           658 => x"88",
           659 => x"3f",
           660 => x"e4",
           661 => x"06",
           662 => x"38",
           663 => x"52",
           664 => x"82",
           665 => x"85",
           666 => x"72",
           667 => x"08",
           668 => x"81",
           669 => x"22",
           670 => x"51",
           671 => x"e0",
           672 => x"51",
           673 => x"f4",
           674 => x"81",
           675 => x"88",
           676 => x"f8",
           677 => x"e0",
           678 => x"2a",
           679 => x"80",
           680 => x"ec",
           681 => x"82",
           682 => x"90",
           683 => x"73",
           684 => x"88",
           685 => x"3f",
           686 => x"05",
           687 => x"51",
           688 => x"82",
           689 => x"11",
           690 => x"e8",
           691 => x"2c",
           692 => x"82",
           693 => x"b0",
           694 => x"e0",
           695 => x"2a",
           696 => x"b0",
           697 => x"22",
           698 => x"a4",
           699 => x"70",
           700 => x"90",
           701 => x"08",
           702 => x"39",
           703 => x"53",
           704 => x"97",
           705 => x"08",
           706 => x"33",
           707 => x"82",
           708 => x"72",
           709 => x"cb",
           710 => x"22",
           711 => x"a4",
           712 => x"ff",
           713 => x"81",
           714 => x"05",
           715 => x"05",
           716 => x"08",
           717 => x"a4",
           718 => x"3f",
           719 => x"f8",
           720 => x"09",
           721 => x"a4",
           722 => x"53",
           723 => x"23",
           724 => x"83",
           725 => x"e0",
           726 => x"e0",
           727 => x"52",
           728 => x"08",
           729 => x"a4",
           730 => x"82",
           731 => x"e0",
           732 => x"08",
           733 => x"08",
           734 => x"a4",
           735 => x"08",
           736 => x"85",
           737 => x"08",
           738 => x"81",
           739 => x"80",
           740 => x"05",
           741 => x"e0",
           742 => x"2b",
           743 => x"25",
           744 => x"05",
           745 => x"d2",
           746 => x"08",
           747 => x"33",
           748 => x"e0",
           749 => x"39",
           750 => x"53",
           751 => x"38",
           752 => x"05",
           753 => x"ec",
           754 => x"08",
           755 => x"a4",
           756 => x"82",
           757 => x"82",
           758 => x"84",
           759 => x"a4",
           760 => x"70",
           761 => x"51",
           762 => x"08",
           763 => x"82",
           764 => x"08",
           765 => x"0d",
           766 => x"a4",
           767 => x"a4",
           768 => x"3f",
           769 => x"98",
           770 => x"a4",
           771 => x"82",
           772 => x"0b",
           773 => x"82",
           774 => x"81",
           775 => x"51",
           776 => x"8d",
           777 => x"f4",
           778 => x"a4",
           779 => x"82",
           780 => x"05",
           781 => x"53",
           782 => x"34",
           783 => x"2e",
           784 => x"fb",
           785 => x"fc",
           786 => x"53",
           787 => x"72",
           788 => x"82",
           789 => x"a5",
           790 => x"fc",
           791 => x"08",
           792 => x"53",
           793 => x"82",
           794 => x"e0",
           795 => x"e0",
           796 => x"e0",
           797 => x"98",
           798 => x"0c",
           799 => x"e0",
           800 => x"82",
           801 => x"e0",
           802 => x"33",
           803 => x"81",
           804 => x"80",
           805 => x"a4",
           806 => x"82",
           807 => x"72",
           808 => x"08",
           809 => x"05",
           810 => x"fc",
           811 => x"72",
           812 => x"08",
           813 => x"8c",
           814 => x"fc",
           815 => x"53",
           816 => x"72",
           817 => x"82",
           818 => x"9f",
           819 => x"08",
           820 => x"0c",
           821 => x"08",
           822 => x"82",
           823 => x"08",
           824 => x"0d",
           825 => x"a4",
           826 => x"82",
           827 => x"0c",
           828 => x"0c",
           829 => x"e0",
           830 => x"a4",
           831 => x"70",
           832 => x"06",
           833 => x"2e",
           834 => x"08",
           835 => x"e0",
           836 => x"33",
           837 => x"51",
           838 => x"38",
           839 => x"82",
           840 => x"54",
           841 => x"9f",
           842 => x"08",
           843 => x"88",
           844 => x"75",
           845 => x"82",
           846 => x"11",
           847 => x"e0",
           848 => x"e0",
           849 => x"80",
           850 => x"05",
           851 => x"08",
           852 => x"08",
           853 => x"08",
           854 => x"98",
           855 => x"a4",
           856 => x"81",
           857 => x"08",
           858 => x"08",
           859 => x"ff",
           860 => x"0c",
           861 => x"82",
           862 => x"e0",
           863 => x"02",
           864 => x"82",
           865 => x"11",
           866 => x"51",
           867 => x"38",
           868 => x"05",
           869 => x"08",
           870 => x"86",
           871 => x"52",
           872 => x"e0",
           873 => x"a4",
           874 => x"12",
           875 => x"71",
           876 => x"88",
           877 => x"8c",
           878 => x"05",
           879 => x"a4",
           880 => x"82",
           881 => x"05",
           882 => x"70",
           883 => x"80",
           884 => x"08",
           885 => x"82",
           886 => x"52",
           887 => x"a9",
           888 => x"08",
           889 => x"53",
           890 => x"51",
           891 => x"82",
           892 => x"d7",
           893 => x"08",
           894 => x"81",
           895 => x"05",
           896 => x"08",
           897 => x"2d",
           898 => x"a4",
           899 => x"a4",
           900 => x"f2",
           901 => x"08",
           902 => x"82",
           903 => x"11",
           904 => x"0c",
           905 => x"08",
           906 => x"82",
           907 => x"07",
           908 => x"05",
           909 => x"f0",
           910 => x"e0",
           911 => x"a4",
           912 => x"a4",
           913 => x"ff",
           914 => x"0c",
           915 => x"05",
           916 => x"12",
           917 => x"08",
           918 => x"a4",
           919 => x"82",
           920 => x"e0",
           921 => x"a4",
           922 => x"82",
           923 => x"e0",
           924 => x"a4",
           925 => x"08",
           926 => x"f8",
           927 => x"05",
           928 => x"e0",
           929 => x"a4",
           930 => x"38",
           931 => x"82",
           932 => x"51",
           933 => x"71",
           934 => x"08",
           935 => x"90",
           936 => x"fc",
           937 => x"05",
           938 => x"08",
           939 => x"0c",
           940 => x"81",
           941 => x"0c",
           942 => x"ff",
           943 => x"0c",
           944 => x"80",
           945 => x"08",
           946 => x"a4",
           947 => x"08",
           948 => x"a4",
           949 => x"08",
           950 => x"f8",
           951 => x"34",
           952 => x"90",
           953 => x"08",
           954 => x"90",
           955 => x"08",
           956 => x"90",
           957 => x"e0",
           958 => x"33",
           959 => x"81",
           960 => x"0c",
           961 => x"52",
           962 => x"08",
           963 => x"a4",
           964 => x"82",
           965 => x"82",
           966 => x"82",
           967 => x"08",
           968 => x"0d",
           969 => x"82",
           970 => x"e0",
           971 => x"33",
           972 => x"81",
           973 => x"0c",
           974 => x"80",
           975 => x"a4",
           976 => x"e0",
           977 => x"a4",
           978 => x"08",
           979 => x"98",
           980 => x"a4",
           981 => x"82",
           982 => x"e0",
           983 => x"a4",
           984 => x"08",
           985 => x"e0",
           986 => x"82",
           987 => x"e0",
           988 => x"70",
           989 => x"05",
           990 => x"fc",
           991 => x"70",
           992 => x"82",
           993 => x"82",
           994 => x"82",
           995 => x"08",
           996 => x"0d",
           997 => x"82",
           998 => x"e0",
           999 => x"a4",
          1000 => x"08",
          1001 => x"38",
          1002 => x"81",
          1003 => x"0c",
          1004 => x"ff",
          1005 => x"0c",
          1006 => x"80",
          1007 => x"f8",
          1008 => x"a4",
          1009 => x"e0",
          1010 => x"a4",
          1011 => x"71",
          1012 => x"08",
          1013 => x"05",
          1014 => x"08",
          1015 => x"0c",
          1016 => x"0c",
          1017 => x"e0",
          1018 => x"a4",
          1019 => x"f4",
          1020 => x"08",
          1021 => x"8c",
          1022 => x"08",
          1023 => x"88",
          1024 => x"06",
          1025 => x"84",
          1026 => x"08",
          1027 => x"e0",
          1028 => x"82",
          1029 => x"81",
          1030 => x"80",
          1031 => x"0c",
          1032 => x"90",
          1033 => x"08",
          1034 => x"90",
          1035 => x"81",
          1036 => x"08",
          1037 => x"a4",
          1038 => x"53",
          1039 => x"a4",
          1040 => x"82",
          1041 => x"05",
          1042 => x"82",
          1043 => x"33",
          1044 => x"82",
          1045 => x"39",
          1046 => x"70",
          1047 => x"08",
          1048 => x"e0",
          1049 => x"52",
          1050 => x"e0",
          1051 => x"a4",
          1052 => x"0c",
          1053 => x"04",
          1054 => x"a4",
          1055 => x"08",
          1056 => x"08",
          1057 => x"82",
          1058 => x"08",
          1059 => x"f8",
          1060 => x"54",
          1061 => x"08",
          1062 => x"0c",
          1063 => x"08",
          1064 => x"08",
          1065 => x"a4",
          1066 => x"08",
          1067 => x"34",
          1068 => x"53",
          1069 => x"52",
          1070 => x"51",
          1071 => x"70",
          1072 => x"54",
          1073 => x"82",
          1074 => x"e0",
          1075 => x"02",
          1076 => x"82",
          1077 => x"e0",
          1078 => x"a4",
          1079 => x"0b",
          1080 => x"80",
          1081 => x"05",
          1082 => x"08",
          1083 => x"a4",
          1084 => x"06",
          1085 => x"82",
          1086 => x"05",
          1087 => x"82",
          1088 => x"2e",
          1089 => x"a4",
          1090 => x"e0",
          1091 => x"a4",
          1092 => x"08",
          1093 => x"a4",
          1094 => x"a4",
          1095 => x"0c",
          1096 => x"04",
          1097 => x"a4",
          1098 => x"08",
          1099 => x"fc",
          1100 => x"05",
          1101 => x"e0",
          1102 => x"82",
          1103 => x"e0",
          1104 => x"82",
          1105 => x"e0",
          1106 => x"a9",
          1107 => x"08",
          1108 => x"05",
          1109 => x"e0",
          1110 => x"82",
          1111 => x"be",
          1112 => x"08",
          1113 => x"3d",
          1114 => x"e0",
          1115 => x"fe",
          1116 => x"05",
          1117 => x"05",
          1118 => x"08",
          1119 => x"3d",
          1120 => x"e0",
          1121 => x"f6",
          1122 => x"08",
          1123 => x"8c",
          1124 => x"e0",
          1125 => x"fc",
          1126 => x"e0",
          1127 => x"39",
          1128 => x"82",
          1129 => x"e0",
          1130 => x"a3",
          1131 => x"08",
          1132 => x"08",
          1133 => x"71",
          1134 => x"0c",
          1135 => x"e4",
          1136 => x"05",
          1137 => x"05",
          1138 => x"08",
          1139 => x"82",
          1140 => x"05",
          1141 => x"05",
          1142 => x"e0",
          1143 => x"39",
          1144 => x"ff",
          1145 => x"f8",
          1146 => x"38",
          1147 => x"70",
          1148 => x"52",
          1149 => x"f8",
          1150 => x"08",
          1151 => x"88",
          1152 => x"05",
          1153 => x"05",
          1154 => x"08",
          1155 => x"31",
          1156 => x"71",
          1157 => x"0c",
          1158 => x"f0",
          1159 => x"05",
          1160 => x"e0",
          1161 => x"e0",
          1162 => x"82",
          1163 => x"2a",
          1164 => x"f4",
          1165 => x"05",
          1166 => x"f0",
          1167 => x"88",
          1168 => x"05",
          1169 => x"08",
          1170 => x"fc",
          1171 => x"82",
          1172 => x"e0",
          1173 => x"82",
          1174 => x"e0",
          1175 => x"a4",
          1176 => x"a4",
          1177 => x"e0",
          1178 => x"a4",
          1179 => x"e0",
          1180 => x"55",
          1181 => x"39",
          1182 => x"10",
          1183 => x"08",
          1184 => x"0c",
          1185 => x"70",
          1186 => x"51",
          1187 => x"08",
          1188 => x"82",
          1189 => x"08",
          1190 => x"0d",
          1191 => x"82",
          1192 => x"e0",
          1193 => x"80",
          1194 => x"82",
          1195 => x"39",
          1196 => x"05",
          1197 => x"08",
          1198 => x"90",
          1199 => x"08",
          1200 => x"08",
          1201 => x"05",
          1202 => x"08",
          1203 => x"82",
          1204 => x"fe",
          1205 => x"88",
          1206 => x"0c",
          1207 => x"08",
          1208 => x"ec",
          1209 => x"05",
          1210 => x"f8",
          1211 => x"fc",
          1212 => x"08",
          1213 => x"f4",
          1214 => x"05",
          1215 => x"05",
          1216 => x"08",
          1217 => x"38",
          1218 => x"05",
          1219 => x"a4",
          1220 => x"08",
          1221 => x"f8",
          1222 => x"08",
          1223 => x"08",
          1224 => x"a4",
          1225 => x"08",
          1226 => x"f8",
          1227 => x"f4",
          1228 => x"05",
          1229 => x"38",
          1230 => x"05",
          1231 => x"a4",
          1232 => x"08",
          1233 => x"f8",
          1234 => x"08",
          1235 => x"08",
          1236 => x"a4",
          1237 => x"08",
          1238 => x"f8",
          1239 => x"f4",
          1240 => x"08",
          1241 => x"08",
          1242 => x"32",
          1243 => x"06",
          1244 => x"11",
          1245 => x"51",
          1246 => x"8a",
          1247 => x"82",
          1248 => x"0c",
          1249 => x"8c",
          1250 => x"88",
          1251 => x"e0",
          1252 => x"8c",
          1253 => x"88",
          1254 => x"98",
          1255 => x"82",
          1256 => x"08",
          1257 => x"0d",
          1258 => x"52",
          1259 => x"51",
          1260 => x"82",
          1261 => x"82",
          1262 => x"08",
          1263 => x"0d",
          1264 => x"05",
          1265 => x"08",
          1266 => x"08",
          1267 => x"82",
          1268 => x"08",
          1269 => x"e0",
          1270 => x"a4",
          1271 => x"08",
          1272 => x"82",
          1273 => x"fa",
          1274 => x"e0",
          1275 => x"82",
          1276 => x"97",
          1277 => x"08",
          1278 => x"31",
          1279 => x"82",
          1280 => x"e0",
          1281 => x"a4",
          1282 => x"71",
          1283 => x"27",
          1284 => x"05",
          1285 => x"05",
          1286 => x"a4",
          1287 => x"71",
          1288 => x"2e",
          1289 => x"82",
          1290 => x"96",
          1291 => x"08",
          1292 => x"05",
          1293 => x"08",
          1294 => x"2a",
          1295 => x"82",
          1296 => x"e0",
          1297 => x"e0",
          1298 => x"82",
          1299 => x"80",
          1300 => x"0c",
          1301 => x"80",
          1302 => x"08",
          1303 => x"08",
          1304 => x"a4",
          1305 => x"73",
          1306 => x"0c",
          1307 => x"10",
          1308 => x"08",
          1309 => x"0c",
          1310 => x"82",
          1311 => x"ff",
          1312 => x"08",
          1313 => x"a4",
          1314 => x"08",
          1315 => x"a4",
          1316 => x"08",
          1317 => x"ec",
          1318 => x"f4",
          1319 => x"08",
          1320 => x"f8",
          1321 => x"08",
          1322 => x"51",
          1323 => x"e0",
          1324 => x"e0",
          1325 => x"e0",
          1326 => x"98",
          1327 => x"0c",
          1328 => x"e0",
          1329 => x"82",
          1330 => x"e0",
          1331 => x"a4",
          1332 => x"a4",
          1333 => x"08",
          1334 => x"fc",
          1335 => x"f4",
          1336 => x"05",
          1337 => x"08",
          1338 => x"05",
          1339 => x"05",
          1340 => x"08",
          1341 => x"32",
          1342 => x"08",
          1343 => x"0c",
          1344 => x"82",
          1345 => x"82",
          1346 => x"e0",
          1347 => x"e0",
          1348 => x"53",
          1349 => x"70",
          1350 => x"32",
          1351 => x"08",
          1352 => x"51",
          1353 => x"0c",
          1354 => x"e0",
          1355 => x"82",
          1356 => x"e0",
          1357 => x"73",
          1358 => x"08",
          1359 => x"72",
          1360 => x"72",
          1361 => x"09",
          1362 => x"08",
          1363 => x"71",
          1364 => x"08",
          1365 => x"09",
          1366 => x"e0",
          1367 => x"a4",
          1368 => x"05",
          1369 => x"33",
          1370 => x"82",
          1371 => x"72",
          1372 => x"38",
          1373 => x"70",
          1374 => x"51",
          1375 => x"f8",
          1376 => x"05",
          1377 => x"0c",
          1378 => x"80",
          1379 => x"08",
          1380 => x"38",
          1381 => x"a4",
          1382 => x"08",
          1383 => x"71",
          1384 => x"82",
          1385 => x"a4",
          1386 => x"f4",
          1387 => x"05",
          1388 => x"70",
          1389 => x"a4",
          1390 => x"82",
          1391 => x"72",
          1392 => x"e0",
          1393 => x"39",
          1394 => x"53",
          1395 => x"a4",
          1396 => x"26",
          1397 => x"e0",
          1398 => x"39",
          1399 => x"05",
          1400 => x"f8",
          1401 => x"38",
          1402 => x"53",
          1403 => x"80",
          1404 => x"0c",
          1405 => x"a4",
          1406 => x"e0",
          1407 => x"a4",
          1408 => x"27",
          1409 => x"f8",
          1410 => x"94",
          1411 => x"33",
          1412 => x"a4",
          1413 => x"08",
          1414 => x"72",
          1415 => x"82",
          1416 => x"90",
          1417 => x"08",
          1418 => x"72",
          1419 => x"82",
          1420 => x"72",
          1421 => x"e0",
          1422 => x"39",
          1423 => x"82",
          1424 => x"54",
          1425 => x"82",
          1426 => x"f7",
          1427 => x"33",
          1428 => x"08",
          1429 => x"33",
          1430 => x"05",
          1431 => x"08",
          1432 => x"08",
          1433 => x"82",
          1434 => x"a5",
          1435 => x"33",
          1436 => x"e0",
          1437 => x"e0",
          1438 => x"a4",
          1439 => x"08",
          1440 => x"0b",
          1441 => x"82",
          1442 => x"e0",
          1443 => x"a4",
          1444 => x"82",
          1445 => x"0b",
          1446 => x"82",
          1447 => x"80",
          1448 => x"05",
          1449 => x"53",
          1450 => x"34",
          1451 => x"2e",
          1452 => x"a4",
          1453 => x"05",
          1454 => x"a4",
          1455 => x"2e",
          1456 => x"82",
          1457 => x"e0",
          1458 => x"81",
          1459 => x"72",
          1460 => x"34",
          1461 => x"53",
          1462 => x"dc",
          1463 => x"08",
          1464 => x"08",
          1465 => x"08",
          1466 => x"f8",
          1467 => x"05",
          1468 => x"08",
          1469 => x"a4",
          1470 => x"84",
          1471 => x"e0",
          1472 => x"a4",
          1473 => x"05",
          1474 => x"33",
          1475 => x"81",
          1476 => x"08",
          1477 => x"88",
          1478 => x"0c",
          1479 => x"e0",
          1480 => x"39",
          1481 => x"53",
          1482 => x"82",
          1483 => x"80",
          1484 => x"33",
          1485 => x"e0",
          1486 => x"b9",
          1487 => x"82",
          1488 => x"d8",
          1489 => x"f4",
          1490 => x"08",
          1491 => x"90",
          1492 => x"33",
          1493 => x"39",
          1494 => x"05",
          1495 => x"e0",
          1496 => x"82",
          1497 => x"e0",
          1498 => x"73",
          1499 => x"08",
          1500 => x"27",
          1501 => x"05",
          1502 => x"e0",
          1503 => x"a4",
          1504 => x"53",
          1505 => x"34",
          1506 => x"53",
          1507 => x"a4",
          1508 => x"53",
          1509 => x"34",
          1510 => x"53",
          1511 => x"82",
          1512 => x"98",
          1513 => x"33",
          1514 => x"54",
          1515 => x"0b",
          1516 => x"80",
          1517 => x"05",
          1518 => x"05",
          1519 => x"05",
          1520 => x"fc",
          1521 => x"05",
          1522 => x"70",
          1523 => x"33",
          1524 => x"fe",
          1525 => x"05",
          1526 => x"82",
          1527 => x"82",
          1528 => x"e0",
          1529 => x"a4",
          1530 => x"81",
          1531 => x"0c",
          1532 => x"82",
          1533 => x"e0",
          1534 => x"70",
          1535 => x"2e",
          1536 => x"79",
          1537 => x"39",
          1538 => x"81",
          1539 => x"39",
          1540 => x"a0",
          1541 => x"3f",
          1542 => x"08",
          1543 => x"df",
          1544 => x"38",
          1545 => x"ff",
          1546 => x"06",
          1547 => x"ff",
          1548 => x"3d",
          1549 => x"98",
          1550 => x"71",
          1551 => x"29",
          1552 => x"04",
          1553 => x"82",
          1554 => x"be",
          1555 => x"90",
          1556 => x"51",
          1557 => x"80",
          1558 => x"d6",
          1559 => x"39",
          1560 => x"82",
          1561 => x"bf",
          1562 => x"51",
          1563 => x"39",
          1564 => x"c0",
          1565 => x"51",
          1566 => x"39",
          1567 => x"c0",
          1568 => x"51",
          1569 => x"8a",
          1570 => x"0d",
          1571 => x"26",
          1572 => x"29",
          1573 => x"51",
          1574 => x"52",
          1575 => x"98",
          1576 => x"c1",
          1577 => x"3d",
          1578 => x"84",
          1579 => x"80",
          1580 => x"25",
          1581 => x"87",
          1582 => x"76",
          1583 => x"93",
          1584 => x"76",
          1585 => x"93",
          1586 => x"82",
          1587 => x"98",
          1588 => x"e0",
          1589 => x"54",
          1590 => x"81",
          1591 => x"57",
          1592 => x"55",
          1593 => x"75",
          1594 => x"d8",
          1595 => x"30",
          1596 => x"70",
          1597 => x"56",
          1598 => x"bc",
          1599 => x"78",
          1600 => x"82",
          1601 => x"f8",
          1602 => x"05",
          1603 => x"7b",
          1604 => x"e0",
          1605 => x"88",
          1606 => x"39",
          1607 => x"54",
          1608 => x"51",
          1609 => x"83",
          1610 => x"0c",
          1611 => x"7f",
          1612 => x"05",
          1613 => x"5d",
          1614 => x"fb",
          1615 => x"ff",
          1616 => x"92",
          1617 => x"8a",
          1618 => x"39",
          1619 => x"51",
          1620 => x"51",
          1621 => x"78",
          1622 => x"89",
          1623 => x"c6",
          1624 => x"8e",
          1625 => x"51",
          1626 => x"c1",
          1627 => x"15",
          1628 => x"72",
          1629 => x"82",
          1630 => x"89",
          1631 => x"8f",
          1632 => x"19",
          1633 => x"33",
          1634 => x"f7",
          1635 => x"ff",
          1636 => x"fb",
          1637 => x"3f",
          1638 => x"ff",
          1639 => x"27",
          1640 => x"55",
          1641 => x"38",
          1642 => x"83",
          1643 => x"81",
          1644 => x"90",
          1645 => x"82",
          1646 => x"39",
          1647 => x"cc",
          1648 => x"39",
          1649 => x"77",
          1650 => x"98",
          1651 => x"2b",
          1652 => x"2e",
          1653 => x"98",
          1654 => x"2b",
          1655 => x"30",
          1656 => x"07",
          1657 => x"59",
          1658 => x"38",
          1659 => x"1e",
          1660 => x"ff",
          1661 => x"3d",
          1662 => x"05",
          1663 => x"82",
          1664 => x"ff",
          1665 => x"51",
          1666 => x"82",
          1667 => x"52",
          1668 => x"3f",
          1669 => x"3f",
          1670 => x"87",
          1671 => x"3f",
          1672 => x"b4",
          1673 => x"b3",
          1674 => x"51",
          1675 => x"51",
          1676 => x"9a",
          1677 => x"72",
          1678 => x"71",
          1679 => x"83",
          1680 => x"3f",
          1681 => x"2a",
          1682 => x"2e",
          1683 => x"82",
          1684 => x"51",
          1685 => x"81",
          1686 => x"38",
          1687 => x"80",
          1688 => x"bb",
          1689 => x"51",
          1690 => x"51",
          1691 => x"99",
          1692 => x"72",
          1693 => x"71",
          1694 => x"8b",
          1695 => x"3f",
          1696 => x"2a",
          1697 => x"2e",
          1698 => x"82",
          1699 => x"51",
          1700 => x"81",
          1701 => x"38",
          1702 => x"d0",
          1703 => x"c3",
          1704 => x"04",
          1705 => x"a3",
          1706 => x"52",
          1707 => x"82",
          1708 => x"81",
          1709 => x"a8",
          1710 => x"98",
          1711 => x"07",
          1712 => x"54",
          1713 => x"0b",
          1714 => x"81",
          1715 => x"f7",
          1716 => x"c7",
          1717 => x"2e",
          1718 => x"c4",
          1719 => x"51",
          1720 => x"0b",
          1721 => x"db",
          1722 => x"81",
          1723 => x"74",
          1724 => x"0b",
          1725 => x"04",
          1726 => x"ff",
          1727 => x"52",
          1728 => x"e0",
          1729 => x"7e",
          1730 => x"3d",
          1731 => x"78",
          1732 => x"52",
          1733 => x"3f",
          1734 => x"38",
          1735 => x"81",
          1736 => x"ff",
          1737 => x"5a",
          1738 => x"3f",
          1739 => x"93",
          1740 => x"70",
          1741 => x"2e",
          1742 => x"b2",
          1743 => x"78",
          1744 => x"ff",
          1745 => x"38",
          1746 => x"83",
          1747 => x"ce",
          1748 => x"8a",
          1749 => x"df",
          1750 => x"78",
          1751 => x"80",
          1752 => x"39",
          1753 => x"78",
          1754 => x"82",
          1755 => x"78",
          1756 => x"86",
          1757 => x"ff",
          1758 => x"e0",
          1759 => x"b5",
          1760 => x"05",
          1761 => x"08",
          1762 => x"fe",
          1763 => x"ec",
          1764 => x"38",
          1765 => x"e8",
          1766 => x"5c",
          1767 => x"62",
          1768 => x"0c",
          1769 => x"39",
          1770 => x"84",
          1771 => x"98",
          1772 => x"3d",
          1773 => x"51",
          1774 => x"80",
          1775 => x"f8",
          1776 => x"9a",
          1777 => x"fd",
          1778 => x"a4",
          1779 => x"81",
          1780 => x"05",
          1781 => x"43",
          1782 => x"53",
          1783 => x"82",
          1784 => x"38",
          1785 => x"84",
          1786 => x"98",
          1787 => x"3d",
          1788 => x"51",
          1789 => x"80",
          1790 => x"51",
          1791 => x"64",
          1792 => x"33",
          1793 => x"38",
          1794 => x"79",
          1795 => x"ef",
          1796 => x"5a",
          1797 => x"fc",
          1798 => x"53",
          1799 => x"82",
          1800 => x"de",
          1801 => x"38",
          1802 => x"39",
          1803 => x"2e",
          1804 => x"bc",
          1805 => x"80",
          1806 => x"45",
          1807 => x"78",
          1808 => x"08",
          1809 => x"59",
          1810 => x"d4",
          1811 => x"08",
          1812 => x"fc",
          1813 => x"f2",
          1814 => x"38",
          1815 => x"2e",
          1816 => x"80",
          1817 => x"78",
          1818 => x"08",
          1819 => x"59",
          1820 => x"c8",
          1821 => x"33",
          1822 => x"de",
          1823 => x"fa",
          1824 => x"82",
          1825 => x"de",
          1826 => x"fe",
          1827 => x"e8",
          1828 => x"2e",
          1829 => x"88",
          1830 => x"32",
          1831 => x"70",
          1832 => x"80",
          1833 => x"38",
          1834 => x"bd",
          1835 => x"53",
          1836 => x"82",
          1837 => x"3d",
          1838 => x"51",
          1839 => x"80",
          1840 => x"fc",
          1841 => x"92",
          1842 => x"a4",
          1843 => x"33",
          1844 => x"3d",
          1845 => x"51",
          1846 => x"e1",
          1847 => x"54",
          1848 => x"c7",
          1849 => x"f8",
          1850 => x"79",
          1851 => x"f8",
          1852 => x"b5",
          1853 => x"05",
          1854 => x"08",
          1855 => x"80",
          1856 => x"05",
          1857 => x"51",
          1858 => x"b5",
          1859 => x"05",
          1860 => x"08",
          1861 => x"fe",
          1862 => x"e0",
          1863 => x"2e",
          1864 => x"05",
          1865 => x"78",
          1866 => x"ff",
          1867 => x"e0",
          1868 => x"61",
          1869 => x"51",
          1870 => x"08",
          1871 => x"9f",
          1872 => x"78",
          1873 => x"26",
          1874 => x"39",
          1875 => x"84",
          1876 => x"98",
          1877 => x"02",
          1878 => x"05",
          1879 => x"82",
          1880 => x"ff",
          1881 => x"53",
          1882 => x"82",
          1883 => x"38",
          1884 => x"84",
          1885 => x"98",
          1886 => x"71",
          1887 => x"3d",
          1888 => x"51",
          1889 => x"e5",
          1890 => x"54",
          1891 => x"ef",
          1892 => x"f8",
          1893 => x"79",
          1894 => x"f6",
          1895 => x"b5",
          1896 => x"05",
          1897 => x"08",
          1898 => x"0c",
          1899 => x"39",
          1900 => x"3f",
          1901 => x"11",
          1902 => x"3f",
          1903 => x"c3",
          1904 => x"ff",
          1905 => x"b5",
          1906 => x"05",
          1907 => x"08",
          1908 => x"82",
          1909 => x"64",
          1910 => x"80",
          1911 => x"08",
          1912 => x"c7",
          1913 => x"51",
          1914 => x"3f",
          1915 => x"ff",
          1916 => x"39",
          1917 => x"3d",
          1918 => x"38",
          1919 => x"3f",
          1920 => x"98",
          1921 => x"e0",
          1922 => x"05",
          1923 => x"08",
          1924 => x"2e",
          1925 => x"51",
          1926 => x"8f",
          1927 => x"82",
          1928 => x"38",
          1929 => x"39",
          1930 => x"39",
          1931 => x"c6",
          1932 => x"52",
          1933 => x"9e",
          1934 => x"3d",
          1935 => x"ab",
          1936 => x"80",
          1937 => x"ff",
          1938 => x"93",
          1939 => x"9c",
          1940 => x"ff",
          1941 => x"82",
          1942 => x"80",
          1943 => x"0a",
          1944 => x"ea",
          1945 => x"e0",
          1946 => x"07",
          1947 => x"5a",
          1948 => x"78",
          1949 => x"38",
          1950 => x"59",
          1951 => x"7e",
          1952 => x"7e",
          1953 => x"82",
          1954 => x"7c",
          1955 => x"82",
          1956 => x"f2",
          1957 => x"82",
          1958 => x"70",
          1959 => x"72",
          1960 => x"08",
          1961 => x"84",
          1962 => x"72",
          1963 => x"87",
          1964 => x"87",
          1965 => x"3f",
          1966 => x"08",
          1967 => x"51",
          1968 => x"08",
          1969 => x"87",
          1970 => x"0b",
          1971 => x"98",
          1972 => x"84",
          1973 => x"fb",
          1974 => x"0c",
          1975 => x"54",
          1976 => x"c7",
          1977 => x"c7",
          1978 => x"e8",
          1979 => x"ec",
          1980 => x"fc",
          1981 => x"80",
          1982 => x"8a",
          1983 => x"09",
          1984 => x"f1",
          1985 => x"09",
          1986 => x"81",
          1987 => x"81",
          1988 => x"52",
          1989 => x"2e",
          1990 => x"9d",
          1991 => x"12",
          1992 => x"a0",
          1993 => x"2e",
          1994 => x"33",
          1995 => x"06",
          1996 => x"70",
          1997 => x"51",
          1998 => x"72",
          1999 => x"0c",
          2000 => x"86",
          2001 => x"53",
          2002 => x"3d",
          2003 => x"3f",
          2004 => x"53",
          2005 => x"98",
          2006 => x"0d",
          2007 => x"53",
          2008 => x"38",
          2009 => x"52",
          2010 => x"13",
          2011 => x"80",
          2012 => x"52",
          2013 => x"13",
          2014 => x"80",
          2015 => x"52",
          2016 => x"8a",
          2017 => x"e7",
          2018 => x"c0",
          2019 => x"98",
          2020 => x"98",
          2021 => x"98",
          2022 => x"98",
          2023 => x"98",
          2024 => x"98",
          2025 => x"0c",
          2026 => x"0b",
          2027 => x"71",
          2028 => x"04",
          2029 => x"98",
          2030 => x"98",
          2031 => x"c0",
          2032 => x"34",
          2033 => x"83",
          2034 => x"5a",
          2035 => x"ac",
          2036 => x"c0",
          2037 => x"34",
          2038 => x"88",
          2039 => x"5a",
          2040 => x"79",
          2041 => x"ff",
          2042 => x"85",
          2043 => x"83",
          2044 => x"7d",
          2045 => x"84",
          2046 => x"0d",
          2047 => x"33",
          2048 => x"81",
          2049 => x"32",
          2050 => x"51",
          2051 => x"84",
          2052 => x"82",
          2053 => x"2c",
          2054 => x"06",
          2055 => x"09",
          2056 => x"83",
          2057 => x"07",
          2058 => x"71",
          2059 => x"04",
          2060 => x"72",
          2061 => x"3f",
          2062 => x"98",
          2063 => x"52",
          2064 => x"e0",
          2065 => x"3d",
          2066 => x"b0",
          2067 => x"55",
          2068 => x"2e",
          2069 => x"70",
          2070 => x"53",
          2071 => x"71",
          2072 => x"70",
          2073 => x"06",
          2074 => x"71",
          2075 => x"70",
          2076 => x"51",
          2077 => x"2e",
          2078 => x"74",
          2079 => x"87",
          2080 => x"8f",
          2081 => x"51",
          2082 => x"83",
          2083 => x"a7",
          2084 => x"81",
          2085 => x"eb",
          2086 => x"ff",
          2087 => x"53",
          2088 => x"94",
          2089 => x"70",
          2090 => x"2e",
          2091 => x"06",
          2092 => x"32",
          2093 => x"2e",
          2094 => x"06",
          2095 => x"81",
          2096 => x"54",
          2097 => x"94",
          2098 => x"82",
          2099 => x"f9",
          2100 => x"70",
          2101 => x"77",
          2102 => x"06",
          2103 => x"81",
          2104 => x"c0",
          2105 => x"38",
          2106 => x"70",
          2107 => x"52",
          2108 => x"2a",
          2109 => x"38",
          2110 => x"51",
          2111 => x"2a",
          2112 => x"be",
          2113 => x"c0",
          2114 => x"38",
          2115 => x"0c",
          2116 => x"06",
          2117 => x"76",
          2118 => x"04",
          2119 => x"70",
          2120 => x"94",
          2121 => x"87",
          2122 => x"82",
          2123 => x"70",
          2124 => x"06",
          2125 => x"80",
          2126 => x"52",
          2127 => x"e0",
          2128 => x"ff",
          2129 => x"ff",
          2130 => x"3d",
          2131 => x"ff",
          2132 => x"52",
          2133 => x"94",
          2134 => x"70",
          2135 => x"70",
          2136 => x"06",
          2137 => x"80",
          2138 => x"52",
          2139 => x"2c",
          2140 => x"0c",
          2141 => x"87",
          2142 => x"8a",
          2143 => x"b4",
          2144 => x"de",
          2145 => x"82",
          2146 => x"08",
          2147 => x"98",
          2148 => x"9e",
          2149 => x"c0",
          2150 => x"87",
          2151 => x"0c",
          2152 => x"d0",
          2153 => x"de",
          2154 => x"82",
          2155 => x"08",
          2156 => x"c0",
          2157 => x"9e",
          2158 => x"c0",
          2159 => x"e8",
          2160 => x"de",
          2161 => x"82",
          2162 => x"08",
          2163 => x"de",
          2164 => x"90",
          2165 => x"52",
          2166 => x"52",
          2167 => x"87",
          2168 => x"0a",
          2169 => x"83",
          2170 => x"34",
          2171 => x"70",
          2172 => x"70",
          2173 => x"82",
          2174 => x"9e",
          2175 => x"51",
          2176 => x"81",
          2177 => x"0b",
          2178 => x"80",
          2179 => x"2e",
          2180 => x"fd",
          2181 => x"08",
          2182 => x"52",
          2183 => x"71",
          2184 => x"c0",
          2185 => x"06",
          2186 => x"38",
          2187 => x"80",
          2188 => x"82",
          2189 => x"80",
          2190 => x"df",
          2191 => x"90",
          2192 => x"52",
          2193 => x"52",
          2194 => x"87",
          2195 => x"80",
          2196 => x"83",
          2197 => x"34",
          2198 => x"70",
          2199 => x"80",
          2200 => x"df",
          2201 => x"70",
          2202 => x"51",
          2203 => x"0b",
          2204 => x"80",
          2205 => x"83",
          2206 => x"34",
          2207 => x"f0",
          2208 => x"70",
          2209 => x"c0",
          2210 => x"52",
          2211 => x"52",
          2212 => x"9e",
          2213 => x"70",
          2214 => x"04",
          2215 => x"ff",
          2216 => x"54",
          2217 => x"b0",
          2218 => x"c4",
          2219 => x"fa",
          2220 => x"82",
          2221 => x"11",
          2222 => x"89",
          2223 => x"73",
          2224 => x"08",
          2225 => x"82",
          2226 => x"82",
          2227 => x"94",
          2228 => x"b8",
          2229 => x"51",
          2230 => x"33",
          2231 => x"de",
          2232 => x"54",
          2233 => x"bf",
          2234 => x"80",
          2235 => x"82",
          2236 => x"c9",
          2237 => x"df",
          2238 => x"38",
          2239 => x"e8",
          2240 => x"87",
          2241 => x"82",
          2242 => x"51",
          2243 => x"33",
          2244 => x"df",
          2245 => x"ff",
          2246 => x"54",
          2247 => x"c8",
          2248 => x"fb",
          2249 => x"82",
          2250 => x"82",
          2251 => x"89",
          2252 => x"b2",
          2253 => x"80",
          2254 => x"ff",
          2255 => x"54",
          2256 => x"fc",
          2257 => x"84",
          2258 => x"dc",
          2259 => x"86",
          2260 => x"82",
          2261 => x"82",
          2262 => x"51",
          2263 => x"51",
          2264 => x"22",
          2265 => x"bf",
          2266 => x"84",
          2267 => x"3f",
          2268 => x"29",
          2269 => x"98",
          2270 => x"86",
          2271 => x"73",
          2272 => x"08",
          2273 => x"ff",
          2274 => x"bd",
          2275 => x"54",
          2276 => x"e4",
          2277 => x"fa",
          2278 => x"82",
          2279 => x"52",
          2280 => x"e0",
          2281 => x"71",
          2282 => x"52",
          2283 => x"3f",
          2284 => x"3d",
          2285 => x"05",
          2286 => x"aa",
          2287 => x"05",
          2288 => x"51",
          2289 => x"39",
          2290 => x"cd",
          2291 => x"51",
          2292 => x"84",
          2293 => x"88",
          2294 => x"96",
          2295 => x"87",
          2296 => x"0d",
          2297 => x"98",
          2298 => x"70",
          2299 => x"51",
          2300 => x"55",
          2301 => x"cd",
          2302 => x"97",
          2303 => x"70",
          2304 => x"81",
          2305 => x"3d",
          2306 => x"84",
          2307 => x"56",
          2308 => x"fb",
          2309 => x"b9",
          2310 => x"51",
          2311 => x"08",
          2312 => x"73",
          2313 => x"72",
          2314 => x"51",
          2315 => x"87",
          2316 => x"02",
          2317 => x"05",
          2318 => x"70",
          2319 => x"08",
          2320 => x"80",
          2321 => x"3f",
          2322 => x"82",
          2323 => x"58",
          2324 => x"98",
          2325 => x"70",
          2326 => x"08",
          2327 => x"38",
          2328 => x"ac",
          2329 => x"05",
          2330 => x"81",
          2331 => x"38",
          2332 => x"80",
          2333 => x"56",
          2334 => x"e0",
          2335 => x"fc",
          2336 => x"51",
          2337 => x"08",
          2338 => x"82",
          2339 => x"3f",
          2340 => x"82",
          2341 => x"52",
          2342 => x"99",
          2343 => x"84",
          2344 => x"38",
          2345 => x"df",
          2346 => x"38",
          2347 => x"df",
          2348 => x"0b",
          2349 => x"04",
          2350 => x"82",
          2351 => x"3f",
          2352 => x"82",
          2353 => x"88",
          2354 => x"3f",
          2355 => x"38",
          2356 => x"e0",
          2357 => x"98",
          2358 => x"08",
          2359 => x"74",
          2360 => x"82",
          2361 => x"3f",
          2362 => x"af",
          2363 => x"0d",
          2364 => x"5a",
          2365 => x"df",
          2366 => x"82",
          2367 => x"0b",
          2368 => x"f8",
          2369 => x"9e",
          2370 => x"2e",
          2371 => x"3f",
          2372 => x"55",
          2373 => x"8e",
          2374 => x"70",
          2375 => x"09",
          2376 => x"51",
          2377 => x"73",
          2378 => x"8c",
          2379 => x"3f",
          2380 => x"38",
          2381 => x"3f",
          2382 => x"38",
          2383 => x"3f",
          2384 => x"3d",
          2385 => x"34",
          2386 => x"a9",
          2387 => x"7e",
          2388 => x"5a",
          2389 => x"a2",
          2390 => x"76",
          2391 => x"70",
          2392 => x"2e",
          2393 => x"26",
          2394 => x"82",
          2395 => x"ff",
          2396 => x"53",
          2397 => x"d9",
          2398 => x"38",
          2399 => x"88",
          2400 => x"39",
          2401 => x"5a",
          2402 => x"51",
          2403 => x"80",
          2404 => x"52",
          2405 => x"98",
          2406 => x"38",
          2407 => x"81",
          2408 => x"ff",
          2409 => x"98",
          2410 => x"0d",
          2411 => x"3d",
          2412 => x"3d",
          2413 => x"e4",
          2414 => x"73",
          2415 => x"83",
          2416 => x"bc",
          2417 => x"73",
          2418 => x"98",
          2419 => x"df",
          2420 => x"2e",
          2421 => x"82",
          2422 => x"3f",
          2423 => x"38",
          2424 => x"3f",
          2425 => x"5b",
          2426 => x"52",
          2427 => x"f8",
          2428 => x"e0",
          2429 => x"80",
          2430 => x"ff",
          2431 => x"55",
          2432 => x"a9",
          2433 => x"70",
          2434 => x"53",
          2435 => x"f8",
          2436 => x"06",
          2437 => x"80",
          2438 => x"ff",
          2439 => x"e0",
          2440 => x"08",
          2441 => x"8f",
          2442 => x"82",
          2443 => x"2c",
          2444 => x"78",
          2445 => x"70",
          2446 => x"d0",
          2447 => x"71",
          2448 => x"cd",
          2449 => x"51",
          2450 => x"5d",
          2451 => x"e9",
          2452 => x"81",
          2453 => x"70",
          2454 => x"80",
          2455 => x"51",
          2456 => x"81",
          2457 => x"38",
          2458 => x"b1",
          2459 => x"80",
          2460 => x"ff",
          2461 => x"97",
          2462 => x"f5",
          2463 => x"ff",
          2464 => x"80",
          2465 => x"81",
          2466 => x"74",
          2467 => x"d0",
          2468 => x"70",
          2469 => x"ec",
          2470 => x"58",
          2471 => x"06",
          2472 => x"08",
          2473 => x"34",
          2474 => x"39",
          2475 => x"f7",
          2476 => x"7d",
          2477 => x"df",
          2478 => x"05",
          2479 => x"33",
          2480 => x"82",
          2481 => x"ab",
          2482 => x"51",
          2483 => x"1a",
          2484 => x"81",
          2485 => x"70",
          2486 => x"51",
          2487 => x"81",
          2488 => x"34",
          2489 => x"34",
          2490 => x"25",
          2491 => x"f7",
          2492 => x"81",
          2493 => x"70",
          2494 => x"51",
          2495 => x"82",
          2496 => x"33",
          2497 => x"81",
          2498 => x"70",
          2499 => x"51",
          2500 => x"f7",
          2501 => x"2c",
          2502 => x"56",
          2503 => x"fb",
          2504 => x"a1",
          2505 => x"80",
          2506 => x"d8",
          2507 => x"de",
          2508 => x"80",
          2509 => x"53",
          2510 => x"9a",
          2511 => x"33",
          2512 => x"80",
          2513 => x"33",
          2514 => x"34",
          2515 => x"34",
          2516 => x"ff",
          2517 => x"70",
          2518 => x"d8",
          2519 => x"25",
          2520 => x"33",
          2521 => x"73",
          2522 => x"81",
          2523 => x"70",
          2524 => x"51",
          2525 => x"fb",
          2526 => x"f1",
          2527 => x"2b",
          2528 => x"57",
          2529 => x"bf",
          2530 => x"51",
          2531 => x"0a",
          2532 => x"2c",
          2533 => x"75",
          2534 => x"82",
          2535 => x"74",
          2536 => x"51",
          2537 => x"52",
          2538 => x"98",
          2539 => x"38",
          2540 => x"2e",
          2541 => x"51",
          2542 => x"34",
          2543 => x"0b",
          2544 => x"98",
          2545 => x"dc",
          2546 => x"38",
          2547 => x"ff",
          2548 => x"ff",
          2549 => x"73",
          2550 => x"f7",
          2551 => x"55",
          2552 => x"14",
          2553 => x"98",
          2554 => x"06",
          2555 => x"38",
          2556 => x"34",
          2557 => x"51",
          2558 => x"0a",
          2559 => x"2c",
          2560 => x"75",
          2561 => x"08",
          2562 => x"82",
          2563 => x"98",
          2564 => x"56",
          2565 => x"82",
          2566 => x"93",
          2567 => x"81",
          2568 => x"f7",
          2569 => x"25",
          2570 => x"dc",
          2571 => x"d8",
          2572 => x"f7",
          2573 => x"81",
          2574 => x"74",
          2575 => x"e9",
          2576 => x"ff",
          2577 => x"54",
          2578 => x"39",
          2579 => x"c1",
          2580 => x"82",
          2581 => x"d8",
          2582 => x"82",
          2583 => x"a6",
          2584 => x"82",
          2585 => x"82",
          2586 => x"05",
          2587 => x"bc",
          2588 => x"84",
          2589 => x"08",
          2590 => x"74",
          2591 => x"98",
          2592 => x"98",
          2593 => x"74",
          2594 => x"ff",
          2595 => x"55",
          2596 => x"51",
          2597 => x"93",
          2598 => x"df",
          2599 => x"38",
          2600 => x"e0",
          2601 => x"e0",
          2602 => x"53",
          2603 => x"3f",
          2604 => x"df",
          2605 => x"80",
          2606 => x"c4",
          2607 => x"d8",
          2608 => x"06",
          2609 => x"ff",
          2610 => x"81",
          2611 => x"f7",
          2612 => x"dc",
          2613 => x"51",
          2614 => x"f7",
          2615 => x"f7",
          2616 => x"27",
          2617 => x"52",
          2618 => x"34",
          2619 => x"90",
          2620 => x"dc",
          2621 => x"38",
          2622 => x"ff",
          2623 => x"ff",
          2624 => x"f4",
          2625 => x"f4",
          2626 => x"0b",
          2627 => x"53",
          2628 => x"a0",
          2629 => x"80",
          2630 => x"81",
          2631 => x"77",
          2632 => x"82",
          2633 => x"34",
          2634 => x"08",
          2635 => x"80",
          2636 => x"70",
          2637 => x"88",
          2638 => x"e0",
          2639 => x"88",
          2640 => x"77",
          2641 => x"89",
          2642 => x"52",
          2643 => x"fb",
          2644 => x"ff",
          2645 => x"e0",
          2646 => x"3d",
          2647 => x"05",
          2648 => x"88",
          2649 => x"83",
          2650 => x"33",
          2651 => x"ae",
          2652 => x"07",
          2653 => x"54",
          2654 => x"77",
          2655 => x"88",
          2656 => x"70",
          2657 => x"82",
          2658 => x"81",
          2659 => x"83",
          2660 => x"56",
          2661 => x"06",
          2662 => x"82",
          2663 => x"72",
          2664 => x"16",
          2665 => x"34",
          2666 => x"82",
          2667 => x"05",
          2668 => x"11",
          2669 => x"71",
          2670 => x"55",
          2671 => x"13",
          2672 => x"2a",
          2673 => x"34",
          2674 => x"08",
          2675 => x"33",
          2676 => x"56",
          2677 => x"33",
          2678 => x"70",
          2679 => x"86",
          2680 => x"e0",
          2681 => x"33",
          2682 => x"ff",
          2683 => x"53",
          2684 => x"34",
          2685 => x"02",
          2686 => x"71",
          2687 => x"12",
          2688 => x"29",
          2689 => x"98",
          2690 => x"53",
          2691 => x"71",
          2692 => x"fe",
          2693 => x"16",
          2694 => x"2b",
          2695 => x"33",
          2696 => x"70",
          2697 => x"52",
          2698 => x"05",
          2699 => x"13",
          2700 => x"88",
          2701 => x"33",
          2702 => x"56",
          2703 => x"81",
          2704 => x"81",
          2705 => x"51",
          2706 => x"81",
          2707 => x"3d",
          2708 => x"05",
          2709 => x"11",
          2710 => x"8b",
          2711 => x"59",
          2712 => x"81",
          2713 => x"8c",
          2714 => x"88",
          2715 => x"73",
          2716 => x"88",
          2717 => x"33",
          2718 => x"56",
          2719 => x"33",
          2720 => x"70",
          2721 => x"82",
          2722 => x"e0",
          2723 => x"12",
          2724 => x"98",
          2725 => x"f7",
          2726 => x"31",
          2727 => x"70",
          2728 => x"e0",
          2729 => x"82",
          2730 => x"2b",
          2731 => x"33",
          2732 => x"90",
          2733 => x"5b",
          2734 => x"8d",
          2735 => x"fe",
          2736 => x"33",
          2737 => x"83",
          2738 => x"53",
          2739 => x"34",
          2740 => x"14",
          2741 => x"84",
          2742 => x"2b",
          2743 => x"56",
          2744 => x"16",
          2745 => x"80",
          2746 => x"14",
          2747 => x"84",
          2748 => x"e0",
          2749 => x"33",
          2750 => x"80",
          2751 => x"56",
          2752 => x"34",
          2753 => x"73",
          2754 => x"f7",
          2755 => x"71",
          2756 => x"04",
          2757 => x"f8",
          2758 => x"ff",
          2759 => x"11",
          2760 => x"07",
          2761 => x"ff",
          2762 => x"38",
          2763 => x"12",
          2764 => x"ff",
          2765 => x"ff",
          2766 => x"56",
          2767 => x"73",
          2768 => x"5b",
          2769 => x"88",
          2770 => x"78",
          2771 => x"79",
          2772 => x"e0",
          2773 => x"33",
          2774 => x"ff",
          2775 => x"73",
          2776 => x"54",
          2777 => x"54",
          2778 => x"7a",
          2779 => x"51",
          2780 => x"80",
          2781 => x"c6",
          2782 => x"86",
          2783 => x"2b",
          2784 => x"55",
          2785 => x"ff",
          2786 => x"54",
          2787 => x"06",
          2788 => x"88",
          2789 => x"1e",
          2790 => x"88",
          2791 => x"5e",
          2792 => x"34",
          2793 => x"08",
          2794 => x"33",
          2795 => x"53",
          2796 => x"86",
          2797 => x"e0",
          2798 => x"11",
          2799 => x"07",
          2800 => x"56",
          2801 => x"16",
          2802 => x"05",
          2803 => x"3d",
          2804 => x"82",
          2805 => x"3f",
          2806 => x"71",
          2807 => x"08",
          2808 => x"3d",
          2809 => x"40",
          2810 => x"88",
          2811 => x"38",
          2812 => x"51",
          2813 => x"54",
          2814 => x"51",
          2815 => x"39",
          2816 => x"98",
          2817 => x"88",
          2818 => x"83",
          2819 => x"11",
          2820 => x"2b",
          2821 => x"ff",
          2822 => x"88",
          2823 => x"71",
          2824 => x"44",
          2825 => x"5b",
          2826 => x"25",
          2827 => x"75",
          2828 => x"54",
          2829 => x"88",
          2830 => x"33",
          2831 => x"90",
          2832 => x"54",
          2833 => x"31",
          2834 => x"77",
          2835 => x"54",
          2836 => x"38",
          2837 => x"ff",
          2838 => x"8e",
          2839 => x"51",
          2840 => x"18",
          2841 => x"79",
          2842 => x"71",
          2843 => x"f4",
          2844 => x"3f",
          2845 => x"06",
          2846 => x"82",
          2847 => x"55",
          2848 => x"88",
          2849 => x"ff",
          2850 => x"15",
          2851 => x"78",
          2852 => x"08",
          2853 => x"71",
          2854 => x"9c",
          2855 => x"3f",
          2856 => x"06",
          2857 => x"82",
          2858 => x"55",
          2859 => x"88",
          2860 => x"19",
          2861 => x"58",
          2862 => x"b0",
          2863 => x"e0",
          2864 => x"53",
          2865 => x"ff",
          2866 => x"3f",
          2867 => x"80",
          2868 => x"3f",
          2869 => x"08",
          2870 => x"7b",
          2871 => x"3d",
          2872 => x"29",
          2873 => x"e0",
          2874 => x"80",
          2875 => x"82",
          2876 => x"3f",
          2877 => x"0d",
          2878 => x"33",
          2879 => x"38",
          2880 => x"82",
          2881 => x"fc",
          2882 => x"84",
          2883 => x"51",
          2884 => x"84",
          2885 => x"51",
          2886 => x"81",
          2887 => x"92",
          2888 => x"0b",
          2889 => x"71",
          2890 => x"80",
          2891 => x"08",
          2892 => x"80",
          2893 => x"c0",
          2894 => x"87",
          2895 => x"82",
          2896 => x"e0",
          2897 => x"3d",
          2898 => x"bf",
          2899 => x"74",
          2900 => x"98",
          2901 => x"81",
          2902 => x"87",
          2903 => x"8c",
          2904 => x"5a",
          2905 => x"c0",
          2906 => x"76",
          2907 => x"81",
          2908 => x"8e",
          2909 => x"81",
          2910 => x"74",
          2911 => x"83",
          2912 => x"8f",
          2913 => x"c0",
          2914 => x"87",
          2915 => x"2e",
          2916 => x"38",
          2917 => x"15",
          2918 => x"52",
          2919 => x"39",
          2920 => x"ff",
          2921 => x"90",
          2922 => x"71",
          2923 => x"38",
          2924 => x"80",
          2925 => x"72",
          2926 => x"04",
          2927 => x"8c",
          2928 => x"5b",
          2929 => x"e1",
          2930 => x"79",
          2931 => x"06",
          2932 => x"87",
          2933 => x"8c",
          2934 => x"59",
          2935 => x"98",
          2936 => x"0c",
          2937 => x"70",
          2938 => x"2e",
          2939 => x"33",
          2940 => x"2a",
          2941 => x"2e",
          2942 => x"52",
          2943 => x"08",
          2944 => x"84",
          2945 => x"87",
          2946 => x"70",
          2947 => x"ff",
          2948 => x"81",
          2949 => x"52",
          2950 => x"80",
          2951 => x"7a",
          2952 => x"80",
          2953 => x"81",
          2954 => x"0c",
          2955 => x"7a",
          2956 => x"88",
          2957 => x"56",
          2958 => x"08",
          2959 => x"fe",
          2960 => x"0c",
          2961 => x"38",
          2962 => x"2b",
          2963 => x"71",
          2964 => x"71",
          2965 => x"39",
          2966 => x"06",
          2967 => x"38",
          2968 => x"e8",
          2969 => x"71",
          2970 => x"92",
          2971 => x"06",
          2972 => x"80",
          2973 => x"0c",
          2974 => x"56",
          2975 => x"82",
          2976 => x"fe",
          2977 => x"33",
          2978 => x"0c",
          2979 => x"3d",
          2980 => x"33",
          2981 => x"81",
          2982 => x"75",
          2983 => x"52",
          2984 => x"0d",
          2985 => x"05",
          2986 => x"70",
          2987 => x"51",
          2988 => x"ff",
          2989 => x"72",
          2990 => x"2a",
          2991 => x"34",
          2992 => x"81",
          2993 => x"70",
          2994 => x"3d",
          2995 => x"70",
          2996 => x"05",
          2997 => x"34",
          2998 => x"0d",
          2999 => x"54",
          3000 => x"54",
          3001 => x"84",
          3002 => x"77",
          3003 => x"05",
          3004 => x"33",
          3005 => x"52",
          3006 => x"80",
          3007 => x"0c",
          3008 => x"74",
          3009 => x"2e",
          3010 => x"52",
          3011 => x"98",
          3012 => x"82",
          3013 => x"77",
          3014 => x"33",
          3015 => x"ff",
          3016 => x"72",
          3017 => x"72",
          3018 => x"98",
          3019 => x"80",
          3020 => x"55",
          3021 => x"0d",
          3022 => x"0b",
          3023 => x"2e",
          3024 => x"08",
          3025 => x"33",
          3026 => x"98",
          3027 => x"38",
          3028 => x"b4",
          3029 => x"a0",
          3030 => x"27",
          3031 => x"82",
          3032 => x"54",
          3033 => x"33",
          3034 => x"5a",
          3035 => x"0d",
          3036 => x"56",
          3037 => x"af",
          3038 => x"e0",
          3039 => x"9f",
          3040 => x"52",
          3041 => x"82",
          3042 => x"ff",
          3043 => x"76",
          3044 => x"04",
          3045 => x"fe",
          3046 => x"82",
          3047 => x"33",
          3048 => x"80",
          3049 => x"81",
          3050 => x"84",
          3051 => x"b8",
          3052 => x"82",
          3053 => x"fb",
          3054 => x"52",
          3055 => x"85",
          3056 => x"fb",
          3057 => x"a0",
          3058 => x"08",
          3059 => x"3f",
          3060 => x"19",
          3061 => x"17",
          3062 => x"18",
          3063 => x"33",
          3064 => x"08",
          3065 => x"82",
          3066 => x"fb",
          3067 => x"08",
          3068 => x"74",
          3069 => x"75",
          3070 => x"53",
          3071 => x"0d",
          3072 => x"08",
          3073 => x"df",
          3074 => x"d7",
          3075 => x"82",
          3076 => x"89",
          3077 => x"bf",
          3078 => x"81",
          3079 => x"89",
          3080 => x"52",
          3081 => x"08",
          3082 => x"14",
          3083 => x"2a",
          3084 => x"57",
          3085 => x"98",
          3086 => x"06",
          3087 => x"78",
          3088 => x"5c",
          3089 => x"38",
          3090 => x"39",
          3091 => x"52",
          3092 => x"98",
          3093 => x"fe",
          3094 => x"cf",
          3095 => x"ff",
          3096 => x"a8",
          3097 => x"91",
          3098 => x"76",
          3099 => x"b8",
          3100 => x"98",
          3101 => x"81",
          3102 => x"3d",
          3103 => x"7e",
          3104 => x"27",
          3105 => x"27",
          3106 => x"79",
          3107 => x"89",
          3108 => x"80",
          3109 => x"81",
          3110 => x"89",
          3111 => x"52",
          3112 => x"08",
          3113 => x"38",
          3114 => x"81",
          3115 => x"77",
          3116 => x"84",
          3117 => x"06",
          3118 => x"81",
          3119 => x"a8",
          3120 => x"d9",
          3121 => x"e0",
          3122 => x"ff",
          3123 => x"54",
          3124 => x"74",
          3125 => x"07",
          3126 => x"39",
          3127 => x"52",
          3128 => x"98",
          3129 => x"d8",
          3130 => x"76",
          3131 => x"05",
          3132 => x"87",
          3133 => x"51",
          3134 => x"59",
          3135 => x"f0",
          3136 => x"06",
          3137 => x"54",
          3138 => x"08",
          3139 => x"51",
          3140 => x"34",
          3141 => x"0d",
          3142 => x"72",
          3143 => x"27",
          3144 => x"9d",
          3145 => x"53",
          3146 => x"82",
          3147 => x"08",
          3148 => x"80",
          3149 => x"82",
          3150 => x"74",
          3151 => x"e0",
          3152 => x"80",
          3153 => x"08",
          3154 => x"08",
          3155 => x"52",
          3156 => x"98",
          3157 => x"11",
          3158 => x"74",
          3159 => x"0c",
          3160 => x"84",
          3161 => x"ff",
          3162 => x"98",
          3163 => x"0d",
          3164 => x"79",
          3165 => x"80",
          3166 => x"26",
          3167 => x"52",
          3168 => x"74",
          3169 => x"38",
          3170 => x"98",
          3171 => x"17",
          3172 => x"c7",
          3173 => x"56",
          3174 => x"77",
          3175 => x"38",
          3176 => x"26",
          3177 => x"51",
          3178 => x"98",
          3179 => x"38",
          3180 => x"98",
          3181 => x"80",
          3182 => x"08",
          3183 => x"ef",
          3184 => x"95",
          3185 => x"27",
          3186 => x"89",
          3187 => x"db",
          3188 => x"17",
          3189 => x"75",
          3190 => x"7a",
          3191 => x"08",
          3192 => x"e0",
          3193 => x"86",
          3194 => x"e0",
          3195 => x"07",
          3196 => x"55",
          3197 => x"2e",
          3198 => x"55",
          3199 => x"76",
          3200 => x"08",
          3201 => x"e0",
          3202 => x"55",
          3203 => x"2e",
          3204 => x"51",
          3205 => x"55",
          3206 => x"9c",
          3207 => x"56",
          3208 => x"15",
          3209 => x"07",
          3210 => x"ff",
          3211 => x"39",
          3212 => x"08",
          3213 => x"74",
          3214 => x"04",
          3215 => x"f3",
          3216 => x"81",
          3217 => x"38",
          3218 => x"82",
          3219 => x"b4",
          3220 => x"52",
          3221 => x"3f",
          3222 => x"8a",
          3223 => x"38",
          3224 => x"81",
          3225 => x"e0",
          3226 => x"15",
          3227 => x"07",
          3228 => x"75",
          3229 => x"04",
          3230 => x"58",
          3231 => x"80",
          3232 => x"80",
          3233 => x"17",
          3234 => x"53",
          3235 => x"08",
          3236 => x"53",
          3237 => x"72",
          3238 => x"08",
          3239 => x"16",
          3240 => x"75",
          3241 => x"f5",
          3242 => x"82",
          3243 => x"81",
          3244 => x"38",
          3245 => x"26",
          3246 => x"73",
          3247 => x"51",
          3248 => x"98",
          3249 => x"17",
          3250 => x"9a",
          3251 => x"74",
          3252 => x"83",
          3253 => x"0c",
          3254 => x"8a",
          3255 => x"70",
          3256 => x"57",
          3257 => x"38",
          3258 => x"08",
          3259 => x"cb",
          3260 => x"81",
          3261 => x"94",
          3262 => x"85",
          3263 => x"73",
          3264 => x"8a",
          3265 => x"06",
          3266 => x"73",
          3267 => x"08",
          3268 => x"98",
          3269 => x"82",
          3270 => x"38",
          3271 => x"26",
          3272 => x"98",
          3273 => x"94",
          3274 => x"3f",
          3275 => x"82",
          3276 => x"38",
          3277 => x"2e",
          3278 => x"08",
          3279 => x"08",
          3280 => x"e0",
          3281 => x"0c",
          3282 => x"82",
          3283 => x"90",
          3284 => x"15",
          3285 => x"0c",
          3286 => x"7b",
          3287 => x"52",
          3288 => x"98",
          3289 => x"ec",
          3290 => x"17",
          3291 => x"82",
          3292 => x"08",
          3293 => x"9c",
          3294 => x"72",
          3295 => x"38",
          3296 => x"72",
          3297 => x"53",
          3298 => x"56",
          3299 => x"38",
          3300 => x"81",
          3301 => x"e0",
          3302 => x"80",
          3303 => x"09",
          3304 => x"82",
          3305 => x"fd",
          3306 => x"eb",
          3307 => x"ff",
          3308 => x"53",
          3309 => x"38",
          3310 => x"e0",
          3311 => x"72",
          3312 => x"04",
          3313 => x"ff",
          3314 => x"55",
          3315 => x"53",
          3316 => x"38",
          3317 => x"eb",
          3318 => x"3d",
          3319 => x"70",
          3320 => x"74",
          3321 => x"70",
          3322 => x"51",
          3323 => x"98",
          3324 => x"0d",
          3325 => x"5f",
          3326 => x"19",
          3327 => x"19",
          3328 => x"82",
          3329 => x"08",
          3330 => x"33",
          3331 => x"82",
          3332 => x"70",
          3333 => x"1a",
          3334 => x"81",
          3335 => x"81",
          3336 => x"ae",
          3337 => x"53",
          3338 => x"82",
          3339 => x"56",
          3340 => x"38",
          3341 => x"81",
          3342 => x"2e",
          3343 => x"86",
          3344 => x"80",
          3345 => x"81",
          3346 => x"1d",
          3347 => x"09",
          3348 => x"33",
          3349 => x"81",
          3350 => x"52",
          3351 => x"08",
          3352 => x"f8",
          3353 => x"8d",
          3354 => x"58",
          3355 => x"05",
          3356 => x"08",
          3357 => x"2e",
          3358 => x"c8",
          3359 => x"75",
          3360 => x"75",
          3361 => x"b0",
          3362 => x"c1",
          3363 => x"81",
          3364 => x"8e",
          3365 => x"73",
          3366 => x"1c",
          3367 => x"39",
          3368 => x"7b",
          3369 => x"82",
          3370 => x"72",
          3371 => x"1a",
          3372 => x"f8",
          3373 => x"82",
          3374 => x"08",
          3375 => x"98",
          3376 => x"90",
          3377 => x"70",
          3378 => x"f6",
          3379 => x"82",
          3380 => x"ff",
          3381 => x"0c",
          3382 => x"a9",
          3383 => x"e0",
          3384 => x"08",
          3385 => x"84",
          3386 => x"bf",
          3387 => x"73",
          3388 => x"82",
          3389 => x"06",
          3390 => x"73",
          3391 => x"81",
          3392 => x"70",
          3393 => x"55",
          3394 => x"70",
          3395 => x"92",
          3396 => x"06",
          3397 => x"58",
          3398 => x"06",
          3399 => x"7d",
          3400 => x"38",
          3401 => x"e5",
          3402 => x"ff",
          3403 => x"76",
          3404 => x"05",
          3405 => x"d2",
          3406 => x"8f",
          3407 => x"ff",
          3408 => x"77",
          3409 => x"51",
          3410 => x"08",
          3411 => x"81",
          3412 => x"74",
          3413 => x"06",
          3414 => x"75",
          3415 => x"b3",
          3416 => x"ff",
          3417 => x"70",
          3418 => x"2e",
          3419 => x"77",
          3420 => x"8b",
          3421 => x"51",
          3422 => x"5c",
          3423 => x"f9",
          3424 => x"ff",
          3425 => x"ab",
          3426 => x"38",
          3427 => x"08",
          3428 => x"08",
          3429 => x"ff",
          3430 => x"51",
          3431 => x"58",
          3432 => x"e8",
          3433 => x"3d",
          3434 => x"08",
          3435 => x"5d",
          3436 => x"73",
          3437 => x"5d",
          3438 => x"70",
          3439 => x"f0",
          3440 => x"92",
          3441 => x"3f",
          3442 => x"54",
          3443 => x"c0",
          3444 => x"1c",
          3445 => x"52",
          3446 => x"27",
          3447 => x"70",
          3448 => x"80",
          3449 => x"06",
          3450 => x"81",
          3451 => x"71",
          3452 => x"56",
          3453 => x"84",
          3454 => x"76",
          3455 => x"55",
          3456 => x"57",
          3457 => x"74",
          3458 => x"76",
          3459 => x"2a",
          3460 => x"3d",
          3461 => x"34",
          3462 => x"54",
          3463 => x"70",
          3464 => x"e0",
          3465 => x"17",
          3466 => x"15",
          3467 => x"89",
          3468 => x"d0",
          3469 => x"54",
          3470 => x"56",
          3471 => x"81",
          3472 => x"78",
          3473 => x"51",
          3474 => x"8b",
          3475 => x"27",
          3476 => x"e4",
          3477 => x"08",
          3478 => x"09",
          3479 => x"cb",
          3480 => x"cb",
          3481 => x"06",
          3482 => x"2e",
          3483 => x"fe",
          3484 => x"19",
          3485 => x"3f",
          3486 => x"98",
          3487 => x"78",
          3488 => x"2b",
          3489 => x"79",
          3490 => x"08",
          3491 => x"38",
          3492 => x"e0",
          3493 => x"1a",
          3494 => x"82",
          3495 => x"08",
          3496 => x"1b",
          3497 => x"5b",
          3498 => x"17",
          3499 => x"34",
          3500 => x"51",
          3501 => x"05",
          3502 => x"2e",
          3503 => x"81",
          3504 => x"d2",
          3505 => x"b9",
          3506 => x"54",
          3507 => x"38",
          3508 => x"74",
          3509 => x"86",
          3510 => x"76",
          3511 => x"52",
          3512 => x"98",
          3513 => x"c9",
          3514 => x"38",
          3515 => x"81",
          3516 => x"e0",
          3517 => x"e0",
          3518 => x"df",
          3519 => x"9c",
          3520 => x"1a",
          3521 => x"55",
          3522 => x"1d",
          3523 => x"0c",
          3524 => x"78",
          3525 => x"08",
          3526 => x"94",
          3527 => x"3f",
          3528 => x"98",
          3529 => x"52",
          3530 => x"98",
          3531 => x"38",
          3532 => x"81",
          3533 => x"77",
          3534 => x"52",
          3535 => x"98",
          3536 => x"2e",
          3537 => x"06",
          3538 => x"98",
          3539 => x"0d",
          3540 => x"80",
          3541 => x"80",
          3542 => x"ff",
          3543 => x"7f",
          3544 => x"5b",
          3545 => x"38",
          3546 => x"5b",
          3547 => x"80",
          3548 => x"53",
          3549 => x"5b",
          3550 => x"81",
          3551 => x"b5",
          3552 => x"80",
          3553 => x"83",
          3554 => x"27",
          3555 => x"74",
          3556 => x"97",
          3557 => x"30",
          3558 => x"72",
          3559 => x"80",
          3560 => x"74",
          3561 => x"80",
          3562 => x"70",
          3563 => x"38",
          3564 => x"79",
          3565 => x"05",
          3566 => x"70",
          3567 => x"08",
          3568 => x"53",
          3569 => x"2e",
          3570 => x"55",
          3571 => x"07",
          3572 => x"26",
          3573 => x"ae",
          3574 => x"17",
          3575 => x"34",
          3576 => x"b5",
          3577 => x"0b",
          3578 => x"72",
          3579 => x"0b",
          3580 => x"39",
          3581 => x"57",
          3582 => x"18",
          3583 => x"bf",
          3584 => x"38",
          3585 => x"53",
          3586 => x"2a",
          3587 => x"72",
          3588 => x"38",
          3589 => x"56",
          3590 => x"34",
          3591 => x"33",
          3592 => x"38",
          3593 => x"82",
          3594 => x"33",
          3595 => x"19",
          3596 => x"33",
          3597 => x"11",
          3598 => x"98",
          3599 => x"87",
          3600 => x"23",
          3601 => x"e0",
          3602 => x"0d",
          3603 => x"41",
          3604 => x"55",
          3605 => x"73",
          3606 => x"2e",
          3607 => x"1f",
          3608 => x"64",
          3609 => x"2e",
          3610 => x"73",
          3611 => x"25",
          3612 => x"38",
          3613 => x"51",
          3614 => x"80",
          3615 => x"51",
          3616 => x"56",
          3617 => x"8c",
          3618 => x"3d",
          3619 => x"e0",
          3620 => x"83",
          3621 => x"27",
          3622 => x"98",
          3623 => x"23",
          3624 => x"83",
          3625 => x"30",
          3626 => x"51",
          3627 => x"80",
          3628 => x"26",
          3629 => x"51",
          3630 => x"81",
          3631 => x"d7",
          3632 => x"23",
          3633 => x"15",
          3634 => x"57",
          3635 => x"38",
          3636 => x"30",
          3637 => x"54",
          3638 => x"27",
          3639 => x"81",
          3640 => x"ae",
          3641 => x"82",
          3642 => x"82",
          3643 => x"81",
          3644 => x"73",
          3645 => x"78",
          3646 => x"0b",
          3647 => x"78",
          3648 => x"70",
          3649 => x"8a",
          3650 => x"54",
          3651 => x"78",
          3652 => x"fe",
          3653 => x"72",
          3654 => x"51",
          3655 => x"2e",
          3656 => x"59",
          3657 => x"55",
          3658 => x"86",
          3659 => x"57",
          3660 => x"83",
          3661 => x"a0",
          3662 => x"1d",
          3663 => x"5d",
          3664 => x"38",
          3665 => x"ae",
          3666 => x"83",
          3667 => x"79",
          3668 => x"73",
          3669 => x"fe",
          3670 => x"2e",
          3671 => x"55",
          3672 => x"38",
          3673 => x"d5",
          3674 => x"5f",
          3675 => x"5f",
          3676 => x"38",
          3677 => x"32",
          3678 => x"54",
          3679 => x"2e",
          3680 => x"39",
          3681 => x"83",
          3682 => x"30",
          3683 => x"07",
          3684 => x"a6",
          3685 => x"7c",
          3686 => x"57",
          3687 => x"5d",
          3688 => x"fc",
          3689 => x"ff",
          3690 => x"57",
          3691 => x"ae",
          3692 => x"ff",
          3693 => x"51",
          3694 => x"75",
          3695 => x"33",
          3696 => x"38",
          3697 => x"38",
          3698 => x"c0",
          3699 => x"2a",
          3700 => x"58",
          3701 => x"38",
          3702 => x"cc",
          3703 => x"8a",
          3704 => x"56",
          3705 => x"99",
          3706 => x"ff",
          3707 => x"38",
          3708 => x"ff",
          3709 => x"a0",
          3710 => x"58",
          3711 => x"73",
          3712 => x"38",
          3713 => x"2e",
          3714 => x"2b",
          3715 => x"54",
          3716 => x"06",
          3717 => x"85",
          3718 => x"2a",
          3719 => x"38",
          3720 => x"85",
          3721 => x"2a",
          3722 => x"2e",
          3723 => x"ab",
          3724 => x"82",
          3725 => x"56",
          3726 => x"38",
          3727 => x"81",
          3728 => x"70",
          3729 => x"54",
          3730 => x"06",
          3731 => x"ff",
          3732 => x"80",
          3733 => x"bb",
          3734 => x"2a",
          3735 => x"38",
          3736 => x"81",
          3737 => x"e1",
          3738 => x"60",
          3739 => x"ef",
          3740 => x"0c",
          3741 => x"0c",
          3742 => x"7c",
          3743 => x"55",
          3744 => x"81",
          3745 => x"33",
          3746 => x"2e",
          3747 => x"2e",
          3748 => x"33",
          3749 => x"52",
          3750 => x"14",
          3751 => x"52",
          3752 => x"0b",
          3753 => x"7a",
          3754 => x"33",
          3755 => x"9f",
          3756 => x"89",
          3757 => x"54",
          3758 => x"26",
          3759 => x"06",
          3760 => x"51",
          3761 => x"85",
          3762 => x"74",
          3763 => x"9f",
          3764 => x"54",
          3765 => x"15",
          3766 => x"ff",
          3767 => x"86",
          3768 => x"51",
          3769 => x"70",
          3770 => x"04",
          3771 => x"83",
          3772 => x"79",
          3773 => x"55",
          3774 => x"84",
          3775 => x"e0",
          3776 => x"83",
          3777 => x"81",
          3778 => x"17",
          3779 => x"09",
          3780 => x"81",
          3781 => x"79",
          3782 => x"74",
          3783 => x"38",
          3784 => x"ee",
          3785 => x"98",
          3786 => x"2e",
          3787 => x"52",
          3788 => x"82",
          3789 => x"08",
          3790 => x"82",
          3791 => x"f2",
          3792 => x"cb",
          3793 => x"60",
          3794 => x"08",
          3795 => x"98",
          3796 => x"98",
          3797 => x"70",
          3798 => x"2e",
          3799 => x"81",
          3800 => x"80",
          3801 => x"c6",
          3802 => x"ff",
          3803 => x"98",
          3804 => x"74",
          3805 => x"8a",
          3806 => x"39",
          3807 => x"e0",
          3808 => x"52",
          3809 => x"82",
          3810 => x"81",
          3811 => x"cb",
          3812 => x"82",
          3813 => x"56",
          3814 => x"74",
          3815 => x"98",
          3816 => x"2e",
          3817 => x"38",
          3818 => x"7b",
          3819 => x"56",
          3820 => x"70",
          3821 => x"83",
          3822 => x"e0",
          3823 => x"05",
          3824 => x"56",
          3825 => x"82",
          3826 => x"9f",
          3827 => x"84",
          3828 => x"55",
          3829 => x"7a",
          3830 => x"51",
          3831 => x"81",
          3832 => x"8d",
          3833 => x"09",
          3834 => x"77",
          3835 => x"38",
          3836 => x"76",
          3837 => x"2e",
          3838 => x"26",
          3839 => x"ca",
          3840 => x"ff",
          3841 => x"09",
          3842 => x"14",
          3843 => x"08",
          3844 => x"38",
          3845 => x"82",
          3846 => x"0c",
          3847 => x"80",
          3848 => x"ff",
          3849 => x"81",
          3850 => x"06",
          3851 => x"52",
          3852 => x"80",
          3853 => x"53",
          3854 => x"83",
          3855 => x"87",
          3856 => x"e0",
          3857 => x"06",
          3858 => x"80",
          3859 => x"e0",
          3860 => x"74",
          3861 => x"ee",
          3862 => x"c6",
          3863 => x"98",
          3864 => x"56",
          3865 => x"14",
          3866 => x"5a",
          3867 => x"8a",
          3868 => x"fe",
          3869 => x"55",
          3870 => x"f3",
          3871 => x"ff",
          3872 => x"74",
          3873 => x"57",
          3874 => x"57",
          3875 => x"82",
          3876 => x"0c",
          3877 => x"a8",
          3878 => x"54",
          3879 => x"af",
          3880 => x"3f",
          3881 => x"06",
          3882 => x"79",
          3883 => x"c7",
          3884 => x"15",
          3885 => x"8d",
          3886 => x"77",
          3887 => x"76",
          3888 => x"70",
          3889 => x"53",
          3890 => x"56",
          3891 => x"38",
          3892 => x"90",
          3893 => x"34",
          3894 => x"92",
          3895 => x"3f",
          3896 => x"06",
          3897 => x"80",
          3898 => x"ca",
          3899 => x"ea",
          3900 => x"34",
          3901 => x"82",
          3902 => x"53",
          3903 => x"06",
          3904 => x"96",
          3905 => x"85",
          3906 => x"38",
          3907 => x"82",
          3908 => x"f2",
          3909 => x"a0",
          3910 => x"98",
          3911 => x"51",
          3912 => x"90",
          3913 => x"f0",
          3914 => x"f0",
          3915 => x"f8",
          3916 => x"15",
          3917 => x"0c",
          3918 => x"77",
          3919 => x"38",
          3920 => x"38",
          3921 => x"38",
          3922 => x"52",
          3923 => x"38",
          3924 => x"3f",
          3925 => x"71",
          3926 => x"83",
          3927 => x"52",
          3928 => x"0d",
          3929 => x"33",
          3930 => x"56",
          3931 => x"82",
          3932 => x"e0",
          3933 => x"05",
          3934 => x"84",
          3935 => x"80",
          3936 => x"75",
          3937 => x"38",
          3938 => x"05",
          3939 => x"08",
          3940 => x"3d",
          3941 => x"84",
          3942 => x"89",
          3943 => x"77",
          3944 => x"05",
          3945 => x"f6",
          3946 => x"82",
          3947 => x"5c",
          3948 => x"ea",
          3949 => x"82",
          3950 => x"d7",
          3951 => x"73",
          3952 => x"9c",
          3953 => x"38",
          3954 => x"2e",
          3955 => x"df",
          3956 => x"9e",
          3957 => x"54",
          3958 => x"70",
          3959 => x"8e",
          3960 => x"88",
          3961 => x"83",
          3962 => x"80",
          3963 => x"51",
          3964 => x"56",
          3965 => x"05",
          3966 => x"0b",
          3967 => x"7a",
          3968 => x"9c",
          3969 => x"81",
          3970 => x"80",
          3971 => x"54",
          3972 => x"05",
          3973 => x"08",
          3974 => x"38",
          3975 => x"b2",
          3976 => x"06",
          3977 => x"38",
          3978 => x"2a",
          3979 => x"2e",
          3980 => x"80",
          3981 => x"39",
          3982 => x"82",
          3983 => x"12",
          3984 => x"81",
          3985 => x"06",
          3986 => x"77",
          3987 => x"08",
          3988 => x"63",
          3989 => x"82",
          3990 => x"88",
          3991 => x"c0",
          3992 => x"e0",
          3993 => x"0c",
          3994 => x"77",
          3995 => x"34",
          3996 => x"94",
          3997 => x"06",
          3998 => x"38",
          3999 => x"84",
          4000 => x"0c",
          4001 => x"52",
          4002 => x"51",
          4003 => x"57",
          4004 => x"38",
          4005 => x"2e",
          4006 => x"75",
          4007 => x"07",
          4008 => x"8a",
          4009 => x"73",
          4010 => x"a9",
          4011 => x"80",
          4012 => x"c4",
          4013 => x"38",
          4014 => x"82",
          4015 => x"84",
          4016 => x"82",
          4017 => x"f2",
          4018 => x"40",
          4019 => x"fc",
          4020 => x"82",
          4021 => x"08",
          4022 => x"80",
          4023 => x"39",
          4024 => x"56",
          4025 => x"39",
          4026 => x"82",
          4027 => x"81",
          4028 => x"94",
          4029 => x"83",
          4030 => x"8c",
          4031 => x"06",
          4032 => x"8a",
          4033 => x"06",
          4034 => x"38",
          4035 => x"19",
          4036 => x"82",
          4037 => x"ff",
          4038 => x"38",
          4039 => x"52",
          4040 => x"98",
          4041 => x"e0",
          4042 => x"57",
          4043 => x"1a",
          4044 => x"75",
          4045 => x"58",
          4046 => x"1b",
          4047 => x"e0",
          4048 => x"11",
          4049 => x"38",
          4050 => x"78",
          4051 => x"16",
          4052 => x"2b",
          4053 => x"77",
          4054 => x"1a",
          4055 => x"84",
          4056 => x"27",
          4057 => x"52",
          4058 => x"98",
          4059 => x"19",
          4060 => x"52",
          4061 => x"76",
          4062 => x"1e",
          4063 => x"5e",
          4064 => x"82",
          4065 => x"f2",
          4066 => x"40",
          4067 => x"fc",
          4068 => x"82",
          4069 => x"08",
          4070 => x"80",
          4071 => x"39",
          4072 => x"81",
          4073 => x"80",
          4074 => x"0b",
          4075 => x"39",
          4076 => x"83",
          4077 => x"56",
          4078 => x"09",
          4079 => x"94",
          4080 => x"56",
          4081 => x"22",
          4082 => x"55",
          4083 => x"18",
          4084 => x"85",
          4085 => x"c6",
          4086 => x"82",
          4087 => x"38",
          4088 => x"ff",
          4089 => x"0c",
          4090 => x"19",
          4091 => x"19",
          4092 => x"74",
          4093 => x"98",
          4094 => x"52",
          4095 => x"e0",
          4096 => x"82",
          4097 => x"5a",
          4098 => x"78",
          4099 => x"55",
          4100 => x"31",
          4101 => x"81",
          4102 => x"82",
          4103 => x"b4",
          4104 => x"79",
          4105 => x"16",
          4106 => x"52",
          4107 => x"7e",
          4108 => x"89",
          4109 => x"08",
          4110 => x"51",
          4111 => x"08",
          4112 => x"0c",
          4113 => x"08",
          4114 => x"57",
          4115 => x"56",
          4116 => x"bc",
          4117 => x"b0",
          4118 => x"08",
          4119 => x"ff",
          4120 => x"83",
          4121 => x"17",
          4122 => x"18",
          4123 => x"58",
          4124 => x"38",
          4125 => x"89",
          4126 => x"55",
          4127 => x"82",
          4128 => x"f8",
          4129 => x"53",
          4130 => x"e0",
          4131 => x"81",
          4132 => x"2a",
          4133 => x"80",
          4134 => x"52",
          4135 => x"e0",
          4136 => x"80",
          4137 => x"33",
          4138 => x"34",
          4139 => x"08",
          4140 => x"52",
          4141 => x"82",
          4142 => x"ff",
          4143 => x"51",
          4144 => x"0b",
          4145 => x"98",
          4146 => x"33",
          4147 => x"17",
          4148 => x"3d",
          4149 => x"52",
          4150 => x"08",
          4151 => x"86",
          4152 => x"ac",
          4153 => x"e0",
          4154 => x"08",
          4155 => x"86",
          4156 => x"3d",
          4157 => x"0b",
          4158 => x"82",
          4159 => x"80",
          4160 => x"3d",
          4161 => x"94",
          4162 => x"e8",
          4163 => x"82",
          4164 => x"58",
          4165 => x"dc",
          4166 => x"82",
          4167 => x"c7",
          4168 => x"73",
          4169 => x"12",
          4170 => x"33",
          4171 => x"55",
          4172 => x"7f",
          4173 => x"82",
          4174 => x"39",
          4175 => x"81",
          4176 => x"e0",
          4177 => x"a3",
          4178 => x"e1",
          4179 => x"80",
          4180 => x"52",
          4181 => x"82",
          4182 => x"08",
          4183 => x"0c",
          4184 => x"3d",
          4185 => x"54",
          4186 => x"52",
          4187 => x"90",
          4188 => x"e0",
          4189 => x"3d",
          4190 => x"3f",
          4191 => x"98",
          4192 => x"08",
          4193 => x"e0",
          4194 => x"52",
          4195 => x"98",
          4196 => x"b3",
          4197 => x"3f",
          4198 => x"98",
          4199 => x"52",
          4200 => x"e0",
          4201 => x"74",
          4202 => x"08",
          4203 => x"c9",
          4204 => x"86",
          4205 => x"81",
          4206 => x"05",
          4207 => x"93",
          4208 => x"56",
          4209 => x"02",
          4210 => x"16",
          4211 => x"38",
          4212 => x"99",
          4213 => x"16",
          4214 => x"3d",
          4215 => x"58",
          4216 => x"eb",
          4217 => x"11",
          4218 => x"39",
          4219 => x"38",
          4220 => x"55",
          4221 => x"f7",
          4222 => x"98",
          4223 => x"56",
          4224 => x"81",
          4225 => x"56",
          4226 => x"78",
          4227 => x"27",
          4228 => x"7a",
          4229 => x"55",
          4230 => x"5c",
          4231 => x"85",
          4232 => x"3d",
          4233 => x"33",
          4234 => x"78",
          4235 => x"82",
          4236 => x"04",
          4237 => x"fc",
          4238 => x"fc",
          4239 => x"e0",
          4240 => x"33",
          4241 => x"08",
          4242 => x"15",
          4243 => x"51",
          4244 => x"94",
          4245 => x"0c",
          4246 => x"79",
          4247 => x"51",
          4248 => x"52",
          4249 => x"82",
          4250 => x"70",
          4251 => x"82",
          4252 => x"76",
          4253 => x"0c",
          4254 => x"58",
          4255 => x"54",
          4256 => x"ff",
          4257 => x"54",
          4258 => x"9d",
          4259 => x"81",
          4260 => x"16",
          4261 => x"2e",
          4262 => x"de",
          4263 => x"18",
          4264 => x"81",
          4265 => x"56",
          4266 => x"74",
          4267 => x"98",
          4268 => x"38",
          4269 => x"73",
          4270 => x"82",
          4271 => x"bf",
          4272 => x"53",
          4273 => x"73",
          4274 => x"15",
          4275 => x"ff",
          4276 => x"73",
          4277 => x"82",
          4278 => x"91",
          4279 => x"81",
          4280 => x"39",
          4281 => x"05",
          4282 => x"08",
          4283 => x"0c",
          4284 => x"72",
          4285 => x"53",
          4286 => x"16",
          4287 => x"0c",
          4288 => x"8b",
          4289 => x"56",
          4290 => x"38",
          4291 => x"8a",
          4292 => x"82",
          4293 => x"08",
          4294 => x"52",
          4295 => x"98",
          4296 => x"c4",
          4297 => x"55",
          4298 => x"16",
          4299 => x"51",
          4300 => x"9c",
          4301 => x"3f",
          4302 => x"77",
          4303 => x"74",
          4304 => x"82",
          4305 => x"09",
          4306 => x"39",
          4307 => x"0c",
          4308 => x"89",
          4309 => x"87",
          4310 => x"e7",
          4311 => x"38",
          4312 => x"3d",
          4313 => x"89",
          4314 => x"54",
          4315 => x"53",
          4316 => x"74",
          4317 => x"73",
          4318 => x"98",
          4319 => x"98",
          4320 => x"82",
          4321 => x"08",
          4322 => x"80",
          4323 => x"a7",
          4324 => x"3f",
          4325 => x"3f",
          4326 => x"30",
          4327 => x"e0",
          4328 => x"72",
          4329 => x"04",
          4330 => x"89",
          4331 => x"de",
          4332 => x"82",
          4333 => x"75",
          4334 => x"08",
          4335 => x"02",
          4336 => x"55",
          4337 => x"55",
          4338 => x"76",
          4339 => x"82",
          4340 => x"f0",
          4341 => x"53",
          4342 => x"51",
          4343 => x"5b",
          4344 => x"7c",
          4345 => x"fe",
          4346 => x"55",
          4347 => x"0c",
          4348 => x"39",
          4349 => x"98",
          4350 => x"2e",
          4351 => x"75",
          4352 => x"05",
          4353 => x"98",
          4354 => x"98",
          4355 => x"98",
          4356 => x"07",
          4357 => x"53",
          4358 => x"26",
          4359 => x"08",
          4360 => x"98",
          4361 => x"58",
          4362 => x"08",
          4363 => x"38",
          4364 => x"5d",
          4365 => x"81",
          4366 => x"a9",
          4367 => x"ff",
          4368 => x"1b",
          4369 => x"39",
          4370 => x"82",
          4371 => x"30",
          4372 => x"5b",
          4373 => x"58",
          4374 => x"0c",
          4375 => x"33",
          4376 => x"34",
          4377 => x"0d",
          4378 => x"fc",
          4379 => x"3f",
          4380 => x"98",
          4381 => x"56",
          4382 => x"70",
          4383 => x"55",
          4384 => x"38",
          4385 => x"08",
          4386 => x"82",
          4387 => x"52",
          4388 => x"e0",
          4389 => x"80",
          4390 => x"51",
          4391 => x"08",
          4392 => x"81",
          4393 => x"09",
          4394 => x"39",
          4395 => x"98",
          4396 => x"98",
          4397 => x"52",
          4398 => x"e0",
          4399 => x"18",
          4400 => x"54",
          4401 => x"85",
          4402 => x"74",
          4403 => x"04",
          4404 => x"ff",
          4405 => x"cf",
          4406 => x"e0",
          4407 => x"a3",
          4408 => x"58",
          4409 => x"55",
          4410 => x"02",
          4411 => x"70",
          4412 => x"73",
          4413 => x"80",
          4414 => x"da",
          4415 => x"87",
          4416 => x"78",
          4417 => x"98",
          4418 => x"51",
          4419 => x"38",
          4420 => x"15",
          4421 => x"82",
          4422 => x"3d",
          4423 => x"82",
          4424 => x"08",
          4425 => x"52",
          4426 => x"e0",
          4427 => x"86",
          4428 => x"e0",
          4429 => x"e0",
          4430 => x"c7",
          4431 => x"e0",
          4432 => x"08",
          4433 => x"80",
          4434 => x"38",
          4435 => x"af",
          4436 => x"74",
          4437 => x"3f",
          4438 => x"e0",
          4439 => x"3d",
          4440 => x"05",
          4441 => x"82",
          4442 => x"08",
          4443 => x"8e",
          4444 => x"82",
          4445 => x"08",
          4446 => x"82",
          4447 => x"06",
          4448 => x"33",
          4449 => x"86",
          4450 => x"74",
          4451 => x"af",
          4452 => x"55",
          4453 => x"87",
          4454 => x"09",
          4455 => x"e0",
          4456 => x"86",
          4457 => x"81",
          4458 => x"78",
          4459 => x"98",
          4460 => x"9f",
          4461 => x"51",
          4462 => x"0b",
          4463 => x"80",
          4464 => x"52",
          4465 => x"3f",
          4466 => x"ff",
          4467 => x"11",
          4468 => x"ee",
          4469 => x"15",
          4470 => x"53",
          4471 => x"81",
          4472 => x"bf",
          4473 => x"82",
          4474 => x"b2",
          4475 => x"a3",
          4476 => x"51",
          4477 => x"0b",
          4478 => x"83",
          4479 => x"3f",
          4480 => x"80",
          4481 => x"a1",
          4482 => x"3d",
          4483 => x"84",
          4484 => x"aa",
          4485 => x"51",
          4486 => x"55",
          4487 => x"78",
          4488 => x"70",
          4489 => x"98",
          4490 => x"be",
          4491 => x"a0",
          4492 => x"38",
          4493 => x"3d",
          4494 => x"3f",
          4495 => x"52",
          4496 => x"08",
          4497 => x"e0",
          4498 => x"97",
          4499 => x"81",
          4500 => x"2e",
          4501 => x"82",
          4502 => x"06",
          4503 => x"92",
          4504 => x"e0",
          4505 => x"93",
          4506 => x"8d",
          4507 => x"af",
          4508 => x"33",
          4509 => x"55",
          4510 => x"54",
          4511 => x"0b",
          4512 => x"84",
          4513 => x"73",
          4514 => x"2e",
          4515 => x"ff",
          4516 => x"52",
          4517 => x"55",
          4518 => x"de",
          4519 => x"51",
          4520 => x"08",
          4521 => x"82",
          4522 => x"16",
          4523 => x"06",
          4524 => x"51",
          4525 => x"0b",
          4526 => x"98",
          4527 => x"3f",
          4528 => x"98",
          4529 => x"98",
          4530 => x"82",
          4531 => x"ec",
          4532 => x"02",
          4533 => x"57",
          4534 => x"97",
          4535 => x"98",
          4536 => x"cf",
          4537 => x"d0",
          4538 => x"98",
          4539 => x"38",
          4540 => x"06",
          4541 => x"a7",
          4542 => x"71",
          4543 => x"55",
          4544 => x"81",
          4545 => x"a2",
          4546 => x"74",
          4547 => x"04",
          4548 => x"94",
          4549 => x"d0",
          4550 => x"82",
          4551 => x"58",
          4552 => x"c4",
          4553 => x"82",
          4554 => x"c7",
          4555 => x"55",
          4556 => x"17",
          4557 => x"96",
          4558 => x"54",
          4559 => x"ff",
          4560 => x"55",
          4561 => x"0d",
          4562 => x"5a",
          4563 => x"9a",
          4564 => x"98",
          4565 => x"82",
          4566 => x"55",
          4567 => x"81",
          4568 => x"2e",
          4569 => x"80",
          4570 => x"ac",
          4571 => x"82",
          4572 => x"52",
          4573 => x"e0",
          4574 => x"bf",
          4575 => x"98",
          4576 => x"81",
          4577 => x"33",
          4578 => x"27",
          4579 => x"80",
          4580 => x"ff",
          4581 => x"56",
          4582 => x"76",
          4583 => x"80",
          4584 => x"78",
          4585 => x"2e",
          4586 => x"38",
          4587 => x"9f",
          4588 => x"82",
          4589 => x"33",
          4590 => x"2e",
          4591 => x"2e",
          4592 => x"05",
          4593 => x"98",
          4594 => x"0c",
          4595 => x"82",
          4596 => x"9d",
          4597 => x"98",
          4598 => x"82",
          4599 => x"53",
          4600 => x"ff",
          4601 => x"51",
          4602 => x"38",
          4603 => x"cc",
          4604 => x"ff",
          4605 => x"08",
          4606 => x"82",
          4607 => x"82",
          4608 => x"55",
          4609 => x"82",
          4610 => x"82",
          4611 => x"75",
          4612 => x"38",
          4613 => x"86",
          4614 => x"27",
          4615 => x"77",
          4616 => x"56",
          4617 => x"81",
          4618 => x"73",
          4619 => x"33",
          4620 => x"81",
          4621 => x"02",
          4622 => x"51",
          4623 => x"87",
          4624 => x"78",
          4625 => x"70",
          4626 => x"e0",
          4627 => x"80",
          4628 => x"ae",
          4629 => x"82",
          4630 => x"c4",
          4631 => x"c6",
          4632 => x"09",
          4633 => x"75",
          4634 => x"74",
          4635 => x"98",
          4636 => x"38",
          4637 => x"66",
          4638 => x"88",
          4639 => x"52",
          4640 => x"54",
          4641 => x"ff",
          4642 => x"54",
          4643 => x"9c",
          4644 => x"62",
          4645 => x"93",
          4646 => x"5e",
          4647 => x"08",
          4648 => x"38",
          4649 => x"38",
          4650 => x"08",
          4651 => x"70",
          4652 => x"55",
          4653 => x"39",
          4654 => x"82",
          4655 => x"89",
          4656 => x"56",
          4657 => x"06",
          4658 => x"82",
          4659 => x"7c",
          4660 => x"27",
          4661 => x"83",
          4662 => x"80",
          4663 => x"c1",
          4664 => x"14",
          4665 => x"82",
          4666 => x"38",
          4667 => x"95",
          4668 => x"81",
          4669 => x"06",
          4670 => x"56",
          4671 => x"b9",
          4672 => x"80",
          4673 => x"7a",
          4674 => x"73",
          4675 => x"ff",
          4676 => x"ff",
          4677 => x"58",
          4678 => x"74",
          4679 => x"73",
          4680 => x"7e",
          4681 => x"2e",
          4682 => x"8c",
          4683 => x"07",
          4684 => x"08",
          4685 => x"75",
          4686 => x"94",
          4687 => x"54",
          4688 => x"82",
          4689 => x"e8",
          4690 => x"80",
          4691 => x"5c",
          4692 => x"0b",
          4693 => x"38",
          4694 => x"f7",
          4695 => x"80",
          4696 => x"e0",
          4697 => x"82",
          4698 => x"12",
          4699 => x"51",
          4700 => x"08",
          4701 => x"57",
          4702 => x"82",
          4703 => x"56",
          4704 => x"05",
          4705 => x"cc",
          4706 => x"68",
          4707 => x"82",
          4708 => x"75",
          4709 => x"81",
          4710 => x"80",
          4711 => x"0a",
          4712 => x"55",
          4713 => x"8b",
          4714 => x"2a",
          4715 => x"59",
          4716 => x"70",
          4717 => x"56",
          4718 => x"80",
          4719 => x"52",
          4720 => x"56",
          4721 => x"83",
          4722 => x"82",
          4723 => x"55",
          4724 => x"09",
          4725 => x"29",
          4726 => x"74",
          4727 => x"17",
          4728 => x"98",
          4729 => x"92",
          4730 => x"b7",
          4731 => x"52",
          4732 => x"56",
          4733 => x"62",
          4734 => x"98",
          4735 => x"bf",
          4736 => x"26",
          4737 => x"8e",
          4738 => x"38",
          4739 => x"af",
          4740 => x"56",
          4741 => x"87",
          4742 => x"38",
          4743 => x"83",
          4744 => x"56",
          4745 => x"38",
          4746 => x"06",
          4747 => x"91",
          4748 => x"22",
          4749 => x"74",
          4750 => x"56",
          4751 => x"57",
          4752 => x"75",
          4753 => x"fe",
          4754 => x"84",
          4755 => x"5e",
          4756 => x"98",
          4757 => x"fd",
          4758 => x"38",
          4759 => x"8c",
          4760 => x"22",
          4761 => x"74",
          4762 => x"56",
          4763 => x"57",
          4764 => x"75",
          4765 => x"fe",
          4766 => x"10",
          4767 => x"9f",
          4768 => x"e0",
          4769 => x"05",
          4770 => x"56",
          4771 => x"81",
          4772 => x"67",
          4773 => x"30",
          4774 => x"59",
          4775 => x"81",
          4776 => x"42",
          4777 => x"90",
          4778 => x"51",
          4779 => x"75",
          4780 => x"67",
          4781 => x"82",
          4782 => x"09",
          4783 => x"08",
          4784 => x"78",
          4785 => x"78",
          4786 => x"82",
          4787 => x"83",
          4788 => x"27",
          4789 => x"55",
          4790 => x"59",
          4791 => x"74",
          4792 => x"88",
          4793 => x"26",
          4794 => x"1a",
          4795 => x"38",
          4796 => x"2e",
          4797 => x"9f",
          4798 => x"06",
          4799 => x"84",
          4800 => x"8f",
          4801 => x"52",
          4802 => x"80",
          4803 => x"3f",
          4804 => x"ff",
          4805 => x"99",
          4806 => x"83",
          4807 => x"80",
          4808 => x"ff",
          4809 => x"ff",
          4810 => x"ff",
          4811 => x"e9",
          4812 => x"51",
          4813 => x"1c",
          4814 => x"8d",
          4815 => x"51",
          4816 => x"1b",
          4817 => x"2e",
          4818 => x"88",
          4819 => x"ff",
          4820 => x"51",
          4821 => x"1b",
          4822 => x"b0",
          4823 => x"52",
          4824 => x"ff",
          4825 => x"0b",
          4826 => x"d1",
          4827 => x"39",
          4828 => x"51",
          4829 => x"ff",
          4830 => x"d1",
          4831 => x"a9",
          4832 => x"d2",
          4833 => x"86",
          4834 => x"1b",
          4835 => x"81",
          4836 => x"ff",
          4837 => x"98",
          4838 => x"09",
          4839 => x"86",
          4840 => x"88",
          4841 => x"7a",
          4842 => x"85",
          4843 => x"87",
          4844 => x"83",
          4845 => x"ff",
          4846 => x"8b",
          4847 => x"51",
          4848 => x"52",
          4849 => x"54",
          4850 => x"ff",
          4851 => x"53",
          4852 => x"3f",
          4853 => x"8c",
          4854 => x"83",
          4855 => x"52",
          4856 => x"52",
          4857 => x"f0",
          4858 => x"87",
          4859 => x"83",
          4860 => x"ff",
          4861 => x"74",
          4862 => x"54",
          4863 => x"86",
          4864 => x"be",
          4865 => x"08",
          4866 => x"76",
          4867 => x"cd",
          4868 => x"ff",
          4869 => x"83",
          4870 => x"26",
          4871 => x"53",
          4872 => x"3f",
          4873 => x"76",
          4874 => x"db",
          4875 => x"38",
          4876 => x"8a",
          4877 => x"38",
          4878 => x"81",
          4879 => x"ff",
          4880 => x"98",
          4881 => x"1b",
          4882 => x"54",
          4883 => x"7f",
          4884 => x"39",
          4885 => x"80",
          4886 => x"7a",
          4887 => x"d5",
          4888 => x"83",
          4889 => x"0b",
          4890 => x"34",
          4891 => x"34",
          4892 => x"75",
          4893 => x"85",
          4894 => x"2a",
          4895 => x"82",
          4896 => x"52",
          4897 => x"3f",
          4898 => x"88",
          4899 => x"52",
          4900 => x"56",
          4901 => x"53",
          4902 => x"3f",
          4903 => x"38",
          4904 => x"56",
          4905 => x"75",
          4906 => x"04",
          4907 => x"80",
          4908 => x"76",
          4909 => x"11",
          4910 => x"79",
          4911 => x"09",
          4912 => x"55",
          4913 => x"70",
          4914 => x"74",
          4915 => x"80",
          4916 => x"76",
          4917 => x"3d",
          4918 => x"84",
          4919 => x"8a",
          4920 => x"52",
          4921 => x"56",
          4922 => x"08",
          4923 => x"75",
          4924 => x"a1",
          4925 => x"53",
          4926 => x"97",
          4927 => x"72",
          4928 => x"56",
          4929 => x"88",
          4930 => x"3d",
          4931 => x"80",
          4932 => x"05",
          4933 => x"08",
          4934 => x"08",
          4935 => x"09",
          4936 => x"55",
          4937 => x"98",
          4938 => x"0d",
          4939 => x"73",
          4940 => x"0c",
          4941 => x"02",
          4942 => x"3d",
          4943 => x"52",
          4944 => x"ff",
          4945 => x"3d",
          4946 => x"22",
          4947 => x"26",
          4948 => x"52",
          4949 => x"27",
          4950 => x"06",
          4951 => x"82",
          4952 => x"9c",
          4953 => x"06",
          4954 => x"38",
          4955 => x"22",
          4956 => x"70",
          4957 => x"e0",
          4958 => x"3d",
          4959 => x"05",
          4960 => x"70",
          4961 => x"9a",
          4962 => x"06",
          4963 => x"38",
          4964 => x"22",
          4965 => x"84",
          4966 => x"51",
          4967 => x"38",
          4968 => x"ec",
          4969 => x"38",
          4970 => x"05",
          4971 => x"72",
          4972 => x"80",
          4973 => x"22",
          4974 => x"70",
          4975 => x"25",
          4976 => x"dc",
          4977 => x"05",
          4978 => x"10",
          4979 => x"80",
          4980 => x"72",
          4981 => x"12",
          4982 => x"39",
          4983 => x"51",
          4984 => x"ff",
          4985 => x"12",
          4986 => x"8c",
          4987 => x"16",
          4988 => x"82",
          4989 => x"00",
          4990 => x"ff",
          4991 => x"00",
          4992 => x"00",
          4993 => x"00",
          4994 => x"00",
          4995 => x"00",
          4996 => x"00",
          4997 => x"00",
          4998 => x"00",
          4999 => x"00",
          5000 => x"00",
          5001 => x"00",
          5002 => x"00",
          5003 => x"00",
          5004 => x"00",
          5005 => x"00",
          5006 => x"00",
          5007 => x"00",
          5008 => x"00",
          5009 => x"00",
          5010 => x"00",
          5011 => x"00",
          5012 => x"00",
          5013 => x"00",
          5014 => x"00",
          5015 => x"00",
          5016 => x"00",
          5017 => x"00",
          5018 => x"00",
          5019 => x"00",
          5020 => x"00",
          5021 => x"00",
          5022 => x"00",
          5023 => x"00",
          5024 => x"00",
          5025 => x"00",
          5026 => x"00",
          5027 => x"00",
          5028 => x"00",
          5029 => x"00",
          5030 => x"00",
          5031 => x"00",
          5032 => x"00",
          5033 => x"00",
          5034 => x"00",
          5035 => x"00",
          5036 => x"00",
          5037 => x"00",
          5038 => x"00",
          5039 => x"00",
          5040 => x"00",
          5041 => x"00",
          5042 => x"00",
          5043 => x"00",
          5044 => x"00",
          5045 => x"00",
          5046 => x"00",
          5047 => x"00",
          5048 => x"00",
          5049 => x"00",
          5050 => x"00",
          5051 => x"00",
          5052 => x"00",
          5053 => x"00",
          5054 => x"00",
          5055 => x"00",
          5056 => x"00",
          5057 => x"00",
          5058 => x"00",
          5059 => x"00",
          5060 => x"00",
          5061 => x"00",
          5062 => x"00",
          5063 => x"00",
          5064 => x"74",
          5065 => x"74",
          5066 => x"74",
          5067 => x"64",
          5068 => x"63",
          5069 => x"61",
          5070 => x"79",
          5071 => x"66",
          5072 => x"70",
          5073 => x"6d",
          5074 => x"68",
          5075 => x"68",
          5076 => x"63",
          5077 => x"6a",
          5078 => x"61",
          5079 => x"74",
          5080 => x"00",
          5081 => x"69",
          5082 => x"69",
          5083 => x"00",
          5084 => x"44",
          5085 => x"6f",
          5086 => x"72",
          5087 => x"6f",
          5088 => x"20",
          5089 => x"64",
          5090 => x"69",
          5091 => x"64",
          5092 => x"61",
          5093 => x"64",
          5094 => x"6c",
          5095 => x"6e",
          5096 => x"41",
          5097 => x"65",
          5098 => x"46",
          5099 => x"65",
          5100 => x"73",
          5101 => x"46",
          5102 => x"64",
          5103 => x"6c",
          5104 => x"53",
          5105 => x"69",
          5106 => x"65",
          5107 => x"44",
          5108 => x"6d",
          5109 => x"69",
          5110 => x"00",
          5111 => x"20",
          5112 => x"62",
          5113 => x"4e",
          5114 => x"74",
          5115 => x"6c",
          5116 => x"20",
          5117 => x"6e",
          5118 => x"46",
          5119 => x"62",
          5120 => x"54",
          5121 => x"20",
          5122 => x"6f",
          5123 => x"6c",
          5124 => x"46",
          5125 => x"6c",
          5126 => x"49",
          5127 => x"69",
          5128 => x"6f",
          5129 => x"54",
          5130 => x"20",
          5131 => x"6c",
          5132 => x"50",
          5133 => x"72",
          5134 => x"72",
          5135 => x"53",
          5136 => x"00",
          5137 => x"6f",
          5138 => x"72",
          5139 => x"20",
          5140 => x"73",
          5141 => x"20",
          5142 => x"65",
          5143 => x"72",
          5144 => x"25",
          5145 => x"3a",
          5146 => x"00",
          5147 => x"20",
          5148 => x"25",
          5149 => x"20",
          5150 => x"7c",
          5151 => x"2a",
          5152 => x"31",
          5153 => x"32",
          5154 => x"63",
          5155 => x"2c",
          5156 => x"32",
          5157 => x"73",
          5158 => x"5a",
          5159 => x"72",
          5160 => x"6e",
          5161 => x"54",
          5162 => x"74",
          5163 => x"50",
          5164 => x"72",
          5165 => x"49",
          5166 => x"20",
          5167 => x"70",
          5168 => x"4c",
          5169 => x"65",
          5170 => x"55",
          5171 => x"20",
          5172 => x"70",
          5173 => x"30",
          5174 => x"65",
          5175 => x"55",
          5176 => x"20",
          5177 => x"70",
          5178 => x"31",
          5179 => x"65",
          5180 => x"53",
          5181 => x"75",
          5182 => x"2e",
          5183 => x"6c",
          5184 => x"65",
          5185 => x"61",
          5186 => x"2e",
          5187 => x"7a",
          5188 => x"68",
          5189 => x"46",
          5190 => x"6f",
          5191 => x"6c",
          5192 => x"63",
          5193 => x"70",
          5194 => x"6e",
          5195 => x"61",
          5196 => x"2a",
          5197 => x"72",
          5198 => x"00",
          5199 => x"69",
          5200 => x"43",
          5201 => x"67",
          5202 => x"25",
          5203 => x"38",
          5204 => x"6c",
          5205 => x"0a",
          5206 => x"20",
          5207 => x"0a",
          5208 => x"65",
          5209 => x"58",
          5210 => x"3f",
          5211 => x"58",
          5212 => x"25",
          5213 => x"38",
          5214 => x"45",
          5215 => x"67",
          5216 => x"20",
          5217 => x"2e",
          5218 => x"69",
          5219 => x"20",
          5220 => x"20",
          5221 => x"43",
          5222 => x"75",
          5223 => x"64",
          5224 => x"0a",
          5225 => x"61",
          5226 => x"70",
          5227 => x"6f",
          5228 => x"43",
          5229 => x"6f",
          5230 => x"2e",
          5231 => x"62",
          5232 => x"25",
          5233 => x"00",
          5234 => x"25",
          5235 => x"25",
          5236 => x"42",
          5237 => x"61",
          5238 => x"4d",
          5239 => x"78",
          5240 => x"2c",
          5241 => x"20",
          5242 => x"20",
          5243 => x"2e",
          5244 => x"69",
          5245 => x"45",
          5246 => x"20",
          5247 => x"70",
          5248 => x"25",
          5249 => x"20",
          5250 => x"64",
          5251 => x"53",
          5252 => x"69",
          5253 => x"6e",
          5254 => x"6f",
          5255 => x"6f",
          5256 => x"3a",
          5257 => x"73",
          5258 => x"65",
          5259 => x"20",
          5260 => x"44",
          5261 => x"30",
          5262 => x"29",
          5263 => x"53",
          5264 => x"20",
          5265 => x"25",
          5266 => x"20",
          5267 => x"20",
          5268 => x"30",
          5269 => x"29",
          5270 => x"42",
          5271 => x"20",
          5272 => x"25",
          5273 => x"20",
          5274 => x"20",
          5275 => x"30",
          5276 => x"29",
          5277 => x"53",
          5278 => x"20",
          5279 => x"65",
          5280 => x"29",
          5281 => x"54",
          5282 => x"20",
          5283 => x"73",
          5284 => x"29",
          5285 => x"49",
          5286 => x"4c",
          5287 => x"65",
          5288 => x"29",
          5289 => x"57",
          5290 => x"20",
          5291 => x"20",
          5292 => x"32",
          5293 => x"49",
          5294 => x"20",
          5295 => x"20",
          5296 => x"41",
          5297 => x"73",
          5298 => x"43",
          5299 => x"74",
          5300 => x"20",
          5301 => x"20",
          5302 => x"00",
          5303 => x"43",
          5304 => x"72",
          5305 => x"20",
          5306 => x"20",
          5307 => x"00",
          5308 => x"53",
          5309 => x"61",
          5310 => x"65",
          5311 => x"20",
          5312 => x"00",
          5313 => x"3a",
          5314 => x"5a",
          5315 => x"20",
          5316 => x"20",
          5317 => x"20",
          5318 => x"00",
          5319 => x"53",
          5320 => x"6c",
          5321 => x"71",
          5322 => x"20",
          5323 => x"34",
          5324 => x"20",
          5325 => x"4d",
          5326 => x"46",
          5327 => x"20",
          5328 => x"64",
          5329 => x"7a",
          5330 => x"57",
          5331 => x"20",
          5332 => x"6c",
          5333 => x"71",
          5334 => x"34",
          5335 => x"53",
          5336 => x"4d",
          5337 => x"46",
          5338 => x"45",
          5339 => x"00",
          5340 => x"6f",
          5341 => x"01",
          5342 => x"00",
          5343 => x"00",
          5344 => x"01",
          5345 => x"00",
          5346 => x"00",
          5347 => x"01",
          5348 => x"00",
          5349 => x"00",
          5350 => x"01",
          5351 => x"00",
          5352 => x"00",
          5353 => x"01",
          5354 => x"00",
          5355 => x"00",
          5356 => x"01",
          5357 => x"00",
          5358 => x"00",
          5359 => x"04",
          5360 => x"00",
          5361 => x"00",
          5362 => x"03",
          5363 => x"00",
          5364 => x"00",
          5365 => x"04",
          5366 => x"00",
          5367 => x"00",
          5368 => x"03",
          5369 => x"00",
          5370 => x"00",
          5371 => x"03",
          5372 => x"00",
          5373 => x"00",
          5374 => x"1b",
          5375 => x"1b",
          5376 => x"1b",
          5377 => x"1b",
          5378 => x"1b",
          5379 => x"10",
          5380 => x"0d",
          5381 => x"08",
          5382 => x"05",
          5383 => x"03",
          5384 => x"01",
          5385 => x"6f",
          5386 => x"00",
          5387 => x"25",
          5388 => x"73",
          5389 => x"65",
          5390 => x"73",
          5391 => x"68",
          5392 => x"66",
          5393 => x"45",
          5394 => x"43",
          5395 => x"70",
          5396 => x"74",
          5397 => x"72",
          5398 => x"20",
          5399 => x"6e",
          5400 => x"22",
          5401 => x"00",
          5402 => x"5b",
          5403 => x"46",
          5404 => x"eb",
          5405 => x"35",
          5406 => x"41",
          5407 => x"41",
          5408 => x"4e",
          5409 => x"20",
          5410 => x"20",
          5411 => x"00",
          5412 => x"00",
          5413 => x"09",
          5414 => x"1e",
          5415 => x"8e",
          5416 => x"49",
          5417 => x"99",
          5418 => x"9c",
          5419 => x"a5",
          5420 => x"ac",
          5421 => x"b4",
          5422 => x"bc",
          5423 => x"c4",
          5424 => x"cc",
          5425 => x"d4",
          5426 => x"dc",
          5427 => x"e4",
          5428 => x"ec",
          5429 => x"f4",
          5430 => x"fc",
          5431 => x"3d",
          5432 => x"3c",
          5433 => x"00",
          5434 => x"01",
          5435 => x"00",
          5436 => x"00",
          5437 => x"00",
          5438 => x"00",
          5439 => x"00",
          5440 => x"00",
          5441 => x"00",
          5442 => x"00",
          5443 => x"00",
          5444 => x"00",
          5445 => x"00",
          5446 => x"00",
          5447 => x"00",
          5448 => x"00",
          5449 => x"25",
          5450 => x"25",
          5451 => x"25",
          5452 => x"25",
          5453 => x"25",
          5454 => x"25",
          5455 => x"25",
          5456 => x"25",
          5457 => x"25",
          5458 => x"25",
          5459 => x"25",
          5460 => x"25",
          5461 => x"03",
          5462 => x"03",
          5463 => x"03",
          5464 => x"22",
          5465 => x"22",
          5466 => x"23",
          5467 => x"00",
          5468 => x"20",
          5469 => x"00",
          5470 => x"00",
          5471 => x"01",
          5472 => x"01",
          5473 => x"01",
          5474 => x"00",
          5475 => x"01",
          5476 => x"01",
          5477 => x"01",
          5478 => x"01",
          5479 => x"01",
          5480 => x"01",
          5481 => x"01",
          5482 => x"01",
          5483 => x"01",
          5484 => x"01",
          5485 => x"01",
          5486 => x"01",
          5487 => x"01",
          5488 => x"01",
          5489 => x"01",
          5490 => x"01",
          5491 => x"01",
          5492 => x"01",
          5493 => x"01",
          5494 => x"01",
          5495 => x"01",
          5496 => x"01",
          5497 => x"02",
          5498 => x"2c",
          5499 => x"2c",
          5500 => x"02",
          5501 => x"00",
          5502 => x"01",
          5503 => x"02",
          5504 => x"02",
          5505 => x"02",
          5506 => x"02",
          5507 => x"02",
          5508 => x"02",
          5509 => x"01",
          5510 => x"02",
          5511 => x"02",
          5512 => x"02",
          5513 => x"02",
          5514 => x"02",
          5515 => x"01",
          5516 => x"02",
          5517 => x"01",
          5518 => x"03",
          5519 => x"03",
          5520 => x"03",
          5521 => x"03",
          5522 => x"03",
          5523 => x"03",
          5524 => x"00",
          5525 => x"03",
          5526 => x"03",
          5527 => x"03",
          5528 => x"01",
          5529 => x"01",
          5530 => x"04",
          5531 => x"00",
          5532 => x"2c",
          5533 => x"01",
          5534 => x"06",
          5535 => x"06",
          5536 => x"00",
          5537 => x"1f",
          5538 => x"1f",
          5539 => x"1f",
          5540 => x"1f",
          5541 => x"1f",
          5542 => x"1f",
          5543 => x"1f",
          5544 => x"1f",
          5545 => x"1f",
          5546 => x"1f",
          5547 => x"06",
          5548 => x"1f",
          5549 => x"00",
          5550 => x"21",
          5551 => x"05",
          5552 => x"01",
          5553 => x"01",
          5554 => x"08",
          5555 => x"00",
          5556 => x"01",
          5557 => x"00",
          5558 => x"01",
          5559 => x"00",
          5560 => x"01",
          5561 => x"00",
          5562 => x"01",
          5563 => x"00",
          5564 => x"01",
          5565 => x"00",
          5566 => x"01",
          5567 => x"00",
          5568 => x"01",
          5569 => x"00",
          5570 => x"01",
          5571 => x"00",
          5572 => x"01",
          5573 => x"00",
          5574 => x"01",
          5575 => x"00",
          5576 => x"01",
          5577 => x"00",
          5578 => x"01",
          5579 => x"00",
          5580 => x"01",
          5581 => x"00",
          5582 => x"01",
          5583 => x"00",
          5584 => x"01",
          5585 => x"00",
          5586 => x"01",
          5587 => x"00",
          5588 => x"01",
          5589 => x"00",
          5590 => x"01",
          5591 => x"00",
          5592 => x"01",
          5593 => x"00",
          5594 => x"01",
          5595 => x"00",
          5596 => x"01",
          5597 => x"00",
          5598 => x"01",
          5599 => x"00",
          5600 => x"01",
          5601 => x"00",
          5602 => x"01",
          5603 => x"00",
          5604 => x"01",
          5605 => x"00",
          5606 => x"00",
          5607 => x"00",
          5608 => x"00",
          5609 => x"00",
          5610 => x"01",
          5611 => x"00",
          5612 => x"00",
          5613 => x"05",
          5614 => x"05",
          5615 => x"01",
          5616 => x"01",
          5617 => x"00",
          5618 => x"00",
          5619 => x"00",
          5620 => x"00",
          5621 => x"00",
          5622 => x"00",
          5623 => x"00",
          5624 => x"00",
          5625 => x"00",
          5626 => x"00",
          5627 => x"00",
          5628 => x"00",
          5629 => x"00",
          5630 => x"00",
          5631 => x"00",
          5632 => x"00",
          5633 => x"00",
          5634 => x"01",
        others => X"00"
    );

    signal RAM0_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM1_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM2_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM3_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM4_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM5_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM6_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM7_DATA         :     std_logic_vector(7 downto 0);         -- Buffer for byte in word to be written.
    signal RAM0_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM1_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM2_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM3_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM4_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM5_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM6_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal RAM7_WREN         :     std_logic;                            -- Write Enable for this particular byte in word.
    signal lowDataA          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataA         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.
    signal lowDataB          :     std_logic_vector(WORD_32BIT_RANGE);   -- Low word in 64 bit output from RAM matrix.
    signal highDataB         :     std_logic_vector(WORD_32BIT_RANGE);   -- High word in 64 bit output from RAM matrix.

begin

    -- Correctly assign the Little Endian value to the correct array, byte writes the data is in '7 downto 0', h-word writes
    -- the data is in '15 downto 0', word writes the data is in '31 downto 0'. Long words (64bits) are treated as two words for Endianness,
    -- and not as one continuous long word, this is because the ZPU is 32bit even when accessing a 64bit chunk.
    --
    RAM0_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '0'
                 else (others => '0');
    RAM1_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '0' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '0' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM4_DATA <= memAWrite(7 downto 0)   when memAAddr(2) = '1'
                 else (others => '0');
    RAM5_DATA <= memAWrite(15 downto 8)  when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);
    RAM6_DATA <= memAWrite(23 downto 16) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(7 downto 0);
    RAM7_DATA <= memAWrite(31 downto 24) when memAAddr(2) = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0'))
                 else
                 memAWrite(15 downto 8)  when memAAddr(2) = '1' and (memAWriteHalfWord = '1')
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "011") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "010") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "01"))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "001") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '0') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "000") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "00"))
                 else '0';
    RAM4_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "111") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM5_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "110") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "11"))
                 else '0';
    RAM6_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "101") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';
    RAM7_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0' and memAAddr(2) = '1') or (memAWriteByte = '1' and memAAddr(2 downto 0) = "100") or (memAWriteHalfWord = '1' and memAAddr(2 downto 1) = "10"))
                 else '0';

    memARead  <= lowDataA  when memAAddr(2) = '0'
                 else
                 highDataA;
    memBRead  <= lowDataB & highDataB;

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM0_DATA;
            else
                lowDataA(7 downto 0)    <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM1_DATA;
            else
                lowDataA(15 downto 8)   <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM2_DATA;
            else
                lowDataA(23 downto 16)  <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM3_DATA;
            else
                lowDataA(31 downto 24)  <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 4 - Port A - bits 39 to 32 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM4_WREN = '1' then
                RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM4_DATA;
            else
                highDataA(7 downto 0)   <= RAM4(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 5 - Port A - bits 47 to 40 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM5_WREN = '1' then
                RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM5_DATA;
            else
                highDataA(15 downto 8)  <= RAM5(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 6 - Port A - bits 56 to 48
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM6_WREN = '1' then
                RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM6_DATA;
            else
                highDataA(23 downto 16) <= RAM6(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- RAM Byte 7 - Port A - bits 63 to 57 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM7_WREN = '1' then
                RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3)))) := RAM7_DATA;
            else
                highDataA(31 downto 24) <= RAM7(to_integer(unsigned(memAAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;


    -- BRAM Byte 0 - Port B - bits 7 downto 0
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(7 downto 0);
                lowDataB(7 downto 0)    <= memBWrite(7 downto 0);
            else
                lowDataB(7 downto 0)    <= RAM0(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 1 - Port B - bits 15 downto 8
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(15 downto 8);
                lowDataB(15 downto 8)    <= memBWrite(15 downto 8);
            else
                lowDataB(15 downto 8)    <= RAM1(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 2 - Port B - bits 23 downto 16
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(23 downto 16);
                lowDataB(23 downto 16)  <= memBWrite(23 downto 16);
            else
                lowDataB(23 downto 16)  <= RAM2(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 3 - Port B - bits 31 downto 24
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(31 downto 24);
                lowDataB(31 downto 24)  <= memBWrite(31 downto 24);
            else
                lowDataB(31 downto 24)  <= RAM3(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 4 - Port B - bits 39 downto 32
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(39 downto 32);
                highDataB(7 downto 0)   <= memBWrite(39 downto 32);
            else
                highDataB(7 downto 0)   <= RAM4(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 5 - Port B - bits 47 downto 40
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(47 downto 40);
                highDataB(15 downto 8)  <= memBWrite(47 downto 40);
            else
                highDataB(15 downto 8)  <= RAM5(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 6 - Port B - bits 55 downto 48
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(55 downto 48);
                highDataB(23 downto 16)  <= memBWrite(55 downto 48);
            else
                highDataB(23 downto 16)  <= RAM6(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

    -- BRAM Byte 7 - Port B - bits 63 downto 56 
    process(clk)
    begin
        if rising_edge(clk) then
            if memBWriteEnable = '1' then
                RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3)))) := memBWrite(63 downto 56);
                highDataB(31 downto 24)  <= memBWrite(63 downto 56);
            else
                highDataB(31 downto 24)  <= RAM7(to_integer(unsigned(memBAddr(addrbits-1 downto 3))));
            end if;
        end if;
    end process;

end arch;
