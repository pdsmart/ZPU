-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBootBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBootBRAM;

architecture arch of SinglePortBootBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"88",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"0b",
            10 => x"08",
            11 => x"8c",
            12 => x"04",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"08",
            17 => x"09",
            18 => x"05",
            19 => x"83",
            20 => x"52",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"08",
            25 => x"73",
            26 => x"81",
            27 => x"83",
            28 => x"06",
            29 => x"ff",
            30 => x"0b",
            31 => x"00",
            32 => x"05",
            33 => x"73",
            34 => x"06",
            35 => x"06",
            36 => x"06",
            37 => x"00",
            38 => x"00",
            39 => x"00",
            40 => x"73",
            41 => x"53",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"09",
            49 => x"06",
            50 => x"72",
            51 => x"72",
            52 => x"31",
            53 => x"06",
            54 => x"51",
            55 => x"00",
            56 => x"73",
            57 => x"53",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"88",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"2b",
            81 => x"04",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"06",
            89 => x"0b",
            90 => x"a7",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"ff",
            97 => x"2a",
            98 => x"0a",
            99 => x"05",
           100 => x"51",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"51",
           105 => x"83",
           106 => x"05",
           107 => x"2b",
           108 => x"72",
           109 => x"51",
           110 => x"00",
           111 => x"00",
           112 => x"05",
           113 => x"70",
           114 => x"06",
           115 => x"53",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"05",
           121 => x"70",
           122 => x"06",
           123 => x"06",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"05",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"81",
           137 => x"51",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"06",
           145 => x"06",
           146 => x"04",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"08",
           153 => x"09",
           154 => x"05",
           155 => x"2a",
           156 => x"52",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"08",
           161 => x"9f",
           162 => x"06",
           163 => x"08",
           164 => x"0b",
           165 => x"00",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"75",
           170 => x"89",
           171 => x"50",
           172 => x"90",
           173 => x"88",
           174 => x"00",
           175 => x"00",
           176 => x"08",
           177 => x"75",
           178 => x"8b",
           179 => x"50",
           180 => x"90",
           181 => x"88",
           182 => x"00",
           183 => x"00",
           184 => x"81",
           185 => x"0a",
           186 => x"05",
           187 => x"06",
           188 => x"74",
           189 => x"06",
           190 => x"51",
           191 => x"00",
           192 => x"81",
           193 => x"0a",
           194 => x"ff",
           195 => x"71",
           196 => x"72",
           197 => x"05",
           198 => x"51",
           199 => x"00",
           200 => x"04",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"52",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"72",
           233 => x"52",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"ff",
           249 => x"51",
           250 => x"00",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"53",
           266 => x"00",
           267 => x"06",
           268 => x"09",
           269 => x"05",
           270 => x"2b",
           271 => x"06",
           272 => x"04",
           273 => x"72",
           274 => x"05",
           275 => x"05",
           276 => x"72",
           277 => x"53",
           278 => x"51",
           279 => x"04",
           280 => x"a0",
           281 => x"38",
           282 => x"84",
           283 => x"0b",
           284 => x"e2",
           285 => x"51",
           286 => x"00",
           287 => x"88",
           288 => x"00",
           289 => x"02",
           290 => x"3d",
           291 => x"94",
           292 => x"08",
           293 => x"88",
           294 => x"82",
           295 => x"08",
           296 => x"54",
           297 => x"94",
           298 => x"08",
           299 => x"fd",
           300 => x"53",
           301 => x"05",
           302 => x"08",
           303 => x"51",
           304 => x"88",
           305 => x"0c",
           306 => x"0d",
           307 => x"94",
           308 => x"0c",
           309 => x"80",
           310 => x"fc",
           311 => x"08",
           312 => x"80",
           313 => x"94",
           314 => x"08",
           315 => x"88",
           316 => x"0b",
           317 => x"05",
           318 => x"fc",
           319 => x"38",
           320 => x"08",
           321 => x"94",
           322 => x"08",
           323 => x"05",
           324 => x"8c",
           325 => x"25",
           326 => x"08",
           327 => x"30",
           328 => x"05",
           329 => x"94",
           330 => x"0c",
           331 => x"05",
           332 => x"81",
           333 => x"f0",
           334 => x"08",
           335 => x"94",
           336 => x"0c",
           337 => x"08",
           338 => x"52",
           339 => x"05",
           340 => x"a7",
           341 => x"70",
           342 => x"05",
           343 => x"08",
           344 => x"80",
           345 => x"94",
           346 => x"08",
           347 => x"f8",
           348 => x"08",
           349 => x"70",
           350 => x"89",
           351 => x"0c",
           352 => x"02",
           353 => x"3d",
           354 => x"94",
           355 => x"0c",
           356 => x"05",
           357 => x"93",
           358 => x"88",
           359 => x"94",
           360 => x"0c",
           361 => x"08",
           362 => x"94",
           363 => x"08",
           364 => x"38",
           365 => x"05",
           366 => x"08",
           367 => x"81",
           368 => x"8c",
           369 => x"94",
           370 => x"08",
           371 => x"88",
           372 => x"08",
           373 => x"54",
           374 => x"05",
           375 => x"8c",
           376 => x"f8",
           377 => x"94",
           378 => x"0c",
           379 => x"05",
           380 => x"0c",
           381 => x"0d",
           382 => x"94",
           383 => x"0c",
           384 => x"81",
           385 => x"fc",
           386 => x"0b",
           387 => x"05",
           388 => x"8c",
           389 => x"08",
           390 => x"27",
           391 => x"08",
           392 => x"80",
           393 => x"80",
           394 => x"8c",
           395 => x"99",
           396 => x"8c",
           397 => x"94",
           398 => x"0c",
           399 => x"05",
           400 => x"08",
           401 => x"c9",
           402 => x"fc",
           403 => x"2e",
           404 => x"94",
           405 => x"08",
           406 => x"05",
           407 => x"38",
           408 => x"05",
           409 => x"8c",
           410 => x"94",
           411 => x"0c",
           412 => x"05",
           413 => x"fc",
           414 => x"94",
           415 => x"0c",
           416 => x"05",
           417 => x"94",
           418 => x"0c",
           419 => x"05",
           420 => x"94",
           421 => x"0c",
           422 => x"94",
           423 => x"08",
           424 => x"38",
           425 => x"05",
           426 => x"08",
           427 => x"51",
           428 => x"08",
           429 => x"70",
           430 => x"05",
           431 => x"08",
           432 => x"88",
           433 => x"0d",
           434 => x"ff",
           435 => x"88",
           436 => x"92",
           437 => x"0b",
           438 => x"8c",
           439 => x"87",
           440 => x"0c",
           441 => x"8c",
           442 => x"06",
           443 => x"80",
           444 => x"87",
           445 => x"08",
           446 => x"38",
           447 => x"8c",
           448 => x"80",
           449 => x"93",
           450 => x"98",
           451 => x"70",
           452 => x"38",
           453 => x"0b",
           454 => x"0b",
           455 => x"f0",
           456 => x"83",
           457 => x"fa",
           458 => x"7b",
           459 => x"56",
           460 => x"0b",
           461 => x"33",
           462 => x"55",
           463 => x"75",
           464 => x"06",
           465 => x"85",
           466 => x"98",
           467 => x"87",
           468 => x"0c",
           469 => x"c0",
           470 => x"87",
           471 => x"08",
           472 => x"70",
           473 => x"52",
           474 => x"2e",
           475 => x"c0",
           476 => x"70",
           477 => x"76",
           478 => x"53",
           479 => x"2e",
           480 => x"80",
           481 => x"71",
           482 => x"05",
           483 => x"14",
           484 => x"55",
           485 => x"51",
           486 => x"8b",
           487 => x"98",
           488 => x"70",
           489 => x"87",
           490 => x"08",
           491 => x"38",
           492 => x"c0",
           493 => x"87",
           494 => x"08",
           495 => x"51",
           496 => x"38",
           497 => x"80",
           498 => x"52",
           499 => x"09",
           500 => x"38",
           501 => x"8c",
           502 => x"72",
           503 => x"06",
           504 => x"52",
           505 => x"88",
           506 => x"fe",
           507 => x"81",
           508 => x"33",
           509 => x"07",
           510 => x"51",
           511 => x"04",
           512 => x"75",
           513 => x"82",
           514 => x"90",
           515 => x"2b",
           516 => x"33",
           517 => x"88",
           518 => x"71",
           519 => x"52",
           520 => x"54",
           521 => x"0d",
           522 => x"0d",
           523 => x"0b",
           524 => x"57",
           525 => x"27",
           526 => x"76",
           527 => x"27",
           528 => x"75",
           529 => x"82",
           530 => x"74",
           531 => x"38",
           532 => x"74",
           533 => x"83",
           534 => x"76",
           535 => x"17",
           536 => x"88",
           537 => x"55",
           538 => x"88",
           539 => x"74",
           540 => x"3f",
           541 => x"ff",
           542 => x"ad",
           543 => x"76",
           544 => x"fc",
           545 => x"87",
           546 => x"08",
           547 => x"3d",
           548 => x"fd",
           549 => x"08",
           550 => x"51",
           551 => x"88",
           552 => x"06",
           553 => x"81",
           554 => x"0c",
           555 => x"04",
           556 => x"0b",
           557 => x"f4",
           558 => x"88",
           559 => x"05",
           560 => x"80",
           561 => x"27",
           562 => x"14",
           563 => x"29",
           564 => x"05",
           565 => x"88",
           566 => x"0d",
           567 => x"0d",
           568 => x"0b",
           569 => x"9f",
           570 => x"33",
           571 => x"71",
           572 => x"81",
           573 => x"94",
           574 => x"ef",
           575 => x"90",
           576 => x"14",
           577 => x"3f",
           578 => x"ff",
           579 => x"07",
           580 => x"3d",
           581 => x"3d",
           582 => x"0b",
           583 => x"08",
           584 => x"75",
           585 => x"08",
           586 => x"2e",
           587 => x"14",
           588 => x"85",
           589 => x"b0",
           590 => x"38",
           591 => x"71",
           592 => x"81",
           593 => x"90",
           594 => x"72",
           595 => x"72",
           596 => x"38",
           597 => x"d8",
           598 => x"52",
           599 => x"14",
           600 => x"90",
           601 => x"52",
           602 => x"86",
           603 => x"fa",
           604 => x"0b",
           605 => x"f4",
           606 => x"81",
           607 => x"ff",
           608 => x"54",
           609 => x"80",
           610 => x"90",
           611 => x"72",
           612 => x"52",
           613 => x"73",
           614 => x"71",
           615 => x"81",
           616 => x"0c",
           617 => x"53",
           618 => x"83",
           619 => x"22",
           620 => x"76",
           621 => x"b5",
           622 => x"33",
           623 => x"84",
           624 => x"71",
           625 => x"51",
           626 => x"81",
           627 => x"08",
           628 => x"83",
           629 => x"88",
           630 => x"96",
           631 => x"8c",
           632 => x"08",
           633 => x"3f",
           634 => x"16",
           635 => x"23",
           636 => x"88",
           637 => x"0d",
           638 => x"0d",
           639 => x"58",
           640 => x"33",
           641 => x"2e",
           642 => x"88",
           643 => x"70",
           644 => x"39",
           645 => x"56",
           646 => x"2e",
           647 => x"84",
           648 => x"43",
           649 => x"1d",
           650 => x"33",
           651 => x"9f",
           652 => x"7b",
           653 => x"3f",
           654 => x"80",
           655 => x"d3",
           656 => x"84",
           657 => x"58",
           658 => x"55",
           659 => x"81",
           660 => x"ff",
           661 => x"ff",
           662 => x"06",
           663 => x"70",
           664 => x"7f",
           665 => x"7a",
           666 => x"81",
           667 => x"13",
           668 => x"af",
           669 => x"a0",
           670 => x"80",
           671 => x"51",
           672 => x"5d",
           673 => x"80",
           674 => x"ae",
           675 => x"06",
           676 => x"55",
           677 => x"75",
           678 => x"80",
           679 => x"79",
           680 => x"30",
           681 => x"70",
           682 => x"07",
           683 => x"51",
           684 => x"75",
           685 => x"58",
           686 => x"ab",
           687 => x"19",
           688 => x"06",
           689 => x"5a",
           690 => x"75",
           691 => x"39",
           692 => x"0c",
           693 => x"a0",
           694 => x"81",
           695 => x"1a",
           696 => x"fc",
           697 => x"08",
           698 => x"a0",
           699 => x"70",
           700 => x"e0",
           701 => x"90",
           702 => x"7c",
           703 => x"3f",
           704 => x"88",
           705 => x"38",
           706 => x"74",
           707 => x"ee",
           708 => x"33",
           709 => x"70",
           710 => x"56",
           711 => x"38",
           712 => x"1e",
           713 => x"59",
           714 => x"ff",
           715 => x"ff",
           716 => x"79",
           717 => x"5b",
           718 => x"81",
           719 => x"71",
           720 => x"56",
           721 => x"2e",
           722 => x"39",
           723 => x"92",
           724 => x"fc",
           725 => x"8e",
           726 => x"56",
           727 => x"38",
           728 => x"56",
           729 => x"8b",
           730 => x"55",
           731 => x"8b",
           732 => x"84",
           733 => x"06",
           734 => x"74",
           735 => x"56",
           736 => x"56",
           737 => x"51",
           738 => x"88",
           739 => x"0c",
           740 => x"75",
           741 => x"3d",
           742 => x"3d",
           743 => x"59",
           744 => x"83",
           745 => x"52",
           746 => x"fb",
           747 => x"88",
           748 => x"38",
           749 => x"b3",
           750 => x"83",
           751 => x"55",
           752 => x"82",
           753 => x"09",
           754 => x"ce",
           755 => x"b6",
           756 => x"76",
           757 => x"3f",
           758 => x"88",
           759 => x"76",
           760 => x"3f",
           761 => x"ff",
           762 => x"74",
           763 => x"2e",
           764 => x"54",
           765 => x"77",
           766 => x"f6",
           767 => x"08",
           768 => x"94",
           769 => x"f7",
           770 => x"08",
           771 => x"06",
           772 => x"82",
           773 => x"38",
           774 => x"88",
           775 => x"0d",
           776 => x"0d",
           777 => x"0b",
           778 => x"9f",
           779 => x"9b",
           780 => x"81",
           781 => x"56",
           782 => x"38",
           783 => x"8d",
           784 => x"57",
           785 => x"3f",
           786 => x"ff",
           787 => x"81",
           788 => x"06",
           789 => x"54",
           790 => x"74",
           791 => x"f5",
           792 => x"08",
           793 => x"3d",
           794 => x"80",
           795 => x"95",
           796 => x"51",
           797 => x"88",
           798 => x"53",
           799 => x"fe",
           800 => x"08",
           801 => x"57",
           802 => x"09",
           803 => x"38",
           804 => x"99",
           805 => x"2e",
           806 => x"56",
           807 => x"a4",
           808 => x"79",
           809 => x"f4",
           810 => x"56",
           811 => x"fd",
           812 => x"e5",
           813 => x"b3",
           814 => x"83",
           815 => x"58",
           816 => x"95",
           817 => x"51",
           818 => x"88",
           819 => x"af",
           820 => x"71",
           821 => x"05",
           822 => x"54",
           823 => x"f6",
           824 => x"08",
           825 => x"06",
           826 => x"1a",
           827 => x"33",
           828 => x"95",
           829 => x"51",
           830 => x"88",
           831 => x"23",
           832 => x"05",
           833 => x"3f",
           834 => x"ff",
           835 => x"75",
           836 => x"3d",
           837 => x"f5",
           838 => x"08",
           839 => x"f5",
           840 => x"08",
           841 => x"06",
           842 => x"79",
           843 => x"22",
           844 => x"82",
           845 => x"72",
           846 => x"59",
           847 => x"ee",
           848 => x"08",
           849 => x"88",
           850 => x"08",
           851 => x"56",
           852 => x"df",
           853 => x"38",
           854 => x"ff",
           855 => x"85",
           856 => x"89",
           857 => x"76",
           858 => x"c1",
           859 => x"34",
           860 => x"09",
           861 => x"38",
           862 => x"05",
           863 => x"3f",
           864 => x"1a",
           865 => x"8c",
           866 => x"90",
           867 => x"83",
           868 => x"8c",
           869 => x"71",
           870 => x"94",
           871 => x"80",
           872 => x"34",
           873 => x"0b",
           874 => x"80",
           875 => x"0c",
           876 => x"04",
           877 => x"0b",
           878 => x"f4",
           879 => x"54",
           880 => x"80",
           881 => x"0b",
           882 => x"98",
           883 => x"45",
           884 => x"3d",
           885 => x"ec",
           886 => x"9d",
           887 => x"54",
           888 => x"c0",
           889 => x"33",
           890 => x"2e",
           891 => x"a7",
           892 => x"84",
           893 => x"06",
           894 => x"73",
           895 => x"38",
           896 => x"39",
           897 => x"d5",
           898 => x"a0",
           899 => x"3d",
           900 => x"f3",
           901 => x"08",
           902 => x"73",
           903 => x"81",
           904 => x"34",
           905 => x"98",
           906 => x"f6",
           907 => x"7f",
           908 => x"0b",
           909 => x"59",
           910 => x"80",
           911 => x"57",
           912 => x"81",
           913 => x"16",
           914 => x"55",
           915 => x"80",
           916 => x"38",
           917 => x"81",
           918 => x"39",
           919 => x"17",
           920 => x"81",
           921 => x"16",
           922 => x"08",
           923 => x"78",
           924 => x"74",
           925 => x"2e",
           926 => x"98",
           927 => x"83",
           928 => x"57",
           929 => x"38",
           930 => x"ff",
           931 => x"2a",
           932 => x"ff",
           933 => x"79",
           934 => x"87",
           935 => x"08",
           936 => x"a4",
           937 => x"f3",
           938 => x"08",
           939 => x"27",
           940 => x"74",
           941 => x"a4",
           942 => x"f3",
           943 => x"08",
           944 => x"80",
           945 => x"38",
           946 => x"a8",
           947 => x"16",
           948 => x"06",
           949 => x"31",
           950 => x"75",
           951 => x"77",
           952 => x"98",
           953 => x"ff",
           954 => x"16",
           955 => x"51",
           956 => x"88",
           957 => x"38",
           958 => x"15",
           959 => x"77",
           960 => x"08",
           961 => x"58",
           962 => x"fe",
           963 => x"19",
           964 => x"39",
           965 => x"88",
           966 => x"0d",
           967 => x"0d",
           968 => x"8c",
           969 => x"84",
           970 => x"51",
           971 => x"88",
           972 => x"87",
           973 => x"08",
           974 => x"84",
           975 => x"51",
           976 => x"73",
           977 => x"87",
           978 => x"0c",
           979 => x"9c",
           980 => x"84",
           981 => x"51",
           982 => x"88",
           983 => x"87",
           984 => x"08",
           985 => x"84",
           986 => x"51",
           987 => x"73",
           988 => x"87",
           989 => x"0c",
           990 => x"0b",
           991 => x"84",
           992 => x"83",
           993 => x"94",
           994 => x"f8",
           995 => x"3f",
           996 => x"38",
           997 => x"fc",
           998 => x"08",
           999 => x"80",
          1000 => x"87",
          1001 => x"0c",
          1002 => x"fc",
          1003 => x"80",
          1004 => x"fc",
          1005 => x"08",
          1006 => x"54",
          1007 => x"86",
          1008 => x"55",
          1009 => x"80",
          1010 => x"80",
          1011 => x"00",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"00",
          1016 => x"54",
          1017 => x"59",
          1018 => x"4d",
          1019 => x"00",
          1020 => x"00",
          2048 => x"a4",
          2049 => x"0b",
          2050 => x"04",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"a4",
          2057 => x"0b",
          2058 => x"04",
          2059 => x"a4",
          2060 => x"0b",
          2061 => x"04",
          2062 => x"a4",
          2063 => x"0b",
          2064 => x"04",
          2065 => x"a4",
          2066 => x"0b",
          2067 => x"04",
          2068 => x"a4",
          2069 => x"0b",
          2070 => x"04",
          2071 => x"a5",
          2072 => x"0b",
          2073 => x"04",
          2074 => x"a5",
          2075 => x"0b",
          2076 => x"04",
          2077 => x"a5",
          2078 => x"0b",
          2079 => x"04",
          2080 => x"a5",
          2081 => x"0b",
          2082 => x"04",
          2083 => x"a6",
          2084 => x"0b",
          2085 => x"04",
          2086 => x"a6",
          2087 => x"0b",
          2088 => x"04",
          2089 => x"a6",
          2090 => x"0b",
          2091 => x"04",
          2092 => x"a6",
          2093 => x"0b",
          2094 => x"04",
          2095 => x"a7",
          2096 => x"0b",
          2097 => x"04",
          2098 => x"a7",
          2099 => x"0b",
          2100 => x"04",
          2101 => x"a7",
          2102 => x"0b",
          2103 => x"04",
          2104 => x"a7",
          2105 => x"0b",
          2106 => x"04",
          2107 => x"a8",
          2108 => x"0b",
          2109 => x"04",
          2110 => x"a8",
          2111 => x"0b",
          2112 => x"04",
          2113 => x"a8",
          2114 => x"0b",
          2115 => x"04",
          2116 => x"a8",
          2117 => x"0b",
          2118 => x"04",
          2119 => x"a9",
          2120 => x"0b",
          2121 => x"04",
          2122 => x"a9",
          2123 => x"0b",
          2124 => x"04",
          2125 => x"a9",
          2126 => x"0b",
          2127 => x"04",
          2128 => x"a9",
          2129 => x"0b",
          2130 => x"04",
          2131 => x"aa",
          2132 => x"0b",
          2133 => x"04",
          2134 => x"aa",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"04",
          2177 => x"0c",
          2178 => x"82",
          2179 => x"83",
          2180 => x"82",
          2181 => x"80",
          2182 => x"82",
          2183 => x"83",
          2184 => x"82",
          2185 => x"80",
          2186 => x"82",
          2187 => x"83",
          2188 => x"82",
          2189 => x"80",
          2190 => x"82",
          2191 => x"83",
          2192 => x"82",
          2193 => x"80",
          2194 => x"82",
          2195 => x"83",
          2196 => x"82",
          2197 => x"80",
          2198 => x"82",
          2199 => x"83",
          2200 => x"82",
          2201 => x"80",
          2202 => x"82",
          2203 => x"83",
          2204 => x"82",
          2205 => x"80",
          2206 => x"82",
          2207 => x"83",
          2208 => x"82",
          2209 => x"80",
          2210 => x"82",
          2211 => x"83",
          2212 => x"82",
          2213 => x"80",
          2214 => x"82",
          2215 => x"83",
          2216 => x"82",
          2217 => x"80",
          2218 => x"82",
          2219 => x"83",
          2220 => x"82",
          2221 => x"80",
          2222 => x"82",
          2223 => x"83",
          2224 => x"82",
          2225 => x"80",
          2226 => x"82",
          2227 => x"83",
          2228 => x"82",
          2229 => x"ba",
          2230 => x"93",
          2231 => x"80",
          2232 => x"93",
          2233 => x"fe",
          2234 => x"90",
          2235 => x"90",
          2236 => x"90",
          2237 => x"2d",
          2238 => x"08",
          2239 => x"04",
          2240 => x"0c",
          2241 => x"82",
          2242 => x"83",
          2243 => x"82",
          2244 => x"b6",
          2245 => x"93",
          2246 => x"80",
          2247 => x"93",
          2248 => x"98",
          2249 => x"93",
          2250 => x"80",
          2251 => x"93",
          2252 => x"a5",
          2253 => x"93",
          2254 => x"80",
          2255 => x"93",
          2256 => x"9d",
          2257 => x"93",
          2258 => x"80",
          2259 => x"93",
          2260 => x"a0",
          2261 => x"93",
          2262 => x"80",
          2263 => x"93",
          2264 => x"aa",
          2265 => x"93",
          2266 => x"80",
          2267 => x"93",
          2268 => x"b3",
          2269 => x"93",
          2270 => x"80",
          2271 => x"93",
          2272 => x"a4",
          2273 => x"93",
          2274 => x"80",
          2275 => x"93",
          2276 => x"ae",
          2277 => x"93",
          2278 => x"80",
          2279 => x"93",
          2280 => x"af",
          2281 => x"93",
          2282 => x"80",
          2283 => x"93",
          2284 => x"af",
          2285 => x"93",
          2286 => x"80",
          2287 => x"93",
          2288 => x"b7",
          2289 => x"93",
          2290 => x"80",
          2291 => x"93",
          2292 => x"b5",
          2293 => x"93",
          2294 => x"80",
          2295 => x"93",
          2296 => x"ba",
          2297 => x"93",
          2298 => x"80",
          2299 => x"93",
          2300 => x"b0",
          2301 => x"93",
          2302 => x"80",
          2303 => x"93",
          2304 => x"bd",
          2305 => x"93",
          2306 => x"80",
          2307 => x"93",
          2308 => x"be",
          2309 => x"93",
          2310 => x"80",
          2311 => x"93",
          2312 => x"a6",
          2313 => x"93",
          2314 => x"80",
          2315 => x"93",
          2316 => x"a6",
          2317 => x"93",
          2318 => x"80",
          2319 => x"93",
          2320 => x"a7",
          2321 => x"93",
          2322 => x"80",
          2323 => x"93",
          2324 => x"b1",
          2325 => x"93",
          2326 => x"80",
          2327 => x"93",
          2328 => x"be",
          2329 => x"93",
          2330 => x"80",
          2331 => x"93",
          2332 => x"c0",
          2333 => x"93",
          2334 => x"80",
          2335 => x"93",
          2336 => x"c4",
          2337 => x"93",
          2338 => x"80",
          2339 => x"93",
          2340 => x"98",
          2341 => x"93",
          2342 => x"80",
          2343 => x"93",
          2344 => x"c7",
          2345 => x"93",
          2346 => x"80",
          2347 => x"93",
          2348 => x"d5",
          2349 => x"93",
          2350 => x"80",
          2351 => x"93",
          2352 => x"d3",
          2353 => x"93",
          2354 => x"80",
          2355 => x"93",
          2356 => x"e9",
          2357 => x"93",
          2358 => x"80",
          2359 => x"93",
          2360 => x"eb",
          2361 => x"93",
          2362 => x"80",
          2363 => x"93",
          2364 => x"ed",
          2365 => x"93",
          2366 => x"80",
          2367 => x"93",
          2368 => x"c3",
          2369 => x"90",
          2370 => x"90",
          2371 => x"90",
          2372 => x"2d",
          2373 => x"08",
          2374 => x"04",
          2375 => x"0c",
          2376 => x"82",
          2377 => x"83",
          2378 => x"82",
          2379 => x"81",
          2380 => x"82",
          2381 => x"83",
          2382 => x"82",
          2383 => x"82",
          2384 => x"8e",
          2385 => x"70",
          2386 => x"0c",
          2387 => x"aa",
          2388 => x"80",
          2389 => x"a3",
          2390 => x"82",
          2391 => x"02",
          2392 => x"0c",
          2393 => x"80",
          2394 => x"90",
          2395 => x"08",
          2396 => x"90",
          2397 => x"08",
          2398 => x"3f",
          2399 => x"08",
          2400 => x"84",
          2401 => x"3d",
          2402 => x"90",
          2403 => x"93",
          2404 => x"82",
          2405 => x"fd",
          2406 => x"53",
          2407 => x"08",
          2408 => x"52",
          2409 => x"08",
          2410 => x"51",
          2411 => x"93",
          2412 => x"82",
          2413 => x"54",
          2414 => x"82",
          2415 => x"04",
          2416 => x"08",
          2417 => x"90",
          2418 => x"0d",
          2419 => x"93",
          2420 => x"05",
          2421 => x"82",
          2422 => x"f8",
          2423 => x"93",
          2424 => x"05",
          2425 => x"90",
          2426 => x"08",
          2427 => x"82",
          2428 => x"fc",
          2429 => x"2e",
          2430 => x"0b",
          2431 => x"08",
          2432 => x"24",
          2433 => x"93",
          2434 => x"05",
          2435 => x"93",
          2436 => x"05",
          2437 => x"90",
          2438 => x"08",
          2439 => x"90",
          2440 => x"0c",
          2441 => x"82",
          2442 => x"fc",
          2443 => x"2e",
          2444 => x"82",
          2445 => x"8c",
          2446 => x"93",
          2447 => x"05",
          2448 => x"38",
          2449 => x"08",
          2450 => x"82",
          2451 => x"8c",
          2452 => x"82",
          2453 => x"88",
          2454 => x"93",
          2455 => x"05",
          2456 => x"90",
          2457 => x"08",
          2458 => x"90",
          2459 => x"0c",
          2460 => x"08",
          2461 => x"81",
          2462 => x"90",
          2463 => x"0c",
          2464 => x"08",
          2465 => x"81",
          2466 => x"90",
          2467 => x"0c",
          2468 => x"82",
          2469 => x"90",
          2470 => x"2e",
          2471 => x"93",
          2472 => x"05",
          2473 => x"93",
          2474 => x"05",
          2475 => x"39",
          2476 => x"08",
          2477 => x"70",
          2478 => x"08",
          2479 => x"51",
          2480 => x"08",
          2481 => x"82",
          2482 => x"85",
          2483 => x"93",
          2484 => x"fc",
          2485 => x"70",
          2486 => x"55",
          2487 => x"72",
          2488 => x"72",
          2489 => x"06",
          2490 => x"2e",
          2491 => x"12",
          2492 => x"2e",
          2493 => x"70",
          2494 => x"33",
          2495 => x"05",
          2496 => x"12",
          2497 => x"2e",
          2498 => x"ea",
          2499 => x"93",
          2500 => x"3d",
          2501 => x"51",
          2502 => x"05",
          2503 => x"70",
          2504 => x"0c",
          2505 => x"05",
          2506 => x"70",
          2507 => x"0c",
          2508 => x"05",
          2509 => x"70",
          2510 => x"0c",
          2511 => x"05",
          2512 => x"70",
          2513 => x"0c",
          2514 => x"71",
          2515 => x"38",
          2516 => x"95",
          2517 => x"84",
          2518 => x"71",
          2519 => x"53",
          2520 => x"52",
          2521 => x"ed",
          2522 => x"ff",
          2523 => x"3d",
          2524 => x"71",
          2525 => x"9f",
          2526 => x"55",
          2527 => x"72",
          2528 => x"74",
          2529 => x"70",
          2530 => x"38",
          2531 => x"71",
          2532 => x"38",
          2533 => x"81",
          2534 => x"ff",
          2535 => x"ff",
          2536 => x"06",
          2537 => x"82",
          2538 => x"86",
          2539 => x"74",
          2540 => x"75",
          2541 => x"90",
          2542 => x"54",
          2543 => x"27",
          2544 => x"71",
          2545 => x"53",
          2546 => x"70",
          2547 => x"0c",
          2548 => x"84",
          2549 => x"72",
          2550 => x"05",
          2551 => x"12",
          2552 => x"26",
          2553 => x"72",
          2554 => x"72",
          2555 => x"05",
          2556 => x"12",
          2557 => x"26",
          2558 => x"53",
          2559 => x"fc",
          2560 => x"70",
          2561 => x"07",
          2562 => x"54",
          2563 => x"80",
          2564 => x"70",
          2565 => x"70",
          2566 => x"ff",
          2567 => x"f8",
          2568 => x"80",
          2569 => x"53",
          2570 => x"a6",
          2571 => x"72",
          2572 => x"05",
          2573 => x"08",
          2574 => x"f7",
          2575 => x"13",
          2576 => x"84",
          2577 => x"06",
          2578 => x"53",
          2579 => x"2e",
          2580 => x"52",
          2581 => x"05",
          2582 => x"70",
          2583 => x"05",
          2584 => x"f0",
          2585 => x"93",
          2586 => x"3d",
          2587 => x"3d",
          2588 => x"71",
          2589 => x"55",
          2590 => x"38",
          2591 => x"70",
          2592 => x"fd",
          2593 => x"70",
          2594 => x"81",
          2595 => x"51",
          2596 => x"9d",
          2597 => x"70",
          2598 => x"f7",
          2599 => x"12",
          2600 => x"84",
          2601 => x"06",
          2602 => x"53",
          2603 => x"e5",
          2604 => x"71",
          2605 => x"80",
          2606 => x"81",
          2607 => x"52",
          2608 => x"38",
          2609 => x"82",
          2610 => x"85",
          2611 => x"fa",
          2612 => x"7a",
          2613 => x"55",
          2614 => x"80",
          2615 => x"38",
          2616 => x"83",
          2617 => x"80",
          2618 => x"38",
          2619 => x"72",
          2620 => x"38",
          2621 => x"33",
          2622 => x"71",
          2623 => x"06",
          2624 => x"80",
          2625 => x"38",
          2626 => x"06",
          2627 => x"2e",
          2628 => x"81",
          2629 => x"ff",
          2630 => x"52",
          2631 => x"09",
          2632 => x"38",
          2633 => x"33",
          2634 => x"81",
          2635 => x"81",
          2636 => x"71",
          2637 => x"52",
          2638 => x"84",
          2639 => x"0d",
          2640 => x"57",
          2641 => x"27",
          2642 => x"08",
          2643 => x"88",
          2644 => x"55",
          2645 => x"39",
          2646 => x"72",
          2647 => x"38",
          2648 => x"09",
          2649 => x"ff",
          2650 => x"f8",
          2651 => x"80",
          2652 => x"51",
          2653 => x"84",
          2654 => x"57",
          2655 => x"27",
          2656 => x"08",
          2657 => x"d0",
          2658 => x"55",
          2659 => x"39",
          2660 => x"93",
          2661 => x"3d",
          2662 => x"3d",
          2663 => x"83",
          2664 => x"2b",
          2665 => x"3f",
          2666 => x"08",
          2667 => x"72",
          2668 => x"54",
          2669 => x"25",
          2670 => x"82",
          2671 => x"84",
          2672 => x"fb",
          2673 => x"70",
          2674 => x"53",
          2675 => x"2e",
          2676 => x"71",
          2677 => x"a0",
          2678 => x"06",
          2679 => x"12",
          2680 => x"71",
          2681 => x"81",
          2682 => x"73",
          2683 => x"ff",
          2684 => x"55",
          2685 => x"83",
          2686 => x"70",
          2687 => x"38",
          2688 => x"73",
          2689 => x"51",
          2690 => x"09",
          2691 => x"38",
          2692 => x"81",
          2693 => x"72",
          2694 => x"51",
          2695 => x"84",
          2696 => x"0d",
          2697 => x"0d",
          2698 => x"08",
          2699 => x"38",
          2700 => x"05",
          2701 => x"9f",
          2702 => x"93",
          2703 => x"38",
          2704 => x"39",
          2705 => x"82",
          2706 => x"86",
          2707 => x"fc",
          2708 => x"82",
          2709 => x"05",
          2710 => x"52",
          2711 => x"81",
          2712 => x"13",
          2713 => x"51",
          2714 => x"9e",
          2715 => x"38",
          2716 => x"51",
          2717 => x"97",
          2718 => x"38",
          2719 => x"51",
          2720 => x"bb",
          2721 => x"38",
          2722 => x"51",
          2723 => x"bb",
          2724 => x"38",
          2725 => x"55",
          2726 => x"87",
          2727 => x"d9",
          2728 => x"22",
          2729 => x"73",
          2730 => x"80",
          2731 => x"0b",
          2732 => x"9c",
          2733 => x"87",
          2734 => x"0c",
          2735 => x"87",
          2736 => x"0c",
          2737 => x"87",
          2738 => x"0c",
          2739 => x"87",
          2740 => x"0c",
          2741 => x"87",
          2742 => x"0c",
          2743 => x"87",
          2744 => x"0c",
          2745 => x"98",
          2746 => x"87",
          2747 => x"0c",
          2748 => x"c0",
          2749 => x"80",
          2750 => x"93",
          2751 => x"3d",
          2752 => x"3d",
          2753 => x"87",
          2754 => x"5d",
          2755 => x"87",
          2756 => x"08",
          2757 => x"23",
          2758 => x"b8",
          2759 => x"82",
          2760 => x"c0",
          2761 => x"5a",
          2762 => x"34",
          2763 => x"b0",
          2764 => x"84",
          2765 => x"c0",
          2766 => x"5a",
          2767 => x"34",
          2768 => x"a8",
          2769 => x"86",
          2770 => x"c0",
          2771 => x"5c",
          2772 => x"23",
          2773 => x"a0",
          2774 => x"8a",
          2775 => x"7d",
          2776 => x"ff",
          2777 => x"7b",
          2778 => x"06",
          2779 => x"33",
          2780 => x"33",
          2781 => x"33",
          2782 => x"33",
          2783 => x"33",
          2784 => x"ff",
          2785 => x"81",
          2786 => x"99",
          2787 => x"3d",
          2788 => x"3d",
          2789 => x"05",
          2790 => x"70",
          2791 => x"52",
          2792 => x"0b",
          2793 => x"34",
          2794 => x"04",
          2795 => x"77",
          2796 => x"8d",
          2797 => x"81",
          2798 => x"55",
          2799 => x"94",
          2800 => x"80",
          2801 => x"87",
          2802 => x"51",
          2803 => x"96",
          2804 => x"06",
          2805 => x"70",
          2806 => x"38",
          2807 => x"70",
          2808 => x"51",
          2809 => x"72",
          2810 => x"81",
          2811 => x"70",
          2812 => x"38",
          2813 => x"70",
          2814 => x"51",
          2815 => x"38",
          2816 => x"06",
          2817 => x"94",
          2818 => x"80",
          2819 => x"87",
          2820 => x"52",
          2821 => x"75",
          2822 => x"0c",
          2823 => x"04",
          2824 => x"02",
          2825 => x"0b",
          2826 => x"fc",
          2827 => x"ff",
          2828 => x"56",
          2829 => x"84",
          2830 => x"2e",
          2831 => x"c0",
          2832 => x"70",
          2833 => x"2a",
          2834 => x"53",
          2835 => x"80",
          2836 => x"71",
          2837 => x"81",
          2838 => x"70",
          2839 => x"81",
          2840 => x"06",
          2841 => x"80",
          2842 => x"71",
          2843 => x"81",
          2844 => x"70",
          2845 => x"73",
          2846 => x"51",
          2847 => x"80",
          2848 => x"2e",
          2849 => x"c0",
          2850 => x"75",
          2851 => x"3d",
          2852 => x"3d",
          2853 => x"80",
          2854 => x"81",
          2855 => x"53",
          2856 => x"2e",
          2857 => x"71",
          2858 => x"81",
          2859 => x"82",
          2860 => x"70",
          2861 => x"59",
          2862 => x"87",
          2863 => x"51",
          2864 => x"86",
          2865 => x"94",
          2866 => x"08",
          2867 => x"70",
          2868 => x"54",
          2869 => x"2e",
          2870 => x"91",
          2871 => x"06",
          2872 => x"d7",
          2873 => x"32",
          2874 => x"51",
          2875 => x"2e",
          2876 => x"93",
          2877 => x"06",
          2878 => x"ff",
          2879 => x"81",
          2880 => x"87",
          2881 => x"52",
          2882 => x"86",
          2883 => x"94",
          2884 => x"72",
          2885 => x"74",
          2886 => x"ff",
          2887 => x"57",
          2888 => x"38",
          2889 => x"84",
          2890 => x"0d",
          2891 => x"0d",
          2892 => x"8d",
          2893 => x"81",
          2894 => x"52",
          2895 => x"84",
          2896 => x"2e",
          2897 => x"c0",
          2898 => x"70",
          2899 => x"2a",
          2900 => x"51",
          2901 => x"80",
          2902 => x"71",
          2903 => x"51",
          2904 => x"80",
          2905 => x"2e",
          2906 => x"c0",
          2907 => x"71",
          2908 => x"ff",
          2909 => x"84",
          2910 => x"3d",
          2911 => x"3d",
          2912 => x"82",
          2913 => x"70",
          2914 => x"52",
          2915 => x"94",
          2916 => x"80",
          2917 => x"87",
          2918 => x"52",
          2919 => x"82",
          2920 => x"06",
          2921 => x"ff",
          2922 => x"2e",
          2923 => x"81",
          2924 => x"87",
          2925 => x"52",
          2926 => x"86",
          2927 => x"94",
          2928 => x"08",
          2929 => x"70",
          2930 => x"53",
          2931 => x"93",
          2932 => x"3d",
          2933 => x"3d",
          2934 => x"9e",
          2935 => x"9c",
          2936 => x"51",
          2937 => x"2e",
          2938 => x"87",
          2939 => x"08",
          2940 => x"0c",
          2941 => x"a8",
          2942 => x"84",
          2943 => x"9e",
          2944 => x"8e",
          2945 => x"c0",
          2946 => x"82",
          2947 => x"87",
          2948 => x"08",
          2949 => x"0c",
          2950 => x"a0",
          2951 => x"94",
          2952 => x"9e",
          2953 => x"8e",
          2954 => x"c0",
          2955 => x"82",
          2956 => x"87",
          2957 => x"08",
          2958 => x"0c",
          2959 => x"b8",
          2960 => x"a4",
          2961 => x"9e",
          2962 => x"8e",
          2963 => x"c0",
          2964 => x"82",
          2965 => x"87",
          2966 => x"08",
          2967 => x"0c",
          2968 => x"80",
          2969 => x"82",
          2970 => x"87",
          2971 => x"08",
          2972 => x"0c",
          2973 => x"88",
          2974 => x"bc",
          2975 => x"9e",
          2976 => x"8e",
          2977 => x"0b",
          2978 => x"34",
          2979 => x"c0",
          2980 => x"70",
          2981 => x"06",
          2982 => x"70",
          2983 => x"38",
          2984 => x"82",
          2985 => x"80",
          2986 => x"9e",
          2987 => x"88",
          2988 => x"51",
          2989 => x"80",
          2990 => x"81",
          2991 => x"8e",
          2992 => x"0b",
          2993 => x"90",
          2994 => x"80",
          2995 => x"52",
          2996 => x"2e",
          2997 => x"52",
          2998 => x"c7",
          2999 => x"87",
          3000 => x"08",
          3001 => x"80",
          3002 => x"52",
          3003 => x"83",
          3004 => x"71",
          3005 => x"34",
          3006 => x"c0",
          3007 => x"70",
          3008 => x"06",
          3009 => x"70",
          3010 => x"38",
          3011 => x"82",
          3012 => x"80",
          3013 => x"9e",
          3014 => x"90",
          3015 => x"51",
          3016 => x"80",
          3017 => x"81",
          3018 => x"8e",
          3019 => x"0b",
          3020 => x"90",
          3021 => x"80",
          3022 => x"52",
          3023 => x"2e",
          3024 => x"52",
          3025 => x"cb",
          3026 => x"87",
          3027 => x"08",
          3028 => x"80",
          3029 => x"52",
          3030 => x"83",
          3031 => x"71",
          3032 => x"34",
          3033 => x"c0",
          3034 => x"70",
          3035 => x"06",
          3036 => x"70",
          3037 => x"38",
          3038 => x"82",
          3039 => x"80",
          3040 => x"9e",
          3041 => x"80",
          3042 => x"51",
          3043 => x"80",
          3044 => x"81",
          3045 => x"8e",
          3046 => x"0b",
          3047 => x"90",
          3048 => x"80",
          3049 => x"52",
          3050 => x"83",
          3051 => x"71",
          3052 => x"34",
          3053 => x"90",
          3054 => x"80",
          3055 => x"2a",
          3056 => x"70",
          3057 => x"34",
          3058 => x"c0",
          3059 => x"70",
          3060 => x"51",
          3061 => x"80",
          3062 => x"81",
          3063 => x"8e",
          3064 => x"c0",
          3065 => x"70",
          3066 => x"70",
          3067 => x"51",
          3068 => x"8e",
          3069 => x"0b",
          3070 => x"90",
          3071 => x"06",
          3072 => x"70",
          3073 => x"38",
          3074 => x"82",
          3075 => x"87",
          3076 => x"08",
          3077 => x"51",
          3078 => x"8e",
          3079 => x"3d",
          3080 => x"3d",
          3081 => x"80",
          3082 => x"3f",
          3083 => x"33",
          3084 => x"2e",
          3085 => x"f7",
          3086 => x"8c",
          3087 => x"a8",
          3088 => x"3f",
          3089 => x"33",
          3090 => x"2e",
          3091 => x"8e",
          3092 => x"8e",
          3093 => x"54",
          3094 => x"c0",
          3095 => x"3f",
          3096 => x"33",
          3097 => x"2e",
          3098 => x"8e",
          3099 => x"8e",
          3100 => x"54",
          3101 => x"dc",
          3102 => x"3f",
          3103 => x"33",
          3104 => x"2e",
          3105 => x"8e",
          3106 => x"8e",
          3107 => x"54",
          3108 => x"f8",
          3109 => x"3f",
          3110 => x"33",
          3111 => x"2e",
          3112 => x"8e",
          3113 => x"8e",
          3114 => x"54",
          3115 => x"94",
          3116 => x"3f",
          3117 => x"33",
          3118 => x"2e",
          3119 => x"8e",
          3120 => x"8e",
          3121 => x"54",
          3122 => x"b0",
          3123 => x"3f",
          3124 => x"33",
          3125 => x"2e",
          3126 => x"8e",
          3127 => x"81",
          3128 => x"8e",
          3129 => x"8e",
          3130 => x"73",
          3131 => x"38",
          3132 => x"33",
          3133 => x"ec",
          3134 => x"3f",
          3135 => x"33",
          3136 => x"2e",
          3137 => x"8e",
          3138 => x"81",
          3139 => x"8e",
          3140 => x"8e",
          3141 => x"73",
          3142 => x"38",
          3143 => x"51",
          3144 => x"82",
          3145 => x"54",
          3146 => x"88",
          3147 => x"c0",
          3148 => x"3f",
          3149 => x"33",
          3150 => x"2e",
          3151 => x"f9",
          3152 => x"84",
          3153 => x"cd",
          3154 => x"80",
          3155 => x"81",
          3156 => x"87",
          3157 => x"8e",
          3158 => x"73",
          3159 => x"38",
          3160 => x"51",
          3161 => x"81",
          3162 => x"87",
          3163 => x"8e",
          3164 => x"81",
          3165 => x"8d",
          3166 => x"8e",
          3167 => x"81",
          3168 => x"8d",
          3169 => x"8e",
          3170 => x"81",
          3171 => x"8d",
          3172 => x"fa",
          3173 => x"b0",
          3174 => x"b4",
          3175 => x"fa",
          3176 => x"88",
          3177 => x"b8",
          3178 => x"84",
          3179 => x"51",
          3180 => x"82",
          3181 => x"bd",
          3182 => x"76",
          3183 => x"54",
          3184 => x"08",
          3185 => x"a4",
          3186 => x"3f",
          3187 => x"33",
          3188 => x"2e",
          3189 => x"8e",
          3190 => x"bd",
          3191 => x"75",
          3192 => x"3f",
          3193 => x"08",
          3194 => x"29",
          3195 => x"54",
          3196 => x"84",
          3197 => x"fb",
          3198 => x"b0",
          3199 => x"c6",
          3200 => x"80",
          3201 => x"82",
          3202 => x"56",
          3203 => x"52",
          3204 => x"c7",
          3205 => x"84",
          3206 => x"c0",
          3207 => x"31",
          3208 => x"93",
          3209 => x"81",
          3210 => x"8b",
          3211 => x"89",
          3212 => x"94",
          3213 => x"0d",
          3214 => x"0d",
          3215 => x"33",
          3216 => x"71",
          3217 => x"38",
          3218 => x"0b",
          3219 => x"d4",
          3220 => x"08",
          3221 => x"a8",
          3222 => x"81",
          3223 => x"97",
          3224 => x"b8",
          3225 => x"81",
          3226 => x"8b",
          3227 => x"c4",
          3228 => x"81",
          3229 => x"85",
          3230 => x"3d",
          3231 => x"88",
          3232 => x"ff",
          3233 => x"c0",
          3234 => x"08",
          3235 => x"72",
          3236 => x"07",
          3237 => x"d8",
          3238 => x"83",
          3239 => x"ff",
          3240 => x"c0",
          3241 => x"08",
          3242 => x"0c",
          3243 => x"0c",
          3244 => x"82",
          3245 => x"06",
          3246 => x"d8",
          3247 => x"51",
          3248 => x"04",
          3249 => x"c0",
          3250 => x"04",
          3251 => x"08",
          3252 => x"84",
          3253 => x"3d",
          3254 => x"94",
          3255 => x"82",
          3256 => x"82",
          3257 => x"82",
          3258 => x"75",
          3259 => x"ff",
          3260 => x"b7",
          3261 => x"38",
          3262 => x"94",
          3263 => x"72",
          3264 => x"0c",
          3265 => x"04",
          3266 => x"79",
          3267 => x"08",
          3268 => x"14",
          3269 => x"08",
          3270 => x"5a",
          3271 => x"57",
          3272 => x"26",
          3273 => x"13",
          3274 => x"53",
          3275 => x"0c",
          3276 => x"84",
          3277 => x"73",
          3278 => x"14",
          3279 => x"12",
          3280 => x"12",
          3281 => x"13",
          3282 => x"14",
          3283 => x"12",
          3284 => x"12",
          3285 => x"15",
          3286 => x"16",
          3287 => x"80",
          3288 => x"90",
          3289 => x"94",
          3290 => x"82",
          3291 => x"89",
          3292 => x"fc",
          3293 => x"8c",
          3294 => x"12",
          3295 => x"53",
          3296 => x"2e",
          3297 => x"a3",
          3298 => x"08",
          3299 => x"55",
          3300 => x"09",
          3301 => x"38",
          3302 => x"15",
          3303 => x"73",
          3304 => x"71",
          3305 => x"71",
          3306 => x"81",
          3307 => x"8e",
          3308 => x"14",
          3309 => x"dc",
          3310 => x"0c",
          3311 => x"ec",
          3312 => x"08",
          3313 => x"0c",
          3314 => x"81",
          3315 => x"06",
          3316 => x"13",
          3317 => x"52",
          3318 => x"2e",
          3319 => x"a4",
          3320 => x"08",
          3321 => x"0c",
          3322 => x"90",
          3323 => x"90",
          3324 => x"94",
          3325 => x"14",
          3326 => x"08",
          3327 => x"0c",
          3328 => x"0c",
          3329 => x"84",
          3330 => x"0d",
          3331 => x"0d",
          3332 => x"57",
          3333 => x"81",
          3334 => x"17",
          3335 => x"8e",
          3336 => x"57",
          3337 => x"2e",
          3338 => x"16",
          3339 => x"80",
          3340 => x"16",
          3341 => x"39",
          3342 => x"17",
          3343 => x"06",
          3344 => x"fd",
          3345 => x"93",
          3346 => x"93",
          3347 => x"70",
          3348 => x"08",
          3349 => x"82",
          3350 => x"09",
          3351 => x"72",
          3352 => x"73",
          3353 => x"58",
          3354 => x"80",
          3355 => x"2e",
          3356 => x"80",
          3357 => x"39",
          3358 => x"51",
          3359 => x"81",
          3360 => x"84",
          3361 => x"82",
          3362 => x"84",
          3363 => x"8e",
          3364 => x"72",
          3365 => x"8c",
          3366 => x"26",
          3367 => x"13",
          3368 => x"39",
          3369 => x"88",
          3370 => x"8c",
          3371 => x"88",
          3372 => x"16",
          3373 => x"12",
          3374 => x"51",
          3375 => x"76",
          3376 => x"84",
          3377 => x"c0",
          3378 => x"84",
          3379 => x"82",
          3380 => x"89",
          3381 => x"ff",
          3382 => x"52",
          3383 => x"87",
          3384 => x"51",
          3385 => x"83",
          3386 => x"fe",
          3387 => x"93",
          3388 => x"72",
          3389 => x"81",
          3390 => x"8d",
          3391 => x"82",
          3392 => x"52",
          3393 => x"90",
          3394 => x"34",
          3395 => x"08",
          3396 => x"93",
          3397 => x"39",
          3398 => x"08",
          3399 => x"2e",
          3400 => x"51",
          3401 => x"3d",
          3402 => x"3d",
          3403 => x"05",
          3404 => x"98",
          3405 => x"93",
          3406 => x"51",
          3407 => x"72",
          3408 => x"0c",
          3409 => x"04",
          3410 => x"75",
          3411 => x"70",
          3412 => x"53",
          3413 => x"2e",
          3414 => x"81",
          3415 => x"81",
          3416 => x"87",
          3417 => x"85",
          3418 => x"fc",
          3419 => x"82",
          3420 => x"78",
          3421 => x"0c",
          3422 => x"33",
          3423 => x"06",
          3424 => x"80",
          3425 => x"72",
          3426 => x"51",
          3427 => x"fe",
          3428 => x"39",
          3429 => x"98",
          3430 => x"0d",
          3431 => x"0d",
          3432 => x"59",
          3433 => x"05",
          3434 => x"75",
          3435 => x"f8",
          3436 => x"2e",
          3437 => x"82",
          3438 => x"70",
          3439 => x"05",
          3440 => x"5b",
          3441 => x"2e",
          3442 => x"85",
          3443 => x"8b",
          3444 => x"2e",
          3445 => x"8a",
          3446 => x"78",
          3447 => x"5a",
          3448 => x"aa",
          3449 => x"06",
          3450 => x"84",
          3451 => x"7b",
          3452 => x"5d",
          3453 => x"59",
          3454 => x"d0",
          3455 => x"89",
          3456 => x"7a",
          3457 => x"10",
          3458 => x"d0",
          3459 => x"81",
          3460 => x"57",
          3461 => x"75",
          3462 => x"70",
          3463 => x"07",
          3464 => x"80",
          3465 => x"30",
          3466 => x"80",
          3467 => x"53",
          3468 => x"55",
          3469 => x"2e",
          3470 => x"84",
          3471 => x"81",
          3472 => x"57",
          3473 => x"2e",
          3474 => x"75",
          3475 => x"76",
          3476 => x"e0",
          3477 => x"ff",
          3478 => x"73",
          3479 => x"81",
          3480 => x"80",
          3481 => x"38",
          3482 => x"2e",
          3483 => x"73",
          3484 => x"8b",
          3485 => x"c2",
          3486 => x"38",
          3487 => x"73",
          3488 => x"81",
          3489 => x"8f",
          3490 => x"d5",
          3491 => x"38",
          3492 => x"24",
          3493 => x"80",
          3494 => x"38",
          3495 => x"73",
          3496 => x"80",
          3497 => x"ef",
          3498 => x"19",
          3499 => x"59",
          3500 => x"33",
          3501 => x"75",
          3502 => x"81",
          3503 => x"70",
          3504 => x"55",
          3505 => x"79",
          3506 => x"90",
          3507 => x"16",
          3508 => x"7b",
          3509 => x"a0",
          3510 => x"3f",
          3511 => x"53",
          3512 => x"e9",
          3513 => x"fc",
          3514 => x"81",
          3515 => x"72",
          3516 => x"b0",
          3517 => x"fb",
          3518 => x"39",
          3519 => x"83",
          3520 => x"59",
          3521 => x"82",
          3522 => x"88",
          3523 => x"8a",
          3524 => x"90",
          3525 => x"75",
          3526 => x"3f",
          3527 => x"79",
          3528 => x"81",
          3529 => x"72",
          3530 => x"38",
          3531 => x"59",
          3532 => x"84",
          3533 => x"58",
          3534 => x"80",
          3535 => x"30",
          3536 => x"80",
          3537 => x"55",
          3538 => x"25",
          3539 => x"80",
          3540 => x"74",
          3541 => x"07",
          3542 => x"0b",
          3543 => x"57",
          3544 => x"51",
          3545 => x"82",
          3546 => x"81",
          3547 => x"53",
          3548 => x"db",
          3549 => x"93",
          3550 => x"89",
          3551 => x"38",
          3552 => x"75",
          3553 => x"84",
          3554 => x"53",
          3555 => x"06",
          3556 => x"53",
          3557 => x"81",
          3558 => x"81",
          3559 => x"70",
          3560 => x"2a",
          3561 => x"76",
          3562 => x"38",
          3563 => x"38",
          3564 => x"70",
          3565 => x"53",
          3566 => x"8e",
          3567 => x"77",
          3568 => x"53",
          3569 => x"81",
          3570 => x"7a",
          3571 => x"55",
          3572 => x"83",
          3573 => x"79",
          3574 => x"81",
          3575 => x"72",
          3576 => x"17",
          3577 => x"27",
          3578 => x"51",
          3579 => x"75",
          3580 => x"72",
          3581 => x"81",
          3582 => x"7a",
          3583 => x"38",
          3584 => x"05",
          3585 => x"ff",
          3586 => x"70",
          3587 => x"57",
          3588 => x"76",
          3589 => x"81",
          3590 => x"72",
          3591 => x"84",
          3592 => x"f9",
          3593 => x"39",
          3594 => x"04",
          3595 => x"86",
          3596 => x"84",
          3597 => x"55",
          3598 => x"fa",
          3599 => x"3d",
          3600 => x"3d",
          3601 => x"93",
          3602 => x"3d",
          3603 => x"75",
          3604 => x"3f",
          3605 => x"08",
          3606 => x"34",
          3607 => x"93",
          3608 => x"3d",
          3609 => x"3d",
          3610 => x"98",
          3611 => x"93",
          3612 => x"3d",
          3613 => x"77",
          3614 => x"a1",
          3615 => x"93",
          3616 => x"3d",
          3617 => x"3d",
          3618 => x"82",
          3619 => x"70",
          3620 => x"55",
          3621 => x"80",
          3622 => x"38",
          3623 => x"08",
          3624 => x"82",
          3625 => x"81",
          3626 => x"72",
          3627 => x"cb",
          3628 => x"2e",
          3629 => x"88",
          3630 => x"70",
          3631 => x"51",
          3632 => x"2e",
          3633 => x"80",
          3634 => x"ff",
          3635 => x"39",
          3636 => x"c8",
          3637 => x"52",
          3638 => x"c0",
          3639 => x"52",
          3640 => x"81",
          3641 => x"51",
          3642 => x"ff",
          3643 => x"15",
          3644 => x"34",
          3645 => x"f3",
          3646 => x"72",
          3647 => x"0c",
          3648 => x"04",
          3649 => x"82",
          3650 => x"75",
          3651 => x"0c",
          3652 => x"52",
          3653 => x"3f",
          3654 => x"9c",
          3655 => x"0d",
          3656 => x"0d",
          3657 => x"56",
          3658 => x"0c",
          3659 => x"70",
          3660 => x"73",
          3661 => x"81",
          3662 => x"81",
          3663 => x"ed",
          3664 => x"2e",
          3665 => x"8e",
          3666 => x"08",
          3667 => x"76",
          3668 => x"56",
          3669 => x"b0",
          3670 => x"06",
          3671 => x"75",
          3672 => x"76",
          3673 => x"70",
          3674 => x"73",
          3675 => x"8b",
          3676 => x"73",
          3677 => x"85",
          3678 => x"82",
          3679 => x"76",
          3680 => x"70",
          3681 => x"ac",
          3682 => x"a0",
          3683 => x"fa",
          3684 => x"53",
          3685 => x"57",
          3686 => x"98",
          3687 => x"39",
          3688 => x"80",
          3689 => x"26",
          3690 => x"86",
          3691 => x"80",
          3692 => x"57",
          3693 => x"74",
          3694 => x"38",
          3695 => x"27",
          3696 => x"14",
          3697 => x"06",
          3698 => x"14",
          3699 => x"06",
          3700 => x"74",
          3701 => x"f9",
          3702 => x"ff",
          3703 => x"89",
          3704 => x"38",
          3705 => x"c5",
          3706 => x"29",
          3707 => x"81",
          3708 => x"76",
          3709 => x"56",
          3710 => x"ba",
          3711 => x"2e",
          3712 => x"30",
          3713 => x"0c",
          3714 => x"82",
          3715 => x"8a",
          3716 => x"f8",
          3717 => x"7c",
          3718 => x"70",
          3719 => x"75",
          3720 => x"55",
          3721 => x"2e",
          3722 => x"87",
          3723 => x"76",
          3724 => x"73",
          3725 => x"81",
          3726 => x"81",
          3727 => x"77",
          3728 => x"70",
          3729 => x"58",
          3730 => x"09",
          3731 => x"c2",
          3732 => x"81",
          3733 => x"75",
          3734 => x"55",
          3735 => x"e2",
          3736 => x"90",
          3737 => x"f8",
          3738 => x"8f",
          3739 => x"81",
          3740 => x"75",
          3741 => x"55",
          3742 => x"81",
          3743 => x"27",
          3744 => x"d0",
          3745 => x"55",
          3746 => x"73",
          3747 => x"80",
          3748 => x"14",
          3749 => x"72",
          3750 => x"e0",
          3751 => x"80",
          3752 => x"39",
          3753 => x"55",
          3754 => x"80",
          3755 => x"e0",
          3756 => x"38",
          3757 => x"81",
          3758 => x"53",
          3759 => x"81",
          3760 => x"53",
          3761 => x"8e",
          3762 => x"70",
          3763 => x"55",
          3764 => x"27",
          3765 => x"77",
          3766 => x"74",
          3767 => x"76",
          3768 => x"77",
          3769 => x"70",
          3770 => x"55",
          3771 => x"77",
          3772 => x"38",
          3773 => x"74",
          3774 => x"55",
          3775 => x"84",
          3776 => x"0d",
          3777 => x"0d",
          3778 => x"70",
          3779 => x"98",
          3780 => x"2c",
          3781 => x"70",
          3782 => x"53",
          3783 => x"51",
          3784 => x"fd",
          3785 => x"55",
          3786 => x"25",
          3787 => x"fd",
          3788 => x"12",
          3789 => x"97",
          3790 => x"33",
          3791 => x"70",
          3792 => x"81",
          3793 => x"81",
          3794 => x"93",
          3795 => x"3d",
          3796 => x"3d",
          3797 => x"84",
          3798 => x"33",
          3799 => x"55",
          3800 => x"2e",
          3801 => x"51",
          3802 => x"a0",
          3803 => x"3f",
          3804 => x"f7",
          3805 => x"ff",
          3806 => x"73",
          3807 => x"ff",
          3808 => x"39",
          3809 => x"c0",
          3810 => x"34",
          3811 => x"04",
          3812 => x"7c",
          3813 => x"b7",
          3814 => x"88",
          3815 => x"33",
          3816 => x"33",
          3817 => x"82",
          3818 => x"70",
          3819 => x"59",
          3820 => x"74",
          3821 => x"38",
          3822 => x"9b",
          3823 => x"d0",
          3824 => x"29",
          3825 => x"05",
          3826 => x"54",
          3827 => x"f0",
          3828 => x"93",
          3829 => x"0c",
          3830 => x"33",
          3831 => x"82",
          3832 => x"70",
          3833 => x"5a",
          3834 => x"a6",
          3835 => x"78",
          3836 => x"d5",
          3837 => x"8f",
          3838 => x"05",
          3839 => x"8f",
          3840 => x"81",
          3841 => x"93",
          3842 => x"38",
          3843 => x"8f",
          3844 => x"80",
          3845 => x"82",
          3846 => x"56",
          3847 => x"ac",
          3848 => x"c8",
          3849 => x"a4",
          3850 => x"fc",
          3851 => x"53",
          3852 => x"51",
          3853 => x"3f",
          3854 => x"08",
          3855 => x"80",
          3856 => x"82",
          3857 => x"51",
          3858 => x"3f",
          3859 => x"04",
          3860 => x"81",
          3861 => x"82",
          3862 => x"51",
          3863 => x"3f",
          3864 => x"08",
          3865 => x"82",
          3866 => x"53",
          3867 => x"88",
          3868 => x"56",
          3869 => x"3f",
          3870 => x"08",
          3871 => x"38",
          3872 => x"ea",
          3873 => x"84",
          3874 => x"0b",
          3875 => x"08",
          3876 => x"82",
          3877 => x"ff",
          3878 => x"55",
          3879 => x"34",
          3880 => x"52",
          3881 => x"fc",
          3882 => x"f6",
          3883 => x"ff",
          3884 => x"06",
          3885 => x"a6",
          3886 => x"d9",
          3887 => x"3d",
          3888 => x"08",
          3889 => x"70",
          3890 => x"52",
          3891 => x"08",
          3892 => x"92",
          3893 => x"84",
          3894 => x"38",
          3895 => x"8f",
          3896 => x"55",
          3897 => x"8b",
          3898 => x"56",
          3899 => x"3f",
          3900 => x"08",
          3901 => x"38",
          3902 => x"f2",
          3903 => x"84",
          3904 => x"58",
          3905 => x"82",
          3906 => x"25",
          3907 => x"93",
          3908 => x"05",
          3909 => x"55",
          3910 => x"74",
          3911 => x"70",
          3912 => x"2a",
          3913 => x"78",
          3914 => x"38",
          3915 => x"38",
          3916 => x"08",
          3917 => x"53",
          3918 => x"aa",
          3919 => x"84",
          3920 => x"88",
          3921 => x"80",
          3922 => x"3f",
          3923 => x"09",
          3924 => x"38",
          3925 => x"51",
          3926 => x"79",
          3927 => x"3f",
          3928 => x"54",
          3929 => x"08",
          3930 => x"58",
          3931 => x"84",
          3932 => x"0d",
          3933 => x"0d",
          3934 => x"5c",
          3935 => x"57",
          3936 => x"73",
          3937 => x"81",
          3938 => x"78",
          3939 => x"56",
          3940 => x"98",
          3941 => x"70",
          3942 => x"33",
          3943 => x"73",
          3944 => x"81",
          3945 => x"75",
          3946 => x"38",
          3947 => x"88",
          3948 => x"d4",
          3949 => x"52",
          3950 => x"3f",
          3951 => x"08",
          3952 => x"74",
          3953 => x"87",
          3954 => x"84",
          3955 => x"38",
          3956 => x"55",
          3957 => x"88",
          3958 => x"2e",
          3959 => x"39",
          3960 => x"ab",
          3961 => x"5a",
          3962 => x"11",
          3963 => x"51",
          3964 => x"82",
          3965 => x"80",
          3966 => x"7a",
          3967 => x"77",
          3968 => x"3f",
          3969 => x"08",
          3970 => x"55",
          3971 => x"74",
          3972 => x"81",
          3973 => x"ff",
          3974 => x"82",
          3975 => x"8e",
          3976 => x"73",
          3977 => x"0c",
          3978 => x"04",
          3979 => x"b0",
          3980 => x"84",
          3981 => x"05",
          3982 => x"80",
          3983 => x"34",
          3984 => x"33",
          3985 => x"cc",
          3986 => x"38",
          3987 => x"33",
          3988 => x"9a",
          3989 => x"eb",
          3990 => x"93",
          3991 => x"8f",
          3992 => x"93",
          3993 => x"2e",
          3994 => x"93",
          3995 => x"f4",
          3996 => x"93",
          3997 => x"bb",
          3998 => x"93",
          3999 => x"2e",
          4000 => x"fd",
          4001 => x"a4",
          4002 => x"39",
          4003 => x"08",
          4004 => x"52",
          4005 => x"52",
          4006 => x"b0",
          4007 => x"84",
          4008 => x"93",
          4009 => x"2e",
          4010 => x"80",
          4011 => x"93",
          4012 => x"d3",
          4013 => x"93",
          4014 => x"80",
          4015 => x"84",
          4016 => x"38",
          4017 => x"08",
          4018 => x"17",
          4019 => x"74",
          4020 => x"74",
          4021 => x"52",
          4022 => x"b4",
          4023 => x"2e",
          4024 => x"ff",
          4025 => x"39",
          4026 => x"8f",
          4027 => x"3d",
          4028 => x"3f",
          4029 => x"08",
          4030 => x"98",
          4031 => x"78",
          4032 => x"38",
          4033 => x"06",
          4034 => x"33",
          4035 => x"70",
          4036 => x"93",
          4037 => x"98",
          4038 => x"2c",
          4039 => x"05",
          4040 => x"81",
          4041 => x"70",
          4042 => x"33",
          4043 => x"51",
          4044 => x"59",
          4045 => x"56",
          4046 => x"80",
          4047 => x"74",
          4048 => x"74",
          4049 => x"29",
          4050 => x"05",
          4051 => x"51",
          4052 => x"24",
          4053 => x"76",
          4054 => x"77",
          4055 => x"3f",
          4056 => x"08",
          4057 => x"54",
          4058 => x"d7",
          4059 => x"93",
          4060 => x"56",
          4061 => x"81",
          4062 => x"81",
          4063 => x"70",
          4064 => x"81",
          4065 => x"51",
          4066 => x"26",
          4067 => x"53",
          4068 => x"51",
          4069 => x"82",
          4070 => x"81",
          4071 => x"73",
          4072 => x"39",
          4073 => x"80",
          4074 => x"38",
          4075 => x"74",
          4076 => x"34",
          4077 => x"70",
          4078 => x"93",
          4079 => x"98",
          4080 => x"2c",
          4081 => x"70",
          4082 => x"fd",
          4083 => x"5e",
          4084 => x"57",
          4085 => x"74",
          4086 => x"81",
          4087 => x"38",
          4088 => x"14",
          4089 => x"80",
          4090 => x"a8",
          4091 => x"82",
          4092 => x"92",
          4093 => x"93",
          4094 => x"82",
          4095 => x"78",
          4096 => x"75",
          4097 => x"54",
          4098 => x"fd",
          4099 => x"84",
          4100 => x"e8",
          4101 => x"08",
          4102 => x"b0",
          4103 => x"7e",
          4104 => x"38",
          4105 => x"33",
          4106 => x"27",
          4107 => x"98",
          4108 => x"2c",
          4109 => x"75",
          4110 => x"74",
          4111 => x"33",
          4112 => x"74",
          4113 => x"29",
          4114 => x"05",
          4115 => x"82",
          4116 => x"56",
          4117 => x"39",
          4118 => x"33",
          4119 => x"54",
          4120 => x"b0",
          4121 => x"54",
          4122 => x"74",
          4123 => x"ac",
          4124 => x"7e",
          4125 => x"81",
          4126 => x"82",
          4127 => x"82",
          4128 => x"70",
          4129 => x"29",
          4130 => x"05",
          4131 => x"82",
          4132 => x"5a",
          4133 => x"74",
          4134 => x"38",
          4135 => x"33",
          4136 => x"c7",
          4137 => x"80",
          4138 => x"80",
          4139 => x"98",
          4140 => x"ac",
          4141 => x"55",
          4142 => x"e0",
          4143 => x"b0",
          4144 => x"2b",
          4145 => x"82",
          4146 => x"5a",
          4147 => x"74",
          4148 => x"9a",
          4149 => x"e8",
          4150 => x"81",
          4151 => x"81",
          4152 => x"70",
          4153 => x"93",
          4154 => x"51",
          4155 => x"24",
          4156 => x"fa",
          4157 => x"b0",
          4158 => x"ff",
          4159 => x"73",
          4160 => x"ea",
          4161 => x"ac",
          4162 => x"54",
          4163 => x"ac",
          4164 => x"54",
          4165 => x"b0",
          4166 => x"e7",
          4167 => x"93",
          4168 => x"98",
          4169 => x"2c",
          4170 => x"33",
          4171 => x"57",
          4172 => x"a7",
          4173 => x"54",
          4174 => x"74",
          4175 => x"51",
          4176 => x"74",
          4177 => x"29",
          4178 => x"05",
          4179 => x"82",
          4180 => x"58",
          4181 => x"75",
          4182 => x"a0",
          4183 => x"3f",
          4184 => x"33",
          4185 => x"70",
          4186 => x"93",
          4187 => x"51",
          4188 => x"74",
          4189 => x"38",
          4190 => x"ef",
          4191 => x"80",
          4192 => x"80",
          4193 => x"98",
          4194 => x"ac",
          4195 => x"55",
          4196 => x"e4",
          4197 => x"39",
          4198 => x"33",
          4199 => x"80",
          4200 => x"51",
          4201 => x"82",
          4202 => x"79",
          4203 => x"3f",
          4204 => x"08",
          4205 => x"54",
          4206 => x"82",
          4207 => x"54",
          4208 => x"84",
          4209 => x"53",
          4210 => x"51",
          4211 => x"84",
          4212 => x"7a",
          4213 => x"39",
          4214 => x"33",
          4215 => x"2e",
          4216 => x"88",
          4217 => x"3f",
          4218 => x"33",
          4219 => x"73",
          4220 => x"34",
          4221 => x"06",
          4222 => x"82",
          4223 => x"82",
          4224 => x"55",
          4225 => x"2e",
          4226 => x"ff",
          4227 => x"82",
          4228 => x"74",
          4229 => x"98",
          4230 => x"ff",
          4231 => x"55",
          4232 => x"a7",
          4233 => x"54",
          4234 => x"74",
          4235 => x"51",
          4236 => x"74",
          4237 => x"29",
          4238 => x"05",
          4239 => x"82",
          4240 => x"58",
          4241 => x"75",
          4242 => x"a0",
          4243 => x"3f",
          4244 => x"33",
          4245 => x"70",
          4246 => x"93",
          4247 => x"51",
          4248 => x"74",
          4249 => x"38",
          4250 => x"ff",
          4251 => x"80",
          4252 => x"80",
          4253 => x"98",
          4254 => x"ac",
          4255 => x"55",
          4256 => x"e4",
          4257 => x"39",
          4258 => x"33",
          4259 => x"06",
          4260 => x"33",
          4261 => x"74",
          4262 => x"d2",
          4263 => x"54",
          4264 => x"b0",
          4265 => x"70",
          4266 => x"e4",
          4267 => x"93",
          4268 => x"81",
          4269 => x"93",
          4270 => x"56",
          4271 => x"26",
          4272 => x"aa",
          4273 => x"38",
          4274 => x"08",
          4275 => x"2e",
          4276 => x"51",
          4277 => x"82",
          4278 => x"82",
          4279 => x"82",
          4280 => x"81",
          4281 => x"05",
          4282 => x"79",
          4283 => x"3f",
          4284 => x"c1",
          4285 => x"29",
          4286 => x"05",
          4287 => x"56",
          4288 => x"2e",
          4289 => x"51",
          4290 => x"82",
          4291 => x"82",
          4292 => x"82",
          4293 => x"81",
          4294 => x"05",
          4295 => x"79",
          4296 => x"3f",
          4297 => x"80",
          4298 => x"08",
          4299 => x"2e",
          4300 => x"74",
          4301 => x"3f",
          4302 => x"7a",
          4303 => x"81",
          4304 => x"82",
          4305 => x"55",
          4306 => x"89",
          4307 => x"ca",
          4308 => x"c8",
          4309 => x"29",
          4310 => x"05",
          4311 => x"56",
          4312 => x"2e",
          4313 => x"51",
          4314 => x"82",
          4315 => x"82",
          4316 => x"82",
          4317 => x"81",
          4318 => x"05",
          4319 => x"79",
          4320 => x"3f",
          4321 => x"73",
          4322 => x"5b",
          4323 => x"08",
          4324 => x"2e",
          4325 => x"74",
          4326 => x"3f",
          4327 => x"08",
          4328 => x"34",
          4329 => x"08",
          4330 => x"81",
          4331 => x"52",
          4332 => x"9f",
          4333 => x"b0",
          4334 => x"ac",
          4335 => x"51",
          4336 => x"f6",
          4337 => x"93",
          4338 => x"81",
          4339 => x"93",
          4340 => x"56",
          4341 => x"27",
          4342 => x"81",
          4343 => x"82",
          4344 => x"74",
          4345 => x"52",
          4346 => x"3f",
          4347 => x"82",
          4348 => x"54",
          4349 => x"f5",
          4350 => x"51",
          4351 => x"82",
          4352 => x"ff",
          4353 => x"82",
          4354 => x"f5",
          4355 => x"0b",
          4356 => x"34",
          4357 => x"93",
          4358 => x"82",
          4359 => x"af",
          4360 => x"ff",
          4361 => x"8f",
          4362 => x"81",
          4363 => x"26",
          4364 => x"8f",
          4365 => x"52",
          4366 => x"84",
          4367 => x"0d",
          4368 => x"0d",
          4369 => x"33",
          4370 => x"9f",
          4371 => x"53",
          4372 => x"81",
          4373 => x"38",
          4374 => x"87",
          4375 => x"11",
          4376 => x"54",
          4377 => x"84",
          4378 => x"54",
          4379 => x"87",
          4380 => x"11",
          4381 => x"0c",
          4382 => x"c0",
          4383 => x"70",
          4384 => x"70",
          4385 => x"51",
          4386 => x"8a",
          4387 => x"98",
          4388 => x"70",
          4389 => x"08",
          4390 => x"06",
          4391 => x"38",
          4392 => x"8c",
          4393 => x"80",
          4394 => x"71",
          4395 => x"14",
          4396 => x"ec",
          4397 => x"70",
          4398 => x"0c",
          4399 => x"04",
          4400 => x"60",
          4401 => x"8c",
          4402 => x"33",
          4403 => x"5b",
          4404 => x"5a",
          4405 => x"82",
          4406 => x"81",
          4407 => x"52",
          4408 => x"38",
          4409 => x"84",
          4410 => x"92",
          4411 => x"c0",
          4412 => x"87",
          4413 => x"13",
          4414 => x"57",
          4415 => x"0b",
          4416 => x"8c",
          4417 => x"0c",
          4418 => x"75",
          4419 => x"2a",
          4420 => x"51",
          4421 => x"80",
          4422 => x"7b",
          4423 => x"7b",
          4424 => x"5d",
          4425 => x"59",
          4426 => x"06",
          4427 => x"73",
          4428 => x"81",
          4429 => x"ff",
          4430 => x"72",
          4431 => x"38",
          4432 => x"8c",
          4433 => x"c3",
          4434 => x"98",
          4435 => x"71",
          4436 => x"38",
          4437 => x"2e",
          4438 => x"76",
          4439 => x"92",
          4440 => x"72",
          4441 => x"06",
          4442 => x"f7",
          4443 => x"5a",
          4444 => x"80",
          4445 => x"70",
          4446 => x"5a",
          4447 => x"80",
          4448 => x"73",
          4449 => x"06",
          4450 => x"38",
          4451 => x"fe",
          4452 => x"fc",
          4453 => x"52",
          4454 => x"83",
          4455 => x"71",
          4456 => x"93",
          4457 => x"3d",
          4458 => x"3d",
          4459 => x"64",
          4460 => x"bf",
          4461 => x"40",
          4462 => x"59",
          4463 => x"58",
          4464 => x"82",
          4465 => x"81",
          4466 => x"52",
          4467 => x"09",
          4468 => x"b1",
          4469 => x"84",
          4470 => x"92",
          4471 => x"c0",
          4472 => x"87",
          4473 => x"13",
          4474 => x"56",
          4475 => x"87",
          4476 => x"0c",
          4477 => x"82",
          4478 => x"58",
          4479 => x"84",
          4480 => x"06",
          4481 => x"71",
          4482 => x"38",
          4483 => x"05",
          4484 => x"0c",
          4485 => x"73",
          4486 => x"81",
          4487 => x"71",
          4488 => x"38",
          4489 => x"8c",
          4490 => x"d0",
          4491 => x"98",
          4492 => x"71",
          4493 => x"38",
          4494 => x"2e",
          4495 => x"76",
          4496 => x"92",
          4497 => x"72",
          4498 => x"06",
          4499 => x"f7",
          4500 => x"59",
          4501 => x"1a",
          4502 => x"06",
          4503 => x"59",
          4504 => x"80",
          4505 => x"73",
          4506 => x"06",
          4507 => x"38",
          4508 => x"fe",
          4509 => x"fc",
          4510 => x"52",
          4511 => x"83",
          4512 => x"71",
          4513 => x"93",
          4514 => x"3d",
          4515 => x"3d",
          4516 => x"84",
          4517 => x"33",
          4518 => x"a7",
          4519 => x"54",
          4520 => x"fa",
          4521 => x"93",
          4522 => x"06",
          4523 => x"72",
          4524 => x"85",
          4525 => x"98",
          4526 => x"56",
          4527 => x"80",
          4528 => x"76",
          4529 => x"74",
          4530 => x"c0",
          4531 => x"54",
          4532 => x"2e",
          4533 => x"d4",
          4534 => x"2e",
          4535 => x"80",
          4536 => x"08",
          4537 => x"70",
          4538 => x"51",
          4539 => x"2e",
          4540 => x"c0",
          4541 => x"52",
          4542 => x"87",
          4543 => x"08",
          4544 => x"38",
          4545 => x"87",
          4546 => x"14",
          4547 => x"70",
          4548 => x"52",
          4549 => x"96",
          4550 => x"92",
          4551 => x"0a",
          4552 => x"39",
          4553 => x"0c",
          4554 => x"39",
          4555 => x"54",
          4556 => x"84",
          4557 => x"0d",
          4558 => x"0d",
          4559 => x"33",
          4560 => x"88",
          4561 => x"93",
          4562 => x"51",
          4563 => x"04",
          4564 => x"75",
          4565 => x"82",
          4566 => x"90",
          4567 => x"2b",
          4568 => x"33",
          4569 => x"88",
          4570 => x"71",
          4571 => x"84",
          4572 => x"54",
          4573 => x"85",
          4574 => x"ff",
          4575 => x"02",
          4576 => x"05",
          4577 => x"70",
          4578 => x"05",
          4579 => x"88",
          4580 => x"72",
          4581 => x"0d",
          4582 => x"0d",
          4583 => x"52",
          4584 => x"81",
          4585 => x"70",
          4586 => x"70",
          4587 => x"05",
          4588 => x"88",
          4589 => x"72",
          4590 => x"54",
          4591 => x"2a",
          4592 => x"34",
          4593 => x"04",
          4594 => x"76",
          4595 => x"54",
          4596 => x"2e",
          4597 => x"70",
          4598 => x"33",
          4599 => x"05",
          4600 => x"11",
          4601 => x"84",
          4602 => x"fe",
          4603 => x"77",
          4604 => x"53",
          4605 => x"81",
          4606 => x"ff",
          4607 => x"f4",
          4608 => x"0d",
          4609 => x"0d",
          4610 => x"56",
          4611 => x"70",
          4612 => x"33",
          4613 => x"05",
          4614 => x"71",
          4615 => x"56",
          4616 => x"72",
          4617 => x"38",
          4618 => x"e2",
          4619 => x"93",
          4620 => x"3d",
          4621 => x"3d",
          4622 => x"54",
          4623 => x"71",
          4624 => x"38",
          4625 => x"70",
          4626 => x"f3",
          4627 => x"82",
          4628 => x"84",
          4629 => x"80",
          4630 => x"84",
          4631 => x"0b",
          4632 => x"0c",
          4633 => x"0d",
          4634 => x"0b",
          4635 => x"56",
          4636 => x"2e",
          4637 => x"81",
          4638 => x"08",
          4639 => x"70",
          4640 => x"33",
          4641 => x"a2",
          4642 => x"84",
          4643 => x"09",
          4644 => x"38",
          4645 => x"08",
          4646 => x"b0",
          4647 => x"a4",
          4648 => x"9c",
          4649 => x"56",
          4650 => x"27",
          4651 => x"16",
          4652 => x"82",
          4653 => x"06",
          4654 => x"54",
          4655 => x"78",
          4656 => x"33",
          4657 => x"3f",
          4658 => x"5a",
          4659 => x"84",
          4660 => x"0d",
          4661 => x"0d",
          4662 => x"56",
          4663 => x"b0",
          4664 => x"af",
          4665 => x"fe",
          4666 => x"93",
          4667 => x"82",
          4668 => x"9f",
          4669 => x"74",
          4670 => x"52",
          4671 => x"51",
          4672 => x"82",
          4673 => x"80",
          4674 => x"ff",
          4675 => x"74",
          4676 => x"76",
          4677 => x"0c",
          4678 => x"04",
          4679 => x"7a",
          4680 => x"fe",
          4681 => x"93",
          4682 => x"82",
          4683 => x"81",
          4684 => x"33",
          4685 => x"2e",
          4686 => x"80",
          4687 => x"17",
          4688 => x"81",
          4689 => x"06",
          4690 => x"84",
          4691 => x"93",
          4692 => x"b4",
          4693 => x"56",
          4694 => x"82",
          4695 => x"84",
          4696 => x"fc",
          4697 => x"8b",
          4698 => x"52",
          4699 => x"a9",
          4700 => x"85",
          4701 => x"84",
          4702 => x"fc",
          4703 => x"17",
          4704 => x"9c",
          4705 => x"91",
          4706 => x"08",
          4707 => x"17",
          4708 => x"3f",
          4709 => x"81",
          4710 => x"19",
          4711 => x"53",
          4712 => x"17",
          4713 => x"82",
          4714 => x"18",
          4715 => x"80",
          4716 => x"33",
          4717 => x"3f",
          4718 => x"08",
          4719 => x"38",
          4720 => x"82",
          4721 => x"8a",
          4722 => x"fb",
          4723 => x"fe",
          4724 => x"08",
          4725 => x"56",
          4726 => x"74",
          4727 => x"38",
          4728 => x"75",
          4729 => x"16",
          4730 => x"53",
          4731 => x"84",
          4732 => x"0d",
          4733 => x"0d",
          4734 => x"08",
          4735 => x"81",
          4736 => x"df",
          4737 => x"15",
          4738 => x"d7",
          4739 => x"33",
          4740 => x"82",
          4741 => x"38",
          4742 => x"89",
          4743 => x"2e",
          4744 => x"bf",
          4745 => x"2e",
          4746 => x"81",
          4747 => x"81",
          4748 => x"89",
          4749 => x"08",
          4750 => x"52",
          4751 => x"3f",
          4752 => x"08",
          4753 => x"74",
          4754 => x"14",
          4755 => x"81",
          4756 => x"2a",
          4757 => x"05",
          4758 => x"57",
          4759 => x"f5",
          4760 => x"84",
          4761 => x"38",
          4762 => x"06",
          4763 => x"33",
          4764 => x"78",
          4765 => x"06",
          4766 => x"5c",
          4767 => x"53",
          4768 => x"38",
          4769 => x"06",
          4770 => x"39",
          4771 => x"a4",
          4772 => x"52",
          4773 => x"bd",
          4774 => x"84",
          4775 => x"38",
          4776 => x"fe",
          4777 => x"b4",
          4778 => x"8d",
          4779 => x"84",
          4780 => x"ff",
          4781 => x"39",
          4782 => x"a4",
          4783 => x"52",
          4784 => x"91",
          4785 => x"84",
          4786 => x"76",
          4787 => x"fc",
          4788 => x"b4",
          4789 => x"f8",
          4790 => x"84",
          4791 => x"06",
          4792 => x"81",
          4793 => x"93",
          4794 => x"3d",
          4795 => x"3d",
          4796 => x"7e",
          4797 => x"82",
          4798 => x"27",
          4799 => x"76",
          4800 => x"27",
          4801 => x"75",
          4802 => x"79",
          4803 => x"38",
          4804 => x"89",
          4805 => x"2e",
          4806 => x"80",
          4807 => x"2e",
          4808 => x"81",
          4809 => x"81",
          4810 => x"89",
          4811 => x"08",
          4812 => x"52",
          4813 => x"3f",
          4814 => x"08",
          4815 => x"84",
          4816 => x"38",
          4817 => x"06",
          4818 => x"81",
          4819 => x"06",
          4820 => x"77",
          4821 => x"2e",
          4822 => x"84",
          4823 => x"06",
          4824 => x"06",
          4825 => x"53",
          4826 => x"81",
          4827 => x"34",
          4828 => x"a4",
          4829 => x"52",
          4830 => x"d9",
          4831 => x"84",
          4832 => x"93",
          4833 => x"94",
          4834 => x"ff",
          4835 => x"05",
          4836 => x"54",
          4837 => x"38",
          4838 => x"74",
          4839 => x"06",
          4840 => x"07",
          4841 => x"74",
          4842 => x"39",
          4843 => x"a4",
          4844 => x"52",
          4845 => x"9d",
          4846 => x"84",
          4847 => x"93",
          4848 => x"d8",
          4849 => x"ff",
          4850 => x"76",
          4851 => x"06",
          4852 => x"05",
          4853 => x"3f",
          4854 => x"87",
          4855 => x"08",
          4856 => x"51",
          4857 => x"82",
          4858 => x"59",
          4859 => x"08",
          4860 => x"f0",
          4861 => x"82",
          4862 => x"06",
          4863 => x"05",
          4864 => x"54",
          4865 => x"3f",
          4866 => x"08",
          4867 => x"74",
          4868 => x"51",
          4869 => x"81",
          4870 => x"34",
          4871 => x"84",
          4872 => x"0d",
          4873 => x"0d",
          4874 => x"72",
          4875 => x"56",
          4876 => x"27",
          4877 => x"98",
          4878 => x"9d",
          4879 => x"2e",
          4880 => x"53",
          4881 => x"51",
          4882 => x"82",
          4883 => x"54",
          4884 => x"08",
          4885 => x"93",
          4886 => x"80",
          4887 => x"54",
          4888 => x"82",
          4889 => x"54",
          4890 => x"74",
          4891 => x"fb",
          4892 => x"93",
          4893 => x"82",
          4894 => x"80",
          4895 => x"38",
          4896 => x"08",
          4897 => x"38",
          4898 => x"08",
          4899 => x"38",
          4900 => x"52",
          4901 => x"d6",
          4902 => x"84",
          4903 => x"98",
          4904 => x"11",
          4905 => x"57",
          4906 => x"74",
          4907 => x"81",
          4908 => x"0c",
          4909 => x"81",
          4910 => x"84",
          4911 => x"55",
          4912 => x"ff",
          4913 => x"54",
          4914 => x"84",
          4915 => x"0d",
          4916 => x"0d",
          4917 => x"08",
          4918 => x"79",
          4919 => x"17",
          4920 => x"80",
          4921 => x"98",
          4922 => x"26",
          4923 => x"58",
          4924 => x"52",
          4925 => x"fd",
          4926 => x"74",
          4927 => x"08",
          4928 => x"38",
          4929 => x"08",
          4930 => x"84",
          4931 => x"82",
          4932 => x"17",
          4933 => x"84",
          4934 => x"c7",
          4935 => x"90",
          4936 => x"56",
          4937 => x"2e",
          4938 => x"77",
          4939 => x"81",
          4940 => x"38",
          4941 => x"98",
          4942 => x"26",
          4943 => x"56",
          4944 => x"51",
          4945 => x"80",
          4946 => x"84",
          4947 => x"09",
          4948 => x"38",
          4949 => x"08",
          4950 => x"84",
          4951 => x"30",
          4952 => x"80",
          4953 => x"07",
          4954 => x"08",
          4955 => x"55",
          4956 => x"ef",
          4957 => x"84",
          4958 => x"95",
          4959 => x"08",
          4960 => x"27",
          4961 => x"98",
          4962 => x"89",
          4963 => x"85",
          4964 => x"db",
          4965 => x"81",
          4966 => x"17",
          4967 => x"89",
          4968 => x"75",
          4969 => x"ac",
          4970 => x"7a",
          4971 => x"3f",
          4972 => x"08",
          4973 => x"38",
          4974 => x"93",
          4975 => x"2e",
          4976 => x"86",
          4977 => x"84",
          4978 => x"93",
          4979 => x"70",
          4980 => x"07",
          4981 => x"7c",
          4982 => x"55",
          4983 => x"f8",
          4984 => x"2e",
          4985 => x"ff",
          4986 => x"55",
          4987 => x"ff",
          4988 => x"76",
          4989 => x"3f",
          4990 => x"08",
          4991 => x"08",
          4992 => x"93",
          4993 => x"80",
          4994 => x"55",
          4995 => x"94",
          4996 => x"2e",
          4997 => x"53",
          4998 => x"51",
          4999 => x"82",
          5000 => x"55",
          5001 => x"75",
          5002 => x"98",
          5003 => x"05",
          5004 => x"56",
          5005 => x"26",
          5006 => x"15",
          5007 => x"84",
          5008 => x"07",
          5009 => x"18",
          5010 => x"ff",
          5011 => x"2e",
          5012 => x"39",
          5013 => x"39",
          5014 => x"08",
          5015 => x"81",
          5016 => x"74",
          5017 => x"0c",
          5018 => x"04",
          5019 => x"7a",
          5020 => x"f3",
          5021 => x"93",
          5022 => x"81",
          5023 => x"84",
          5024 => x"38",
          5025 => x"51",
          5026 => x"82",
          5027 => x"82",
          5028 => x"b0",
          5029 => x"84",
          5030 => x"52",
          5031 => x"52",
          5032 => x"3f",
          5033 => x"39",
          5034 => x"8a",
          5035 => x"75",
          5036 => x"38",
          5037 => x"19",
          5038 => x"81",
          5039 => x"ed",
          5040 => x"93",
          5041 => x"2e",
          5042 => x"15",
          5043 => x"70",
          5044 => x"07",
          5045 => x"53",
          5046 => x"75",
          5047 => x"0c",
          5048 => x"04",
          5049 => x"7a",
          5050 => x"58",
          5051 => x"f0",
          5052 => x"80",
          5053 => x"9f",
          5054 => x"80",
          5055 => x"90",
          5056 => x"17",
          5057 => x"aa",
          5058 => x"53",
          5059 => x"88",
          5060 => x"08",
          5061 => x"38",
          5062 => x"53",
          5063 => x"17",
          5064 => x"72",
          5065 => x"fe",
          5066 => x"08",
          5067 => x"80",
          5068 => x"16",
          5069 => x"2b",
          5070 => x"75",
          5071 => x"73",
          5072 => x"f5",
          5073 => x"93",
          5074 => x"82",
          5075 => x"ff",
          5076 => x"81",
          5077 => x"84",
          5078 => x"38",
          5079 => x"82",
          5080 => x"26",
          5081 => x"58",
          5082 => x"73",
          5083 => x"39",
          5084 => x"51",
          5085 => x"82",
          5086 => x"98",
          5087 => x"94",
          5088 => x"17",
          5089 => x"58",
          5090 => x"9a",
          5091 => x"81",
          5092 => x"74",
          5093 => x"98",
          5094 => x"83",
          5095 => x"b4",
          5096 => x"0c",
          5097 => x"82",
          5098 => x"8a",
          5099 => x"f8",
          5100 => x"70",
          5101 => x"08",
          5102 => x"57",
          5103 => x"0a",
          5104 => x"38",
          5105 => x"15",
          5106 => x"08",
          5107 => x"72",
          5108 => x"cb",
          5109 => x"ff",
          5110 => x"81",
          5111 => x"13",
          5112 => x"94",
          5113 => x"74",
          5114 => x"85",
          5115 => x"22",
          5116 => x"73",
          5117 => x"38",
          5118 => x"8a",
          5119 => x"05",
          5120 => x"06",
          5121 => x"8a",
          5122 => x"73",
          5123 => x"3f",
          5124 => x"08",
          5125 => x"81",
          5126 => x"84",
          5127 => x"ff",
          5128 => x"82",
          5129 => x"ff",
          5130 => x"38",
          5131 => x"82",
          5132 => x"26",
          5133 => x"7b",
          5134 => x"98",
          5135 => x"55",
          5136 => x"94",
          5137 => x"73",
          5138 => x"3f",
          5139 => x"08",
          5140 => x"82",
          5141 => x"80",
          5142 => x"38",
          5143 => x"93",
          5144 => x"2e",
          5145 => x"55",
          5146 => x"08",
          5147 => x"38",
          5148 => x"08",
          5149 => x"fb",
          5150 => x"93",
          5151 => x"38",
          5152 => x"0c",
          5153 => x"51",
          5154 => x"82",
          5155 => x"98",
          5156 => x"90",
          5157 => x"16",
          5158 => x"15",
          5159 => x"74",
          5160 => x"0c",
          5161 => x"04",
          5162 => x"7b",
          5163 => x"5b",
          5164 => x"52",
          5165 => x"ac",
          5166 => x"84",
          5167 => x"93",
          5168 => x"ec",
          5169 => x"84",
          5170 => x"17",
          5171 => x"51",
          5172 => x"82",
          5173 => x"54",
          5174 => x"08",
          5175 => x"82",
          5176 => x"9c",
          5177 => x"33",
          5178 => x"72",
          5179 => x"09",
          5180 => x"38",
          5181 => x"93",
          5182 => x"72",
          5183 => x"55",
          5184 => x"53",
          5185 => x"8e",
          5186 => x"56",
          5187 => x"09",
          5188 => x"38",
          5189 => x"93",
          5190 => x"81",
          5191 => x"fd",
          5192 => x"93",
          5193 => x"82",
          5194 => x"80",
          5195 => x"38",
          5196 => x"09",
          5197 => x"38",
          5198 => x"82",
          5199 => x"8b",
          5200 => x"fd",
          5201 => x"9a",
          5202 => x"eb",
          5203 => x"93",
          5204 => x"ff",
          5205 => x"70",
          5206 => x"53",
          5207 => x"09",
          5208 => x"38",
          5209 => x"eb",
          5210 => x"93",
          5211 => x"2b",
          5212 => x"72",
          5213 => x"0c",
          5214 => x"04",
          5215 => x"77",
          5216 => x"ff",
          5217 => x"9a",
          5218 => x"55",
          5219 => x"76",
          5220 => x"53",
          5221 => x"09",
          5222 => x"38",
          5223 => x"52",
          5224 => x"eb",
          5225 => x"3d",
          5226 => x"3d",
          5227 => x"5b",
          5228 => x"08",
          5229 => x"15",
          5230 => x"81",
          5231 => x"15",
          5232 => x"51",
          5233 => x"82",
          5234 => x"58",
          5235 => x"08",
          5236 => x"9c",
          5237 => x"33",
          5238 => x"86",
          5239 => x"80",
          5240 => x"13",
          5241 => x"06",
          5242 => x"06",
          5243 => x"72",
          5244 => x"82",
          5245 => x"53",
          5246 => x"2e",
          5247 => x"53",
          5248 => x"a9",
          5249 => x"74",
          5250 => x"72",
          5251 => x"38",
          5252 => x"99",
          5253 => x"84",
          5254 => x"06",
          5255 => x"88",
          5256 => x"06",
          5257 => x"54",
          5258 => x"a0",
          5259 => x"74",
          5260 => x"3f",
          5261 => x"08",
          5262 => x"84",
          5263 => x"98",
          5264 => x"fa",
          5265 => x"80",
          5266 => x"0c",
          5267 => x"84",
          5268 => x"0d",
          5269 => x"0d",
          5270 => x"57",
          5271 => x"73",
          5272 => x"3f",
          5273 => x"08",
          5274 => x"84",
          5275 => x"98",
          5276 => x"75",
          5277 => x"3f",
          5278 => x"08",
          5279 => x"84",
          5280 => x"a0",
          5281 => x"84",
          5282 => x"14",
          5283 => x"db",
          5284 => x"a0",
          5285 => x"14",
          5286 => x"ac",
          5287 => x"83",
          5288 => x"82",
          5289 => x"87",
          5290 => x"fd",
          5291 => x"70",
          5292 => x"08",
          5293 => x"55",
          5294 => x"3f",
          5295 => x"08",
          5296 => x"13",
          5297 => x"73",
          5298 => x"83",
          5299 => x"3d",
          5300 => x"3d",
          5301 => x"57",
          5302 => x"89",
          5303 => x"17",
          5304 => x"81",
          5305 => x"70",
          5306 => x"55",
          5307 => x"08",
          5308 => x"81",
          5309 => x"52",
          5310 => x"a8",
          5311 => x"2e",
          5312 => x"84",
          5313 => x"52",
          5314 => x"09",
          5315 => x"38",
          5316 => x"81",
          5317 => x"81",
          5318 => x"73",
          5319 => x"55",
          5320 => x"55",
          5321 => x"c5",
          5322 => x"88",
          5323 => x"0b",
          5324 => x"9c",
          5325 => x"8b",
          5326 => x"17",
          5327 => x"08",
          5328 => x"52",
          5329 => x"82",
          5330 => x"76",
          5331 => x"51",
          5332 => x"82",
          5333 => x"86",
          5334 => x"12",
          5335 => x"3f",
          5336 => x"08",
          5337 => x"88",
          5338 => x"f3",
          5339 => x"70",
          5340 => x"80",
          5341 => x"51",
          5342 => x"af",
          5343 => x"81",
          5344 => x"dc",
          5345 => x"74",
          5346 => x"38",
          5347 => x"88",
          5348 => x"39",
          5349 => x"80",
          5350 => x"56",
          5351 => x"af",
          5352 => x"06",
          5353 => x"56",
          5354 => x"32",
          5355 => x"80",
          5356 => x"51",
          5357 => x"dc",
          5358 => x"1c",
          5359 => x"33",
          5360 => x"9f",
          5361 => x"ff",
          5362 => x"1c",
          5363 => x"7a",
          5364 => x"3f",
          5365 => x"08",
          5366 => x"39",
          5367 => x"a0",
          5368 => x"5e",
          5369 => x"52",
          5370 => x"ff",
          5371 => x"59",
          5372 => x"33",
          5373 => x"ae",
          5374 => x"06",
          5375 => x"78",
          5376 => x"81",
          5377 => x"32",
          5378 => x"9f",
          5379 => x"26",
          5380 => x"53",
          5381 => x"73",
          5382 => x"17",
          5383 => x"34",
          5384 => x"db",
          5385 => x"32",
          5386 => x"9f",
          5387 => x"54",
          5388 => x"2e",
          5389 => x"80",
          5390 => x"75",
          5391 => x"bd",
          5392 => x"7e",
          5393 => x"a0",
          5394 => x"bd",
          5395 => x"82",
          5396 => x"18",
          5397 => x"1a",
          5398 => x"a0",
          5399 => x"fc",
          5400 => x"32",
          5401 => x"80",
          5402 => x"30",
          5403 => x"71",
          5404 => x"51",
          5405 => x"55",
          5406 => x"ac",
          5407 => x"81",
          5408 => x"78",
          5409 => x"51",
          5410 => x"af",
          5411 => x"06",
          5412 => x"55",
          5413 => x"32",
          5414 => x"80",
          5415 => x"51",
          5416 => x"db",
          5417 => x"39",
          5418 => x"09",
          5419 => x"38",
          5420 => x"7c",
          5421 => x"54",
          5422 => x"a2",
          5423 => x"32",
          5424 => x"ae",
          5425 => x"72",
          5426 => x"9f",
          5427 => x"51",
          5428 => x"74",
          5429 => x"88",
          5430 => x"fe",
          5431 => x"98",
          5432 => x"80",
          5433 => x"75",
          5434 => x"81",
          5435 => x"33",
          5436 => x"51",
          5437 => x"82",
          5438 => x"80",
          5439 => x"78",
          5440 => x"81",
          5441 => x"5a",
          5442 => x"d2",
          5443 => x"84",
          5444 => x"80",
          5445 => x"1c",
          5446 => x"27",
          5447 => x"79",
          5448 => x"74",
          5449 => x"7a",
          5450 => x"74",
          5451 => x"39",
          5452 => x"ff",
          5453 => x"fe",
          5454 => x"84",
          5455 => x"ff",
          5456 => x"73",
          5457 => x"38",
          5458 => x"81",
          5459 => x"54",
          5460 => x"75",
          5461 => x"17",
          5462 => x"39",
          5463 => x"0c",
          5464 => x"99",
          5465 => x"54",
          5466 => x"2e",
          5467 => x"84",
          5468 => x"34",
          5469 => x"76",
          5470 => x"8b",
          5471 => x"81",
          5472 => x"56",
          5473 => x"80",
          5474 => x"1b",
          5475 => x"08",
          5476 => x"51",
          5477 => x"82",
          5478 => x"56",
          5479 => x"08",
          5480 => x"98",
          5481 => x"76",
          5482 => x"3f",
          5483 => x"08",
          5484 => x"84",
          5485 => x"38",
          5486 => x"70",
          5487 => x"73",
          5488 => x"be",
          5489 => x"33",
          5490 => x"73",
          5491 => x"8b",
          5492 => x"83",
          5493 => x"06",
          5494 => x"73",
          5495 => x"53",
          5496 => x"51",
          5497 => x"82",
          5498 => x"80",
          5499 => x"75",
          5500 => x"f3",
          5501 => x"9f",
          5502 => x"1c",
          5503 => x"74",
          5504 => x"38",
          5505 => x"09",
          5506 => x"e7",
          5507 => x"2a",
          5508 => x"77",
          5509 => x"51",
          5510 => x"2e",
          5511 => x"81",
          5512 => x"80",
          5513 => x"38",
          5514 => x"ab",
          5515 => x"55",
          5516 => x"75",
          5517 => x"73",
          5518 => x"55",
          5519 => x"82",
          5520 => x"06",
          5521 => x"ab",
          5522 => x"33",
          5523 => x"70",
          5524 => x"55",
          5525 => x"2e",
          5526 => x"1b",
          5527 => x"06",
          5528 => x"52",
          5529 => x"db",
          5530 => x"84",
          5531 => x"0c",
          5532 => x"74",
          5533 => x"0c",
          5534 => x"04",
          5535 => x"7c",
          5536 => x"08",
          5537 => x"55",
          5538 => x"59",
          5539 => x"81",
          5540 => x"70",
          5541 => x"33",
          5542 => x"52",
          5543 => x"2e",
          5544 => x"ee",
          5545 => x"2e",
          5546 => x"81",
          5547 => x"33",
          5548 => x"81",
          5549 => x"52",
          5550 => x"26",
          5551 => x"14",
          5552 => x"06",
          5553 => x"52",
          5554 => x"80",
          5555 => x"0b",
          5556 => x"59",
          5557 => x"7a",
          5558 => x"70",
          5559 => x"33",
          5560 => x"05",
          5561 => x"9f",
          5562 => x"53",
          5563 => x"89",
          5564 => x"70",
          5565 => x"54",
          5566 => x"12",
          5567 => x"26",
          5568 => x"12",
          5569 => x"06",
          5570 => x"30",
          5571 => x"51",
          5572 => x"2e",
          5573 => x"85",
          5574 => x"be",
          5575 => x"74",
          5576 => x"30",
          5577 => x"9f",
          5578 => x"2a",
          5579 => x"54",
          5580 => x"2e",
          5581 => x"15",
          5582 => x"55",
          5583 => x"ff",
          5584 => x"39",
          5585 => x"86",
          5586 => x"7c",
          5587 => x"51",
          5588 => x"93",
          5589 => x"70",
          5590 => x"0c",
          5591 => x"04",
          5592 => x"78",
          5593 => x"83",
          5594 => x"0b",
          5595 => x"79",
          5596 => x"e2",
          5597 => x"55",
          5598 => x"08",
          5599 => x"84",
          5600 => x"df",
          5601 => x"93",
          5602 => x"ff",
          5603 => x"83",
          5604 => x"d4",
          5605 => x"81",
          5606 => x"38",
          5607 => x"17",
          5608 => x"74",
          5609 => x"09",
          5610 => x"38",
          5611 => x"81",
          5612 => x"30",
          5613 => x"79",
          5614 => x"54",
          5615 => x"74",
          5616 => x"09",
          5617 => x"38",
          5618 => x"ff",
          5619 => x"ea",
          5620 => x"b1",
          5621 => x"84",
          5622 => x"93",
          5623 => x"2e",
          5624 => x"53",
          5625 => x"52",
          5626 => x"51",
          5627 => x"82",
          5628 => x"55",
          5629 => x"08",
          5630 => x"38",
          5631 => x"82",
          5632 => x"88",
          5633 => x"f2",
          5634 => x"02",
          5635 => x"cb",
          5636 => x"55",
          5637 => x"60",
          5638 => x"3f",
          5639 => x"08",
          5640 => x"80",
          5641 => x"84",
          5642 => x"fc",
          5643 => x"84",
          5644 => x"82",
          5645 => x"70",
          5646 => x"8c",
          5647 => x"2e",
          5648 => x"73",
          5649 => x"81",
          5650 => x"33",
          5651 => x"80",
          5652 => x"81",
          5653 => x"d7",
          5654 => x"93",
          5655 => x"ff",
          5656 => x"06",
          5657 => x"98",
          5658 => x"2e",
          5659 => x"74",
          5660 => x"81",
          5661 => x"8a",
          5662 => x"ac",
          5663 => x"39",
          5664 => x"77",
          5665 => x"81",
          5666 => x"33",
          5667 => x"3f",
          5668 => x"08",
          5669 => x"70",
          5670 => x"55",
          5671 => x"86",
          5672 => x"80",
          5673 => x"74",
          5674 => x"81",
          5675 => x"8a",
          5676 => x"f4",
          5677 => x"53",
          5678 => x"fd",
          5679 => x"93",
          5680 => x"ff",
          5681 => x"82",
          5682 => x"06",
          5683 => x"8c",
          5684 => x"58",
          5685 => x"f6",
          5686 => x"58",
          5687 => x"2e",
          5688 => x"fa",
          5689 => x"e8",
          5690 => x"84",
          5691 => x"78",
          5692 => x"5a",
          5693 => x"90",
          5694 => x"75",
          5695 => x"38",
          5696 => x"3d",
          5697 => x"70",
          5698 => x"08",
          5699 => x"7a",
          5700 => x"38",
          5701 => x"51",
          5702 => x"82",
          5703 => x"81",
          5704 => x"81",
          5705 => x"38",
          5706 => x"83",
          5707 => x"38",
          5708 => x"84",
          5709 => x"38",
          5710 => x"81",
          5711 => x"38",
          5712 => x"db",
          5713 => x"93",
          5714 => x"ff",
          5715 => x"72",
          5716 => x"09",
          5717 => x"d0",
          5718 => x"14",
          5719 => x"3f",
          5720 => x"08",
          5721 => x"06",
          5722 => x"38",
          5723 => x"51",
          5724 => x"82",
          5725 => x"58",
          5726 => x"0c",
          5727 => x"33",
          5728 => x"80",
          5729 => x"ff",
          5730 => x"ff",
          5731 => x"55",
          5732 => x"81",
          5733 => x"38",
          5734 => x"06",
          5735 => x"80",
          5736 => x"52",
          5737 => x"8a",
          5738 => x"80",
          5739 => x"ff",
          5740 => x"53",
          5741 => x"86",
          5742 => x"83",
          5743 => x"c5",
          5744 => x"f5",
          5745 => x"84",
          5746 => x"93",
          5747 => x"15",
          5748 => x"06",
          5749 => x"76",
          5750 => x"80",
          5751 => x"da",
          5752 => x"93",
          5753 => x"ff",
          5754 => x"74",
          5755 => x"d4",
          5756 => x"dc",
          5757 => x"84",
          5758 => x"c2",
          5759 => x"b9",
          5760 => x"84",
          5761 => x"ff",
          5762 => x"56",
          5763 => x"83",
          5764 => x"14",
          5765 => x"71",
          5766 => x"5a",
          5767 => x"26",
          5768 => x"8a",
          5769 => x"74",
          5770 => x"ff",
          5771 => x"82",
          5772 => x"55",
          5773 => x"08",
          5774 => x"ec",
          5775 => x"84",
          5776 => x"ff",
          5777 => x"83",
          5778 => x"74",
          5779 => x"26",
          5780 => x"57",
          5781 => x"26",
          5782 => x"57",
          5783 => x"56",
          5784 => x"82",
          5785 => x"15",
          5786 => x"0c",
          5787 => x"0c",
          5788 => x"a4",
          5789 => x"1d",
          5790 => x"54",
          5791 => x"2e",
          5792 => x"af",
          5793 => x"14",
          5794 => x"3f",
          5795 => x"08",
          5796 => x"06",
          5797 => x"72",
          5798 => x"79",
          5799 => x"80",
          5800 => x"d9",
          5801 => x"93",
          5802 => x"15",
          5803 => x"2b",
          5804 => x"8d",
          5805 => x"2e",
          5806 => x"77",
          5807 => x"0c",
          5808 => x"76",
          5809 => x"38",
          5810 => x"70",
          5811 => x"81",
          5812 => x"53",
          5813 => x"89",
          5814 => x"56",
          5815 => x"08",
          5816 => x"38",
          5817 => x"15",
          5818 => x"8c",
          5819 => x"80",
          5820 => x"34",
          5821 => x"09",
          5822 => x"92",
          5823 => x"14",
          5824 => x"3f",
          5825 => x"08",
          5826 => x"06",
          5827 => x"2e",
          5828 => x"80",
          5829 => x"1b",
          5830 => x"db",
          5831 => x"93",
          5832 => x"ea",
          5833 => x"84",
          5834 => x"34",
          5835 => x"51",
          5836 => x"82",
          5837 => x"83",
          5838 => x"53",
          5839 => x"d5",
          5840 => x"06",
          5841 => x"b4",
          5842 => x"84",
          5843 => x"84",
          5844 => x"85",
          5845 => x"09",
          5846 => x"38",
          5847 => x"51",
          5848 => x"82",
          5849 => x"86",
          5850 => x"f2",
          5851 => x"06",
          5852 => x"9c",
          5853 => x"d8",
          5854 => x"84",
          5855 => x"0c",
          5856 => x"51",
          5857 => x"82",
          5858 => x"8c",
          5859 => x"74",
          5860 => x"c4",
          5861 => x"53",
          5862 => x"c4",
          5863 => x"15",
          5864 => x"94",
          5865 => x"56",
          5866 => x"84",
          5867 => x"0d",
          5868 => x"0d",
          5869 => x"55",
          5870 => x"b9",
          5871 => x"53",
          5872 => x"b1",
          5873 => x"52",
          5874 => x"a9",
          5875 => x"22",
          5876 => x"57",
          5877 => x"2e",
          5878 => x"99",
          5879 => x"33",
          5880 => x"3f",
          5881 => x"08",
          5882 => x"71",
          5883 => x"74",
          5884 => x"83",
          5885 => x"78",
          5886 => x"52",
          5887 => x"84",
          5888 => x"0d",
          5889 => x"0d",
          5890 => x"33",
          5891 => x"3d",
          5892 => x"56",
          5893 => x"8b",
          5894 => x"82",
          5895 => x"24",
          5896 => x"93",
          5897 => x"29",
          5898 => x"05",
          5899 => x"55",
          5900 => x"84",
          5901 => x"34",
          5902 => x"80",
          5903 => x"80",
          5904 => x"75",
          5905 => x"75",
          5906 => x"38",
          5907 => x"3d",
          5908 => x"05",
          5909 => x"3f",
          5910 => x"08",
          5911 => x"93",
          5912 => x"3d",
          5913 => x"3d",
          5914 => x"84",
          5915 => x"05",
          5916 => x"89",
          5917 => x"2e",
          5918 => x"77",
          5919 => x"54",
          5920 => x"05",
          5921 => x"84",
          5922 => x"f6",
          5923 => x"93",
          5924 => x"82",
          5925 => x"84",
          5926 => x"5c",
          5927 => x"3d",
          5928 => x"ed",
          5929 => x"93",
          5930 => x"82",
          5931 => x"92",
          5932 => x"d7",
          5933 => x"98",
          5934 => x"73",
          5935 => x"38",
          5936 => x"9c",
          5937 => x"80",
          5938 => x"38",
          5939 => x"95",
          5940 => x"2e",
          5941 => x"aa",
          5942 => x"ea",
          5943 => x"93",
          5944 => x"9e",
          5945 => x"05",
          5946 => x"54",
          5947 => x"38",
          5948 => x"70",
          5949 => x"54",
          5950 => x"8e",
          5951 => x"83",
          5952 => x"88",
          5953 => x"83",
          5954 => x"83",
          5955 => x"06",
          5956 => x"80",
          5957 => x"38",
          5958 => x"51",
          5959 => x"82",
          5960 => x"56",
          5961 => x"0a",
          5962 => x"05",
          5963 => x"3f",
          5964 => x"0b",
          5965 => x"80",
          5966 => x"7a",
          5967 => x"3f",
          5968 => x"9c",
          5969 => x"d1",
          5970 => x"81",
          5971 => x"34",
          5972 => x"80",
          5973 => x"b0",
          5974 => x"54",
          5975 => x"52",
          5976 => x"05",
          5977 => x"3f",
          5978 => x"08",
          5979 => x"84",
          5980 => x"38",
          5981 => x"82",
          5982 => x"b2",
          5983 => x"84",
          5984 => x"06",
          5985 => x"73",
          5986 => x"38",
          5987 => x"ad",
          5988 => x"2a",
          5989 => x"51",
          5990 => x"2e",
          5991 => x"81",
          5992 => x"80",
          5993 => x"87",
          5994 => x"39",
          5995 => x"51",
          5996 => x"82",
          5997 => x"7b",
          5998 => x"12",
          5999 => x"82",
          6000 => x"81",
          6001 => x"83",
          6002 => x"06",
          6003 => x"80",
          6004 => x"77",
          6005 => x"58",
          6006 => x"08",
          6007 => x"63",
          6008 => x"63",
          6009 => x"57",
          6010 => x"82",
          6011 => x"82",
          6012 => x"88",
          6013 => x"9c",
          6014 => x"d2",
          6015 => x"93",
          6016 => x"93",
          6017 => x"1b",
          6018 => x"0c",
          6019 => x"22",
          6020 => x"77",
          6021 => x"80",
          6022 => x"34",
          6023 => x"1a",
          6024 => x"94",
          6025 => x"85",
          6026 => x"06",
          6027 => x"80",
          6028 => x"38",
          6029 => x"08",
          6030 => x"84",
          6031 => x"84",
          6032 => x"0c",
          6033 => x"70",
          6034 => x"52",
          6035 => x"39",
          6036 => x"51",
          6037 => x"82",
          6038 => x"57",
          6039 => x"08",
          6040 => x"38",
          6041 => x"93",
          6042 => x"2e",
          6043 => x"83",
          6044 => x"75",
          6045 => x"74",
          6046 => x"07",
          6047 => x"54",
          6048 => x"8a",
          6049 => x"75",
          6050 => x"73",
          6051 => x"98",
          6052 => x"a9",
          6053 => x"ff",
          6054 => x"80",
          6055 => x"76",
          6056 => x"d6",
          6057 => x"93",
          6058 => x"38",
          6059 => x"39",
          6060 => x"82",
          6061 => x"05",
          6062 => x"84",
          6063 => x"0c",
          6064 => x"82",
          6065 => x"97",
          6066 => x"f2",
          6067 => x"63",
          6068 => x"40",
          6069 => x"7e",
          6070 => x"fc",
          6071 => x"51",
          6072 => x"82",
          6073 => x"55",
          6074 => x"08",
          6075 => x"19",
          6076 => x"80",
          6077 => x"74",
          6078 => x"39",
          6079 => x"81",
          6080 => x"56",
          6081 => x"82",
          6082 => x"39",
          6083 => x"1a",
          6084 => x"82",
          6085 => x"0b",
          6086 => x"81",
          6087 => x"39",
          6088 => x"94",
          6089 => x"55",
          6090 => x"83",
          6091 => x"7b",
          6092 => x"89",
          6093 => x"08",
          6094 => x"06",
          6095 => x"81",
          6096 => x"8a",
          6097 => x"05",
          6098 => x"06",
          6099 => x"a8",
          6100 => x"38",
          6101 => x"55",
          6102 => x"19",
          6103 => x"51",
          6104 => x"82",
          6105 => x"55",
          6106 => x"ff",
          6107 => x"ff",
          6108 => x"38",
          6109 => x"0c",
          6110 => x"52",
          6111 => x"cb",
          6112 => x"84",
          6113 => x"ff",
          6114 => x"93",
          6115 => x"7c",
          6116 => x"57",
          6117 => x"80",
          6118 => x"1a",
          6119 => x"22",
          6120 => x"75",
          6121 => x"38",
          6122 => x"58",
          6123 => x"53",
          6124 => x"1b",
          6125 => x"88",
          6126 => x"84",
          6127 => x"38",
          6128 => x"33",
          6129 => x"80",
          6130 => x"b0",
          6131 => x"31",
          6132 => x"27",
          6133 => x"80",
          6134 => x"52",
          6135 => x"77",
          6136 => x"7d",
          6137 => x"e0",
          6138 => x"2b",
          6139 => x"76",
          6140 => x"94",
          6141 => x"ff",
          6142 => x"71",
          6143 => x"7b",
          6144 => x"38",
          6145 => x"19",
          6146 => x"51",
          6147 => x"82",
          6148 => x"fe",
          6149 => x"53",
          6150 => x"83",
          6151 => x"b4",
          6152 => x"51",
          6153 => x"7b",
          6154 => x"08",
          6155 => x"76",
          6156 => x"08",
          6157 => x"0c",
          6158 => x"f3",
          6159 => x"75",
          6160 => x"0c",
          6161 => x"04",
          6162 => x"60",
          6163 => x"40",
          6164 => x"80",
          6165 => x"3d",
          6166 => x"77",
          6167 => x"3f",
          6168 => x"08",
          6169 => x"84",
          6170 => x"91",
          6171 => x"74",
          6172 => x"38",
          6173 => x"b8",
          6174 => x"33",
          6175 => x"70",
          6176 => x"56",
          6177 => x"74",
          6178 => x"a4",
          6179 => x"82",
          6180 => x"34",
          6181 => x"98",
          6182 => x"91",
          6183 => x"56",
          6184 => x"94",
          6185 => x"11",
          6186 => x"76",
          6187 => x"75",
          6188 => x"80",
          6189 => x"38",
          6190 => x"70",
          6191 => x"56",
          6192 => x"fd",
          6193 => x"11",
          6194 => x"77",
          6195 => x"5c",
          6196 => x"38",
          6197 => x"88",
          6198 => x"74",
          6199 => x"52",
          6200 => x"18",
          6201 => x"51",
          6202 => x"82",
          6203 => x"55",
          6204 => x"08",
          6205 => x"ab",
          6206 => x"2e",
          6207 => x"74",
          6208 => x"95",
          6209 => x"19",
          6210 => x"08",
          6211 => x"88",
          6212 => x"55",
          6213 => x"9c",
          6214 => x"09",
          6215 => x"38",
          6216 => x"c1",
          6217 => x"84",
          6218 => x"38",
          6219 => x"52",
          6220 => x"97",
          6221 => x"84",
          6222 => x"fe",
          6223 => x"93",
          6224 => x"7c",
          6225 => x"57",
          6226 => x"80",
          6227 => x"1b",
          6228 => x"22",
          6229 => x"75",
          6230 => x"38",
          6231 => x"59",
          6232 => x"53",
          6233 => x"1a",
          6234 => x"be",
          6235 => x"84",
          6236 => x"38",
          6237 => x"08",
          6238 => x"56",
          6239 => x"9b",
          6240 => x"53",
          6241 => x"77",
          6242 => x"7d",
          6243 => x"16",
          6244 => x"3f",
          6245 => x"0b",
          6246 => x"78",
          6247 => x"80",
          6248 => x"18",
          6249 => x"08",
          6250 => x"7e",
          6251 => x"3f",
          6252 => x"08",
          6253 => x"7e",
          6254 => x"0c",
          6255 => x"19",
          6256 => x"08",
          6257 => x"84",
          6258 => x"57",
          6259 => x"27",
          6260 => x"56",
          6261 => x"52",
          6262 => x"f9",
          6263 => x"84",
          6264 => x"38",
          6265 => x"52",
          6266 => x"83",
          6267 => x"b4",
          6268 => x"d4",
          6269 => x"81",
          6270 => x"34",
          6271 => x"7e",
          6272 => x"0c",
          6273 => x"1a",
          6274 => x"94",
          6275 => x"1b",
          6276 => x"5e",
          6277 => x"27",
          6278 => x"55",
          6279 => x"0c",
          6280 => x"90",
          6281 => x"c0",
          6282 => x"90",
          6283 => x"56",
          6284 => x"84",
          6285 => x"0d",
          6286 => x"0d",
          6287 => x"fc",
          6288 => x"52",
          6289 => x"3f",
          6290 => x"08",
          6291 => x"84",
          6292 => x"38",
          6293 => x"70",
          6294 => x"81",
          6295 => x"55",
          6296 => x"80",
          6297 => x"16",
          6298 => x"51",
          6299 => x"82",
          6300 => x"57",
          6301 => x"08",
          6302 => x"a4",
          6303 => x"11",
          6304 => x"55",
          6305 => x"16",
          6306 => x"08",
          6307 => x"75",
          6308 => x"e8",
          6309 => x"08",
          6310 => x"51",
          6311 => x"82",
          6312 => x"52",
          6313 => x"c9",
          6314 => x"52",
          6315 => x"c9",
          6316 => x"54",
          6317 => x"15",
          6318 => x"cc",
          6319 => x"93",
          6320 => x"17",
          6321 => x"06",
          6322 => x"90",
          6323 => x"82",
          6324 => x"8a",
          6325 => x"fc",
          6326 => x"70",
          6327 => x"d9",
          6328 => x"84",
          6329 => x"93",
          6330 => x"38",
          6331 => x"05",
          6332 => x"f1",
          6333 => x"93",
          6334 => x"82",
          6335 => x"87",
          6336 => x"84",
          6337 => x"72",
          6338 => x"0c",
          6339 => x"04",
          6340 => x"84",
          6341 => x"e4",
          6342 => x"80",
          6343 => x"84",
          6344 => x"38",
          6345 => x"08",
          6346 => x"34",
          6347 => x"82",
          6348 => x"83",
          6349 => x"ef",
          6350 => x"53",
          6351 => x"05",
          6352 => x"51",
          6353 => x"82",
          6354 => x"55",
          6355 => x"08",
          6356 => x"76",
          6357 => x"93",
          6358 => x"51",
          6359 => x"82",
          6360 => x"55",
          6361 => x"08",
          6362 => x"80",
          6363 => x"70",
          6364 => x"56",
          6365 => x"89",
          6366 => x"94",
          6367 => x"b2",
          6368 => x"05",
          6369 => x"2a",
          6370 => x"51",
          6371 => x"80",
          6372 => x"76",
          6373 => x"52",
          6374 => x"3f",
          6375 => x"08",
          6376 => x"8e",
          6377 => x"84",
          6378 => x"09",
          6379 => x"38",
          6380 => x"82",
          6381 => x"93",
          6382 => x"e4",
          6383 => x"6f",
          6384 => x"7a",
          6385 => x"9e",
          6386 => x"05",
          6387 => x"51",
          6388 => x"82",
          6389 => x"57",
          6390 => x"08",
          6391 => x"7b",
          6392 => x"94",
          6393 => x"55",
          6394 => x"73",
          6395 => x"ed",
          6396 => x"93",
          6397 => x"55",
          6398 => x"82",
          6399 => x"57",
          6400 => x"08",
          6401 => x"68",
          6402 => x"c9",
          6403 => x"93",
          6404 => x"82",
          6405 => x"82",
          6406 => x"52",
          6407 => x"a3",
          6408 => x"84",
          6409 => x"52",
          6410 => x"b8",
          6411 => x"84",
          6412 => x"93",
          6413 => x"a2",
          6414 => x"74",
          6415 => x"3f",
          6416 => x"08",
          6417 => x"84",
          6418 => x"69",
          6419 => x"d9",
          6420 => x"82",
          6421 => x"2e",
          6422 => x"52",
          6423 => x"cf",
          6424 => x"84",
          6425 => x"93",
          6426 => x"2e",
          6427 => x"84",
          6428 => x"06",
          6429 => x"57",
          6430 => x"76",
          6431 => x"9e",
          6432 => x"05",
          6433 => x"dc",
          6434 => x"90",
          6435 => x"81",
          6436 => x"56",
          6437 => x"80",
          6438 => x"02",
          6439 => x"81",
          6440 => x"70",
          6441 => x"56",
          6442 => x"81",
          6443 => x"78",
          6444 => x"38",
          6445 => x"99",
          6446 => x"81",
          6447 => x"18",
          6448 => x"18",
          6449 => x"58",
          6450 => x"33",
          6451 => x"ee",
          6452 => x"6f",
          6453 => x"af",
          6454 => x"8d",
          6455 => x"2e",
          6456 => x"8a",
          6457 => x"6f",
          6458 => x"af",
          6459 => x"0b",
          6460 => x"33",
          6461 => x"81",
          6462 => x"70",
          6463 => x"52",
          6464 => x"56",
          6465 => x"8d",
          6466 => x"70",
          6467 => x"51",
          6468 => x"f5",
          6469 => x"54",
          6470 => x"a7",
          6471 => x"74",
          6472 => x"38",
          6473 => x"73",
          6474 => x"81",
          6475 => x"81",
          6476 => x"39",
          6477 => x"81",
          6478 => x"74",
          6479 => x"81",
          6480 => x"91",
          6481 => x"6e",
          6482 => x"59",
          6483 => x"7a",
          6484 => x"5c",
          6485 => x"26",
          6486 => x"7a",
          6487 => x"93",
          6488 => x"3d",
          6489 => x"3d",
          6490 => x"8d",
          6491 => x"54",
          6492 => x"55",
          6493 => x"82",
          6494 => x"53",
          6495 => x"08",
          6496 => x"91",
          6497 => x"72",
          6498 => x"8c",
          6499 => x"73",
          6500 => x"38",
          6501 => x"70",
          6502 => x"81",
          6503 => x"57",
          6504 => x"73",
          6505 => x"08",
          6506 => x"94",
          6507 => x"75",
          6508 => x"97",
          6509 => x"11",
          6510 => x"2b",
          6511 => x"73",
          6512 => x"38",
          6513 => x"16",
          6514 => x"8f",
          6515 => x"84",
          6516 => x"78",
          6517 => x"55",
          6518 => x"ff",
          6519 => x"84",
          6520 => x"96",
          6521 => x"70",
          6522 => x"94",
          6523 => x"71",
          6524 => x"08",
          6525 => x"53",
          6526 => x"15",
          6527 => x"a6",
          6528 => x"74",
          6529 => x"3f",
          6530 => x"08",
          6531 => x"84",
          6532 => x"81",
          6533 => x"93",
          6534 => x"2e",
          6535 => x"82",
          6536 => x"88",
          6537 => x"98",
          6538 => x"80",
          6539 => x"38",
          6540 => x"80",
          6541 => x"77",
          6542 => x"08",
          6543 => x"0c",
          6544 => x"70",
          6545 => x"81",
          6546 => x"5a",
          6547 => x"2e",
          6548 => x"52",
          6549 => x"f9",
          6550 => x"84",
          6551 => x"93",
          6552 => x"38",
          6553 => x"08",
          6554 => x"73",
          6555 => x"c7",
          6556 => x"93",
          6557 => x"73",
          6558 => x"38",
          6559 => x"af",
          6560 => x"73",
          6561 => x"27",
          6562 => x"98",
          6563 => x"a0",
          6564 => x"08",
          6565 => x"0c",
          6566 => x"06",
          6567 => x"2e",
          6568 => x"52",
          6569 => x"a3",
          6570 => x"84",
          6571 => x"82",
          6572 => x"34",
          6573 => x"c4",
          6574 => x"91",
          6575 => x"53",
          6576 => x"89",
          6577 => x"84",
          6578 => x"94",
          6579 => x"8c",
          6580 => x"27",
          6581 => x"8c",
          6582 => x"15",
          6583 => x"07",
          6584 => x"16",
          6585 => x"ff",
          6586 => x"80",
          6587 => x"77",
          6588 => x"2e",
          6589 => x"9c",
          6590 => x"53",
          6591 => x"84",
          6592 => x"0d",
          6593 => x"0d",
          6594 => x"54",
          6595 => x"81",
          6596 => x"53",
          6597 => x"05",
          6598 => x"84",
          6599 => x"e7",
          6600 => x"84",
          6601 => x"93",
          6602 => x"ea",
          6603 => x"0c",
          6604 => x"51",
          6605 => x"82",
          6606 => x"55",
          6607 => x"08",
          6608 => x"ab",
          6609 => x"98",
          6610 => x"80",
          6611 => x"38",
          6612 => x"70",
          6613 => x"81",
          6614 => x"57",
          6615 => x"ad",
          6616 => x"08",
          6617 => x"d3",
          6618 => x"93",
          6619 => x"17",
          6620 => x"86",
          6621 => x"17",
          6622 => x"75",
          6623 => x"3f",
          6624 => x"08",
          6625 => x"2e",
          6626 => x"85",
          6627 => x"86",
          6628 => x"2e",
          6629 => x"76",
          6630 => x"73",
          6631 => x"0c",
          6632 => x"04",
          6633 => x"76",
          6634 => x"05",
          6635 => x"53",
          6636 => x"82",
          6637 => x"87",
          6638 => x"84",
          6639 => x"86",
          6640 => x"fb",
          6641 => x"79",
          6642 => x"05",
          6643 => x"56",
          6644 => x"3f",
          6645 => x"08",
          6646 => x"84",
          6647 => x"38",
          6648 => x"82",
          6649 => x"52",
          6650 => x"f8",
          6651 => x"84",
          6652 => x"ca",
          6653 => x"84",
          6654 => x"51",
          6655 => x"82",
          6656 => x"53",
          6657 => x"08",
          6658 => x"81",
          6659 => x"80",
          6660 => x"82",
          6661 => x"a6",
          6662 => x"73",
          6663 => x"3f",
          6664 => x"51",
          6665 => x"82",
          6666 => x"84",
          6667 => x"70",
          6668 => x"2c",
          6669 => x"84",
          6670 => x"51",
          6671 => x"82",
          6672 => x"87",
          6673 => x"ee",
          6674 => x"57",
          6675 => x"3d",
          6676 => x"3d",
          6677 => x"af",
          6678 => x"84",
          6679 => x"93",
          6680 => x"38",
          6681 => x"51",
          6682 => x"82",
          6683 => x"55",
          6684 => x"08",
          6685 => x"80",
          6686 => x"70",
          6687 => x"58",
          6688 => x"85",
          6689 => x"8d",
          6690 => x"2e",
          6691 => x"52",
          6692 => x"be",
          6693 => x"93",
          6694 => x"3d",
          6695 => x"3d",
          6696 => x"55",
          6697 => x"92",
          6698 => x"52",
          6699 => x"de",
          6700 => x"93",
          6701 => x"82",
          6702 => x"82",
          6703 => x"74",
          6704 => x"98",
          6705 => x"11",
          6706 => x"59",
          6707 => x"75",
          6708 => x"38",
          6709 => x"81",
          6710 => x"5b",
          6711 => x"82",
          6712 => x"39",
          6713 => x"08",
          6714 => x"59",
          6715 => x"09",
          6716 => x"38",
          6717 => x"57",
          6718 => x"3d",
          6719 => x"c1",
          6720 => x"93",
          6721 => x"2e",
          6722 => x"93",
          6723 => x"2e",
          6724 => x"93",
          6725 => x"70",
          6726 => x"08",
          6727 => x"7a",
          6728 => x"7f",
          6729 => x"54",
          6730 => x"77",
          6731 => x"80",
          6732 => x"15",
          6733 => x"84",
          6734 => x"75",
          6735 => x"52",
          6736 => x"52",
          6737 => x"8d",
          6738 => x"84",
          6739 => x"93",
          6740 => x"d6",
          6741 => x"33",
          6742 => x"1a",
          6743 => x"54",
          6744 => x"09",
          6745 => x"38",
          6746 => x"ff",
          6747 => x"82",
          6748 => x"83",
          6749 => x"70",
          6750 => x"25",
          6751 => x"59",
          6752 => x"9b",
          6753 => x"51",
          6754 => x"3f",
          6755 => x"08",
          6756 => x"70",
          6757 => x"25",
          6758 => x"59",
          6759 => x"75",
          6760 => x"7a",
          6761 => x"ff",
          6762 => x"7c",
          6763 => x"90",
          6764 => x"11",
          6765 => x"56",
          6766 => x"15",
          6767 => x"93",
          6768 => x"3d",
          6769 => x"3d",
          6770 => x"3d",
          6771 => x"70",
          6772 => x"dd",
          6773 => x"84",
          6774 => x"93",
          6775 => x"a8",
          6776 => x"33",
          6777 => x"a0",
          6778 => x"33",
          6779 => x"70",
          6780 => x"55",
          6781 => x"73",
          6782 => x"8e",
          6783 => x"08",
          6784 => x"18",
          6785 => x"80",
          6786 => x"38",
          6787 => x"08",
          6788 => x"08",
          6789 => x"c4",
          6790 => x"93",
          6791 => x"88",
          6792 => x"80",
          6793 => x"17",
          6794 => x"51",
          6795 => x"3f",
          6796 => x"08",
          6797 => x"81",
          6798 => x"81",
          6799 => x"84",
          6800 => x"09",
          6801 => x"38",
          6802 => x"39",
          6803 => x"77",
          6804 => x"84",
          6805 => x"08",
          6806 => x"98",
          6807 => x"82",
          6808 => x"52",
          6809 => x"bd",
          6810 => x"84",
          6811 => x"17",
          6812 => x"0c",
          6813 => x"80",
          6814 => x"73",
          6815 => x"75",
          6816 => x"38",
          6817 => x"34",
          6818 => x"82",
          6819 => x"89",
          6820 => x"e2",
          6821 => x"53",
          6822 => x"a4",
          6823 => x"3d",
          6824 => x"3f",
          6825 => x"08",
          6826 => x"84",
          6827 => x"38",
          6828 => x"3d",
          6829 => x"3d",
          6830 => x"d1",
          6831 => x"93",
          6832 => x"82",
          6833 => x"81",
          6834 => x"80",
          6835 => x"70",
          6836 => x"81",
          6837 => x"56",
          6838 => x"81",
          6839 => x"98",
          6840 => x"74",
          6841 => x"38",
          6842 => x"05",
          6843 => x"06",
          6844 => x"55",
          6845 => x"38",
          6846 => x"51",
          6847 => x"82",
          6848 => x"74",
          6849 => x"81",
          6850 => x"56",
          6851 => x"80",
          6852 => x"54",
          6853 => x"08",
          6854 => x"2e",
          6855 => x"73",
          6856 => x"84",
          6857 => x"52",
          6858 => x"52",
          6859 => x"3f",
          6860 => x"08",
          6861 => x"84",
          6862 => x"38",
          6863 => x"08",
          6864 => x"cc",
          6865 => x"93",
          6866 => x"82",
          6867 => x"86",
          6868 => x"80",
          6869 => x"93",
          6870 => x"2e",
          6871 => x"93",
          6872 => x"c0",
          6873 => x"ce",
          6874 => x"93",
          6875 => x"93",
          6876 => x"70",
          6877 => x"08",
          6878 => x"51",
          6879 => x"80",
          6880 => x"73",
          6881 => x"38",
          6882 => x"52",
          6883 => x"95",
          6884 => x"84",
          6885 => x"8c",
          6886 => x"ff",
          6887 => x"82",
          6888 => x"55",
          6889 => x"84",
          6890 => x"0d",
          6891 => x"0d",
          6892 => x"3d",
          6893 => x"9a",
          6894 => x"cb",
          6895 => x"84",
          6896 => x"93",
          6897 => x"b0",
          6898 => x"69",
          6899 => x"70",
          6900 => x"97",
          6901 => x"84",
          6902 => x"93",
          6903 => x"38",
          6904 => x"94",
          6905 => x"84",
          6906 => x"09",
          6907 => x"88",
          6908 => x"df",
          6909 => x"85",
          6910 => x"51",
          6911 => x"74",
          6912 => x"78",
          6913 => x"8a",
          6914 => x"57",
          6915 => x"82",
          6916 => x"75",
          6917 => x"93",
          6918 => x"38",
          6919 => x"93",
          6920 => x"2e",
          6921 => x"83",
          6922 => x"82",
          6923 => x"ff",
          6924 => x"06",
          6925 => x"54",
          6926 => x"73",
          6927 => x"82",
          6928 => x"52",
          6929 => x"a4",
          6930 => x"84",
          6931 => x"93",
          6932 => x"9a",
          6933 => x"a0",
          6934 => x"51",
          6935 => x"3f",
          6936 => x"0b",
          6937 => x"78",
          6938 => x"bf",
          6939 => x"88",
          6940 => x"80",
          6941 => x"ff",
          6942 => x"75",
          6943 => x"11",
          6944 => x"f8",
          6945 => x"78",
          6946 => x"80",
          6947 => x"ff",
          6948 => x"78",
          6949 => x"80",
          6950 => x"7f",
          6951 => x"d4",
          6952 => x"c9",
          6953 => x"54",
          6954 => x"15",
          6955 => x"cb",
          6956 => x"93",
          6957 => x"82",
          6958 => x"b2",
          6959 => x"b2",
          6960 => x"96",
          6961 => x"b5",
          6962 => x"53",
          6963 => x"51",
          6964 => x"64",
          6965 => x"8b",
          6966 => x"54",
          6967 => x"15",
          6968 => x"ff",
          6969 => x"82",
          6970 => x"54",
          6971 => x"53",
          6972 => x"51",
          6973 => x"3f",
          6974 => x"84",
          6975 => x"0d",
          6976 => x"0d",
          6977 => x"05",
          6978 => x"3f",
          6979 => x"3d",
          6980 => x"52",
          6981 => x"d5",
          6982 => x"93",
          6983 => x"82",
          6984 => x"82",
          6985 => x"4d",
          6986 => x"52",
          6987 => x"52",
          6988 => x"3f",
          6989 => x"08",
          6990 => x"84",
          6991 => x"38",
          6992 => x"05",
          6993 => x"06",
          6994 => x"73",
          6995 => x"a0",
          6996 => x"08",
          6997 => x"ff",
          6998 => x"ff",
          6999 => x"ac",
          7000 => x"92",
          7001 => x"54",
          7002 => x"3f",
          7003 => x"52",
          7004 => x"f7",
          7005 => x"84",
          7006 => x"93",
          7007 => x"38",
          7008 => x"09",
          7009 => x"38",
          7010 => x"08",
          7011 => x"88",
          7012 => x"39",
          7013 => x"08",
          7014 => x"81",
          7015 => x"38",
          7016 => x"b1",
          7017 => x"84",
          7018 => x"93",
          7019 => x"c8",
          7020 => x"93",
          7021 => x"ff",
          7022 => x"8d",
          7023 => x"b4",
          7024 => x"af",
          7025 => x"17",
          7026 => x"33",
          7027 => x"70",
          7028 => x"55",
          7029 => x"38",
          7030 => x"54",
          7031 => x"34",
          7032 => x"0b",
          7033 => x"8b",
          7034 => x"84",
          7035 => x"06",
          7036 => x"73",
          7037 => x"e5",
          7038 => x"2e",
          7039 => x"75",
          7040 => x"c6",
          7041 => x"93",
          7042 => x"78",
          7043 => x"bb",
          7044 => x"82",
          7045 => x"80",
          7046 => x"38",
          7047 => x"08",
          7048 => x"ff",
          7049 => x"82",
          7050 => x"79",
          7051 => x"58",
          7052 => x"93",
          7053 => x"c0",
          7054 => x"33",
          7055 => x"2e",
          7056 => x"99",
          7057 => x"75",
          7058 => x"c6",
          7059 => x"54",
          7060 => x"15",
          7061 => x"82",
          7062 => x"9c",
          7063 => x"c8",
          7064 => x"93",
          7065 => x"82",
          7066 => x"8c",
          7067 => x"ff",
          7068 => x"82",
          7069 => x"55",
          7070 => x"84",
          7071 => x"0d",
          7072 => x"0d",
          7073 => x"05",
          7074 => x"05",
          7075 => x"33",
          7076 => x"53",
          7077 => x"05",
          7078 => x"51",
          7079 => x"82",
          7080 => x"55",
          7081 => x"08",
          7082 => x"78",
          7083 => x"95",
          7084 => x"51",
          7085 => x"82",
          7086 => x"55",
          7087 => x"08",
          7088 => x"80",
          7089 => x"81",
          7090 => x"86",
          7091 => x"38",
          7092 => x"61",
          7093 => x"12",
          7094 => x"7a",
          7095 => x"51",
          7096 => x"74",
          7097 => x"78",
          7098 => x"83",
          7099 => x"51",
          7100 => x"3f",
          7101 => x"08",
          7102 => x"93",
          7103 => x"3d",
          7104 => x"3d",
          7105 => x"82",
          7106 => x"d0",
          7107 => x"3d",
          7108 => x"3f",
          7109 => x"08",
          7110 => x"84",
          7111 => x"38",
          7112 => x"52",
          7113 => x"05",
          7114 => x"3f",
          7115 => x"08",
          7116 => x"84",
          7117 => x"02",
          7118 => x"33",
          7119 => x"54",
          7120 => x"a6",
          7121 => x"22",
          7122 => x"71",
          7123 => x"53",
          7124 => x"51",
          7125 => x"3f",
          7126 => x"0b",
          7127 => x"76",
          7128 => x"b8",
          7129 => x"84",
          7130 => x"82",
          7131 => x"93",
          7132 => x"ea",
          7133 => x"6b",
          7134 => x"53",
          7135 => x"05",
          7136 => x"51",
          7137 => x"82",
          7138 => x"82",
          7139 => x"30",
          7140 => x"84",
          7141 => x"25",
          7142 => x"79",
          7143 => x"85",
          7144 => x"75",
          7145 => x"73",
          7146 => x"f9",
          7147 => x"80",
          7148 => x"8d",
          7149 => x"54",
          7150 => x"3f",
          7151 => x"08",
          7152 => x"84",
          7153 => x"38",
          7154 => x"51",
          7155 => x"82",
          7156 => x"57",
          7157 => x"08",
          7158 => x"93",
          7159 => x"93",
          7160 => x"5b",
          7161 => x"18",
          7162 => x"18",
          7163 => x"74",
          7164 => x"81",
          7165 => x"78",
          7166 => x"8b",
          7167 => x"54",
          7168 => x"75",
          7169 => x"38",
          7170 => x"1b",
          7171 => x"55",
          7172 => x"2e",
          7173 => x"39",
          7174 => x"09",
          7175 => x"38",
          7176 => x"80",
          7177 => x"70",
          7178 => x"25",
          7179 => x"80",
          7180 => x"38",
          7181 => x"bc",
          7182 => x"11",
          7183 => x"ff",
          7184 => x"82",
          7185 => x"57",
          7186 => x"08",
          7187 => x"70",
          7188 => x"80",
          7189 => x"83",
          7190 => x"80",
          7191 => x"84",
          7192 => x"a7",
          7193 => x"b4",
          7194 => x"ad",
          7195 => x"93",
          7196 => x"0c",
          7197 => x"84",
          7198 => x"0d",
          7199 => x"0d",
          7200 => x"3d",
          7201 => x"52",
          7202 => x"ce",
          7203 => x"93",
          7204 => x"93",
          7205 => x"54",
          7206 => x"08",
          7207 => x"8b",
          7208 => x"8b",
          7209 => x"59",
          7210 => x"3f",
          7211 => x"33",
          7212 => x"06",
          7213 => x"57",
          7214 => x"81",
          7215 => x"58",
          7216 => x"06",
          7217 => x"4e",
          7218 => x"ff",
          7219 => x"82",
          7220 => x"80",
          7221 => x"6c",
          7222 => x"53",
          7223 => x"ae",
          7224 => x"93",
          7225 => x"2e",
          7226 => x"88",
          7227 => x"6d",
          7228 => x"55",
          7229 => x"93",
          7230 => x"ff",
          7231 => x"83",
          7232 => x"51",
          7233 => x"26",
          7234 => x"15",
          7235 => x"ff",
          7236 => x"80",
          7237 => x"87",
          7238 => x"f0",
          7239 => x"74",
          7240 => x"38",
          7241 => x"80",
          7242 => x"ae",
          7243 => x"93",
          7244 => x"38",
          7245 => x"27",
          7246 => x"89",
          7247 => x"8b",
          7248 => x"27",
          7249 => x"55",
          7250 => x"81",
          7251 => x"8f",
          7252 => x"2a",
          7253 => x"70",
          7254 => x"34",
          7255 => x"74",
          7256 => x"05",
          7257 => x"17",
          7258 => x"70",
          7259 => x"52",
          7260 => x"73",
          7261 => x"c8",
          7262 => x"33",
          7263 => x"73",
          7264 => x"81",
          7265 => x"80",
          7266 => x"02",
          7267 => x"76",
          7268 => x"51",
          7269 => x"2e",
          7270 => x"87",
          7271 => x"57",
          7272 => x"79",
          7273 => x"80",
          7274 => x"70",
          7275 => x"ba",
          7276 => x"93",
          7277 => x"82",
          7278 => x"80",
          7279 => x"52",
          7280 => x"bf",
          7281 => x"93",
          7282 => x"82",
          7283 => x"8d",
          7284 => x"c4",
          7285 => x"e5",
          7286 => x"c6",
          7287 => x"84",
          7288 => x"09",
          7289 => x"cc",
          7290 => x"76",
          7291 => x"c4",
          7292 => x"74",
          7293 => x"b0",
          7294 => x"84",
          7295 => x"93",
          7296 => x"38",
          7297 => x"93",
          7298 => x"67",
          7299 => x"db",
          7300 => x"88",
          7301 => x"34",
          7302 => x"52",
          7303 => x"ab",
          7304 => x"54",
          7305 => x"15",
          7306 => x"ff",
          7307 => x"82",
          7308 => x"54",
          7309 => x"82",
          7310 => x"9c",
          7311 => x"f2",
          7312 => x"62",
          7313 => x"80",
          7314 => x"93",
          7315 => x"55",
          7316 => x"5e",
          7317 => x"3f",
          7318 => x"08",
          7319 => x"84",
          7320 => x"38",
          7321 => x"58",
          7322 => x"38",
          7323 => x"97",
          7324 => x"08",
          7325 => x"38",
          7326 => x"70",
          7327 => x"81",
          7328 => x"55",
          7329 => x"87",
          7330 => x"39",
          7331 => x"90",
          7332 => x"82",
          7333 => x"8a",
          7334 => x"89",
          7335 => x"7f",
          7336 => x"56",
          7337 => x"3f",
          7338 => x"06",
          7339 => x"72",
          7340 => x"82",
          7341 => x"05",
          7342 => x"7c",
          7343 => x"55",
          7344 => x"27",
          7345 => x"16",
          7346 => x"83",
          7347 => x"76",
          7348 => x"80",
          7349 => x"79",
          7350 => x"99",
          7351 => x"7f",
          7352 => x"14",
          7353 => x"83",
          7354 => x"82",
          7355 => x"81",
          7356 => x"38",
          7357 => x"08",
          7358 => x"95",
          7359 => x"84",
          7360 => x"81",
          7361 => x"7b",
          7362 => x"06",
          7363 => x"39",
          7364 => x"56",
          7365 => x"09",
          7366 => x"b9",
          7367 => x"80",
          7368 => x"80",
          7369 => x"78",
          7370 => x"7a",
          7371 => x"38",
          7372 => x"73",
          7373 => x"81",
          7374 => x"ff",
          7375 => x"74",
          7376 => x"ff",
          7377 => x"82",
          7378 => x"58",
          7379 => x"08",
          7380 => x"74",
          7381 => x"16",
          7382 => x"73",
          7383 => x"39",
          7384 => x"7e",
          7385 => x"0c",
          7386 => x"2e",
          7387 => x"88",
          7388 => x"8c",
          7389 => x"1a",
          7390 => x"07",
          7391 => x"1b",
          7392 => x"08",
          7393 => x"16",
          7394 => x"75",
          7395 => x"38",
          7396 => x"90",
          7397 => x"15",
          7398 => x"54",
          7399 => x"34",
          7400 => x"82",
          7401 => x"90",
          7402 => x"e9",
          7403 => x"6d",
          7404 => x"80",
          7405 => x"9d",
          7406 => x"5c",
          7407 => x"3f",
          7408 => x"0b",
          7409 => x"08",
          7410 => x"38",
          7411 => x"08",
          7412 => x"93",
          7413 => x"08",
          7414 => x"80",
          7415 => x"80",
          7416 => x"93",
          7417 => x"ff",
          7418 => x"52",
          7419 => x"a0",
          7420 => x"93",
          7421 => x"ff",
          7422 => x"06",
          7423 => x"56",
          7424 => x"38",
          7425 => x"70",
          7426 => x"55",
          7427 => x"8b",
          7428 => x"3d",
          7429 => x"83",
          7430 => x"ff",
          7431 => x"82",
          7432 => x"99",
          7433 => x"74",
          7434 => x"38",
          7435 => x"80",
          7436 => x"ff",
          7437 => x"55",
          7438 => x"83",
          7439 => x"78",
          7440 => x"38",
          7441 => x"26",
          7442 => x"81",
          7443 => x"8b",
          7444 => x"79",
          7445 => x"80",
          7446 => x"93",
          7447 => x"39",
          7448 => x"6e",
          7449 => x"89",
          7450 => x"48",
          7451 => x"83",
          7452 => x"61",
          7453 => x"25",
          7454 => x"55",
          7455 => x"8a",
          7456 => x"3d",
          7457 => x"81",
          7458 => x"ff",
          7459 => x"81",
          7460 => x"84",
          7461 => x"38",
          7462 => x"70",
          7463 => x"93",
          7464 => x"56",
          7465 => x"38",
          7466 => x"55",
          7467 => x"75",
          7468 => x"38",
          7469 => x"70",
          7470 => x"ff",
          7471 => x"83",
          7472 => x"78",
          7473 => x"89",
          7474 => x"81",
          7475 => x"06",
          7476 => x"80",
          7477 => x"77",
          7478 => x"74",
          7479 => x"8d",
          7480 => x"06",
          7481 => x"2e",
          7482 => x"77",
          7483 => x"93",
          7484 => x"74",
          7485 => x"cb",
          7486 => x"7d",
          7487 => x"81",
          7488 => x"38",
          7489 => x"66",
          7490 => x"81",
          7491 => x"94",
          7492 => x"74",
          7493 => x"38",
          7494 => x"98",
          7495 => x"94",
          7496 => x"82",
          7497 => x"57",
          7498 => x"80",
          7499 => x"76",
          7500 => x"38",
          7501 => x"51",
          7502 => x"3f",
          7503 => x"08",
          7504 => x"87",
          7505 => x"2a",
          7506 => x"5c",
          7507 => x"93",
          7508 => x"80",
          7509 => x"44",
          7510 => x"0a",
          7511 => x"ec",
          7512 => x"39",
          7513 => x"66",
          7514 => x"81",
          7515 => x"84",
          7516 => x"74",
          7517 => x"38",
          7518 => x"98",
          7519 => x"84",
          7520 => x"82",
          7521 => x"57",
          7522 => x"80",
          7523 => x"76",
          7524 => x"38",
          7525 => x"51",
          7526 => x"3f",
          7527 => x"08",
          7528 => x"57",
          7529 => x"08",
          7530 => x"96",
          7531 => x"82",
          7532 => x"10",
          7533 => x"08",
          7534 => x"72",
          7535 => x"59",
          7536 => x"ff",
          7537 => x"5d",
          7538 => x"44",
          7539 => x"11",
          7540 => x"70",
          7541 => x"71",
          7542 => x"06",
          7543 => x"52",
          7544 => x"40",
          7545 => x"09",
          7546 => x"38",
          7547 => x"18",
          7548 => x"39",
          7549 => x"79",
          7550 => x"70",
          7551 => x"58",
          7552 => x"76",
          7553 => x"38",
          7554 => x"7d",
          7555 => x"70",
          7556 => x"55",
          7557 => x"3f",
          7558 => x"08",
          7559 => x"2e",
          7560 => x"9b",
          7561 => x"84",
          7562 => x"f5",
          7563 => x"38",
          7564 => x"38",
          7565 => x"59",
          7566 => x"38",
          7567 => x"7d",
          7568 => x"81",
          7569 => x"38",
          7570 => x"0b",
          7571 => x"08",
          7572 => x"78",
          7573 => x"1a",
          7574 => x"c0",
          7575 => x"74",
          7576 => x"39",
          7577 => x"55",
          7578 => x"8f",
          7579 => x"fd",
          7580 => x"93",
          7581 => x"f5",
          7582 => x"78",
          7583 => x"79",
          7584 => x"80",
          7585 => x"f1",
          7586 => x"39",
          7587 => x"81",
          7588 => x"06",
          7589 => x"55",
          7590 => x"27",
          7591 => x"81",
          7592 => x"56",
          7593 => x"38",
          7594 => x"80",
          7595 => x"ff",
          7596 => x"8b",
          7597 => x"ac",
          7598 => x"ff",
          7599 => x"84",
          7600 => x"1b",
          7601 => x"b3",
          7602 => x"1c",
          7603 => x"ff",
          7604 => x"8e",
          7605 => x"a1",
          7606 => x"0b",
          7607 => x"7d",
          7608 => x"30",
          7609 => x"84",
          7610 => x"51",
          7611 => x"51",
          7612 => x"3f",
          7613 => x"83",
          7614 => x"90",
          7615 => x"ff",
          7616 => x"93",
          7617 => x"a0",
          7618 => x"39",
          7619 => x"1b",
          7620 => x"85",
          7621 => x"95",
          7622 => x"52",
          7623 => x"ff",
          7624 => x"81",
          7625 => x"1b",
          7626 => x"cf",
          7627 => x"9c",
          7628 => x"a0",
          7629 => x"83",
          7630 => x"06",
          7631 => x"82",
          7632 => x"52",
          7633 => x"51",
          7634 => x"3f",
          7635 => x"1b",
          7636 => x"c5",
          7637 => x"ac",
          7638 => x"a0",
          7639 => x"52",
          7640 => x"ff",
          7641 => x"86",
          7642 => x"51",
          7643 => x"3f",
          7644 => x"80",
          7645 => x"a9",
          7646 => x"1c",
          7647 => x"81",
          7648 => x"80",
          7649 => x"ae",
          7650 => x"b2",
          7651 => x"1b",
          7652 => x"85",
          7653 => x"ff",
          7654 => x"96",
          7655 => x"9f",
          7656 => x"80",
          7657 => x"34",
          7658 => x"1c",
          7659 => x"81",
          7660 => x"ab",
          7661 => x"a0",
          7662 => x"d4",
          7663 => x"fe",
          7664 => x"59",
          7665 => x"3f",
          7666 => x"53",
          7667 => x"51",
          7668 => x"3f",
          7669 => x"93",
          7670 => x"e7",
          7671 => x"2e",
          7672 => x"80",
          7673 => x"54",
          7674 => x"53",
          7675 => x"51",
          7676 => x"3f",
          7677 => x"80",
          7678 => x"ff",
          7679 => x"84",
          7680 => x"d2",
          7681 => x"ff",
          7682 => x"86",
          7683 => x"f2",
          7684 => x"1b",
          7685 => x"81",
          7686 => x"52",
          7687 => x"51",
          7688 => x"3f",
          7689 => x"ec",
          7690 => x"9e",
          7691 => x"d4",
          7692 => x"51",
          7693 => x"3f",
          7694 => x"87",
          7695 => x"52",
          7696 => x"9a",
          7697 => x"54",
          7698 => x"7a",
          7699 => x"ff",
          7700 => x"65",
          7701 => x"7a",
          7702 => x"8f",
          7703 => x"80",
          7704 => x"2e",
          7705 => x"9a",
          7706 => x"7a",
          7707 => x"a9",
          7708 => x"84",
          7709 => x"9e",
          7710 => x"0a",
          7711 => x"51",
          7712 => x"ff",
          7713 => x"7d",
          7714 => x"38",
          7715 => x"52",
          7716 => x"9e",
          7717 => x"55",
          7718 => x"62",
          7719 => x"74",
          7720 => x"75",
          7721 => x"7e",
          7722 => x"fe",
          7723 => x"84",
          7724 => x"38",
          7725 => x"82",
          7726 => x"52",
          7727 => x"9e",
          7728 => x"16",
          7729 => x"56",
          7730 => x"38",
          7731 => x"77",
          7732 => x"8d",
          7733 => x"7d",
          7734 => x"38",
          7735 => x"57",
          7736 => x"83",
          7737 => x"76",
          7738 => x"7a",
          7739 => x"ff",
          7740 => x"82",
          7741 => x"81",
          7742 => x"16",
          7743 => x"56",
          7744 => x"38",
          7745 => x"83",
          7746 => x"86",
          7747 => x"ff",
          7748 => x"38",
          7749 => x"82",
          7750 => x"81",
          7751 => x"06",
          7752 => x"fe",
          7753 => x"53",
          7754 => x"51",
          7755 => x"3f",
          7756 => x"52",
          7757 => x"9c",
          7758 => x"be",
          7759 => x"75",
          7760 => x"81",
          7761 => x"0b",
          7762 => x"77",
          7763 => x"75",
          7764 => x"60",
          7765 => x"80",
          7766 => x"75",
          7767 => x"fb",
          7768 => x"85",
          7769 => x"93",
          7770 => x"2a",
          7771 => x"75",
          7772 => x"82",
          7773 => x"87",
          7774 => x"52",
          7775 => x"51",
          7776 => x"3f",
          7777 => x"ca",
          7778 => x"9c",
          7779 => x"54",
          7780 => x"52",
          7781 => x"98",
          7782 => x"56",
          7783 => x"08",
          7784 => x"53",
          7785 => x"51",
          7786 => x"3f",
          7787 => x"93",
          7788 => x"38",
          7789 => x"56",
          7790 => x"56",
          7791 => x"93",
          7792 => x"75",
          7793 => x"0c",
          7794 => x"04",
          7795 => x"7d",
          7796 => x"80",
          7797 => x"05",
          7798 => x"76",
          7799 => x"38",
          7800 => x"11",
          7801 => x"53",
          7802 => x"79",
          7803 => x"3f",
          7804 => x"09",
          7805 => x"38",
          7806 => x"55",
          7807 => x"db",
          7808 => x"70",
          7809 => x"34",
          7810 => x"74",
          7811 => x"81",
          7812 => x"80",
          7813 => x"55",
          7814 => x"76",
          7815 => x"93",
          7816 => x"3d",
          7817 => x"3d",
          7818 => x"84",
          7819 => x"33",
          7820 => x"8a",
          7821 => x"06",
          7822 => x"52",
          7823 => x"3f",
          7824 => x"56",
          7825 => x"be",
          7826 => x"08",
          7827 => x"05",
          7828 => x"75",
          7829 => x"56",
          7830 => x"a1",
          7831 => x"fc",
          7832 => x"53",
          7833 => x"76",
          7834 => x"dc",
          7835 => x"32",
          7836 => x"72",
          7837 => x"70",
          7838 => x"56",
          7839 => x"18",
          7840 => x"88",
          7841 => x"3d",
          7842 => x"3d",
          7843 => x"11",
          7844 => x"80",
          7845 => x"38",
          7846 => x"05",
          7847 => x"8c",
          7848 => x"08",
          7849 => x"3f",
          7850 => x"08",
          7851 => x"16",
          7852 => x"09",
          7853 => x"38",
          7854 => x"55",
          7855 => x"55",
          7856 => x"84",
          7857 => x"0d",
          7858 => x"0d",
          7859 => x"cc",
          7860 => x"73",
          7861 => x"93",
          7862 => x"0c",
          7863 => x"04",
          7864 => x"02",
          7865 => x"33",
          7866 => x"3d",
          7867 => x"54",
          7868 => x"52",
          7869 => x"ae",
          7870 => x"ff",
          7871 => x"3d",
          7872 => x"3d",
          7873 => x"08",
          7874 => x"59",
          7875 => x"80",
          7876 => x"39",
          7877 => x"0c",
          7878 => x"54",
          7879 => x"74",
          7880 => x"a0",
          7881 => x"06",
          7882 => x"15",
          7883 => x"80",
          7884 => x"29",
          7885 => x"05",
          7886 => x"56",
          7887 => x"3f",
          7888 => x"08",
          7889 => x"08",
          7890 => x"76",
          7891 => x"fe",
          7892 => x"82",
          7893 => x"8b",
          7894 => x"33",
          7895 => x"2e",
          7896 => x"81",
          7897 => x"ff",
          7898 => x"98",
          7899 => x"38",
          7900 => x"82",
          7901 => x"8a",
          7902 => x"ff",
          7903 => x"52",
          7904 => x"81",
          7905 => x"84",
          7906 => x"98",
          7907 => x"08",
          7908 => x"cc",
          7909 => x"39",
          7910 => x"51",
          7911 => x"82",
          7912 => x"80",
          7913 => x"83",
          7914 => x"eb",
          7915 => x"90",
          7916 => x"39",
          7917 => x"51",
          7918 => x"82",
          7919 => x"80",
          7920 => x"83",
          7921 => x"cf",
          7922 => x"dc",
          7923 => x"39",
          7924 => x"51",
          7925 => x"82",
          7926 => x"bb",
          7927 => x"a8",
          7928 => x"82",
          7929 => x"af",
          7930 => x"e8",
          7931 => x"82",
          7932 => x"a3",
          7933 => x"9c",
          7934 => x"82",
          7935 => x"97",
          7936 => x"c8",
          7937 => x"82",
          7938 => x"8b",
          7939 => x"f8",
          7940 => x"82",
          7941 => x"fe",
          7942 => x"83",
          7943 => x"fb",
          7944 => x"79",
          7945 => x"87",
          7946 => x"38",
          7947 => x"87",
          7948 => x"91",
          7949 => x"52",
          7950 => x"d2",
          7951 => x"93",
          7952 => x"75",
          7953 => x"93",
          7954 => x"84",
          7955 => x"53",
          7956 => x"86",
          7957 => x"f7",
          7958 => x"3d",
          7959 => x"3d",
          7960 => x"84",
          7961 => x"05",
          7962 => x"80",
          7963 => x"70",
          7964 => x"25",
          7965 => x"59",
          7966 => x"87",
          7967 => x"38",
          7968 => x"76",
          7969 => x"ff",
          7970 => x"93",
          7971 => x"80",
          7972 => x"76",
          7973 => x"70",
          7974 => x"bf",
          7975 => x"93",
          7976 => x"82",
          7977 => x"b8",
          7978 => x"84",
          7979 => x"98",
          7980 => x"93",
          7981 => x"96",
          7982 => x"54",
          7983 => x"77",
          7984 => x"c4",
          7985 => x"93",
          7986 => x"82",
          7987 => x"90",
          7988 => x"74",
          7989 => x"38",
          7990 => x"19",
          7991 => x"39",
          7992 => x"05",
          7993 => x"3f",
          7994 => x"78",
          7995 => x"7b",
          7996 => x"2a",
          7997 => x"57",
          7998 => x"80",
          7999 => x"82",
          8000 => x"87",
          8001 => x"08",
          8002 => x"fe",
          8003 => x"56",
          8004 => x"84",
          8005 => x"0d",
          8006 => x"0d",
          8007 => x"05",
          8008 => x"57",
          8009 => x"80",
          8010 => x"79",
          8011 => x"3f",
          8012 => x"08",
          8013 => x"80",
          8014 => x"75",
          8015 => x"38",
          8016 => x"55",
          8017 => x"93",
          8018 => x"52",
          8019 => x"2d",
          8020 => x"08",
          8021 => x"77",
          8022 => x"93",
          8023 => x"3d",
          8024 => x"3d",
          8025 => x"63",
          8026 => x"80",
          8027 => x"73",
          8028 => x"41",
          8029 => x"5e",
          8030 => x"52",
          8031 => x"51",
          8032 => x"3f",
          8033 => x"51",
          8034 => x"3f",
          8035 => x"79",
          8036 => x"38",
          8037 => x"89",
          8038 => x"2e",
          8039 => x"c6",
          8040 => x"53",
          8041 => x"8e",
          8042 => x"52",
          8043 => x"51",
          8044 => x"3f",
          8045 => x"86",
          8046 => x"ef",
          8047 => x"15",
          8048 => x"39",
          8049 => x"72",
          8050 => x"38",
          8051 => x"82",
          8052 => x"fe",
          8053 => x"89",
          8054 => x"d4",
          8055 => x"e8",
          8056 => x"55",
          8057 => x"18",
          8058 => x"27",
          8059 => x"33",
          8060 => x"e0",
          8061 => x"b4",
          8062 => x"82",
          8063 => x"fe",
          8064 => x"81",
          8065 => x"51",
          8066 => x"3f",
          8067 => x"82",
          8068 => x"fe",
          8069 => x"80",
          8070 => x"27",
          8071 => x"18",
          8072 => x"53",
          8073 => x"7a",
          8074 => x"81",
          8075 => x"9f",
          8076 => x"38",
          8077 => x"73",
          8078 => x"ff",
          8079 => x"72",
          8080 => x"38",
          8081 => x"26",
          8082 => x"51",
          8083 => x"51",
          8084 => x"3f",
          8085 => x"c1",
          8086 => x"f0",
          8087 => x"e8",
          8088 => x"79",
          8089 => x"fe",
          8090 => x"82",
          8091 => x"98",
          8092 => x"2c",
          8093 => x"a0",
          8094 => x"06",
          8095 => x"dd",
          8096 => x"93",
          8097 => x"2b",
          8098 => x"70",
          8099 => x"30",
          8100 => x"70",
          8101 => x"07",
          8102 => x"06",
          8103 => x"59",
          8104 => x"80",
          8105 => x"38",
          8106 => x"09",
          8107 => x"38",
          8108 => x"39",
          8109 => x"72",
          8110 => x"be",
          8111 => x"72",
          8112 => x"0c",
          8113 => x"04",
          8114 => x"02",
          8115 => x"82",
          8116 => x"82",
          8117 => x"55",
          8118 => x"3f",
          8119 => x"22",
          8120 => x"d5",
          8121 => x"88",
          8122 => x"94",
          8123 => x"b5",
          8124 => x"87",
          8125 => x"f2",
          8126 => x"80",
          8127 => x"fe",
          8128 => x"86",
          8129 => x"fe",
          8130 => x"c0",
          8131 => x"53",
          8132 => x"3f",
          8133 => x"d8",
          8134 => x"87",
          8135 => x"da",
          8136 => x"51",
          8137 => x"3f",
          8138 => x"70",
          8139 => x"52",
          8140 => x"95",
          8141 => x"fe",
          8142 => x"82",
          8143 => x"fe",
          8144 => x"80",
          8145 => x"ca",
          8146 => x"2a",
          8147 => x"51",
          8148 => x"2e",
          8149 => x"51",
          8150 => x"3f",
          8151 => x"51",
          8152 => x"3f",
          8153 => x"d8",
          8154 => x"83",
          8155 => x"06",
          8156 => x"80",
          8157 => x"81",
          8158 => x"96",
          8159 => x"f8",
          8160 => x"8e",
          8161 => x"fe",
          8162 => x"72",
          8163 => x"81",
          8164 => x"71",
          8165 => x"38",
          8166 => x"d7",
          8167 => x"88",
          8168 => x"d9",
          8169 => x"51",
          8170 => x"3f",
          8171 => x"70",
          8172 => x"52",
          8173 => x"95",
          8174 => x"fe",
          8175 => x"82",
          8176 => x"fe",
          8177 => x"80",
          8178 => x"c6",
          8179 => x"2a",
          8180 => x"51",
          8181 => x"2e",
          8182 => x"51",
          8183 => x"3f",
          8184 => x"51",
          8185 => x"3f",
          8186 => x"d7",
          8187 => x"87",
          8188 => x"06",
          8189 => x"80",
          8190 => x"81",
          8191 => x"92",
          8192 => x"c8",
          8193 => x"8a",
          8194 => x"fe",
          8195 => x"72",
          8196 => x"81",
          8197 => x"71",
          8198 => x"38",
          8199 => x"d6",
          8200 => x"88",
          8201 => x"d8",
          8202 => x"51",
          8203 => x"3f",
          8204 => x"3f",
          8205 => x"04",
          8206 => x"77",
          8207 => x"a3",
          8208 => x"55",
          8209 => x"52",
          8210 => x"ce",
          8211 => x"8f",
          8212 => x"73",
          8213 => x"53",
          8214 => x"52",
          8215 => x"51",
          8216 => x"3f",
          8217 => x"08",
          8218 => x"93",
          8219 => x"80",
          8220 => x"31",
          8221 => x"73",
          8222 => x"34",
          8223 => x"33",
          8224 => x"2e",
          8225 => x"ac",
          8226 => x"9c",
          8227 => x"75",
          8228 => x"3f",
          8229 => x"08",
          8230 => x"38",
          8231 => x"08",
          8232 => x"a4",
          8233 => x"82",
          8234 => x"c4",
          8235 => x"0b",
          8236 => x"34",
          8237 => x"33",
          8238 => x"2e",
          8239 => x"89",
          8240 => x"75",
          8241 => x"e4",
          8242 => x"82",
          8243 => x"87",
          8244 => x"ce",
          8245 => x"70",
          8246 => x"98",
          8247 => x"81",
          8248 => x"ff",
          8249 => x"82",
          8250 => x"81",
          8251 => x"78",
          8252 => x"81",
          8253 => x"82",
          8254 => x"96",
          8255 => x"59",
          8256 => x"3f",
          8257 => x"52",
          8258 => x"51",
          8259 => x"3f",
          8260 => x"08",
          8261 => x"38",
          8262 => x"51",
          8263 => x"81",
          8264 => x"82",
          8265 => x"fe",
          8266 => x"96",
          8267 => x"5a",
          8268 => x"79",
          8269 => x"3f",
          8270 => x"84",
          8271 => x"c2",
          8272 => x"84",
          8273 => x"70",
          8274 => x"59",
          8275 => x"2e",
          8276 => x"78",
          8277 => x"80",
          8278 => x"ab",
          8279 => x"38",
          8280 => x"a4",
          8281 => x"2e",
          8282 => x"78",
          8283 => x"38",
          8284 => x"ff",
          8285 => x"a5",
          8286 => x"2e",
          8287 => x"78",
          8288 => x"b1",
          8289 => x"39",
          8290 => x"85",
          8291 => x"bd",
          8292 => x"78",
          8293 => x"af",
          8294 => x"2e",
          8295 => x"8e",
          8296 => x"bf",
          8297 => x"38",
          8298 => x"2e",
          8299 => x"8e",
          8300 => x"80",
          8301 => x"c2",
          8302 => x"d5",
          8303 => x"78",
          8304 => x"8c",
          8305 => x"80",
          8306 => x"38",
          8307 => x"2e",
          8308 => x"78",
          8309 => x"8b",
          8310 => x"c1",
          8311 => x"d1",
          8312 => x"38",
          8313 => x"2e",
          8314 => x"8e",
          8315 => x"81",
          8316 => x"86",
          8317 => x"82",
          8318 => x"78",
          8319 => x"8d",
          8320 => x"80",
          8321 => x"b4",
          8322 => x"39",
          8323 => x"2e",
          8324 => x"78",
          8325 => x"8d",
          8326 => x"81",
          8327 => x"ff",
          8328 => x"ff",
          8329 => x"fe",
          8330 => x"82",
          8331 => x"88",
          8332 => x"ec",
          8333 => x"39",
          8334 => x"fc",
          8335 => x"84",
          8336 => x"ed",
          8337 => x"93",
          8338 => x"2e",
          8339 => x"63",
          8340 => x"80",
          8341 => x"cb",
          8342 => x"02",
          8343 => x"33",
          8344 => x"dd",
          8345 => x"84",
          8346 => x"06",
          8347 => x"38",
          8348 => x"51",
          8349 => x"3f",
          8350 => x"a7",
          8351 => x"8c",
          8352 => x"39",
          8353 => x"80",
          8354 => x"84",
          8355 => x"ed",
          8356 => x"93",
          8357 => x"2e",
          8358 => x"80",
          8359 => x"02",
          8360 => x"33",
          8361 => x"e6",
          8362 => x"84",
          8363 => x"8a",
          8364 => x"bf",
          8365 => x"ff",
          8366 => x"ff",
          8367 => x"fe",
          8368 => x"82",
          8369 => x"80",
          8370 => x"63",
          8371 => x"d3",
          8372 => x"fe",
          8373 => x"ff",
          8374 => x"fe",
          8375 => x"82",
          8376 => x"86",
          8377 => x"84",
          8378 => x"53",
          8379 => x"52",
          8380 => x"ea",
          8381 => x"80",
          8382 => x"53",
          8383 => x"84",
          8384 => x"94",
          8385 => x"ff",
          8386 => x"82",
          8387 => x"81",
          8388 => x"89",
          8389 => x"e4",
          8390 => x"5d",
          8391 => x"b4",
          8392 => x"05",
          8393 => x"9b",
          8394 => x"84",
          8395 => x"ff",
          8396 => x"5b",
          8397 => x"3f",
          8398 => x"93",
          8399 => x"7a",
          8400 => x"3f",
          8401 => x"b4",
          8402 => x"05",
          8403 => x"f3",
          8404 => x"84",
          8405 => x"ff",
          8406 => x"5b",
          8407 => x"3f",
          8408 => x"08",
          8409 => x"84",
          8410 => x"fe",
          8411 => x"82",
          8412 => x"b5",
          8413 => x"05",
          8414 => x"cd",
          8415 => x"8e",
          8416 => x"93",
          8417 => x"56",
          8418 => x"93",
          8419 => x"ff",
          8420 => x"53",
          8421 => x"51",
          8422 => x"82",
          8423 => x"80",
          8424 => x"38",
          8425 => x"08",
          8426 => x"3f",
          8427 => x"b4",
          8428 => x"11",
          8429 => x"05",
          8430 => x"e5",
          8431 => x"84",
          8432 => x"fa",
          8433 => x"3d",
          8434 => x"53",
          8435 => x"51",
          8436 => x"3f",
          8437 => x"08",
          8438 => x"c7",
          8439 => x"fe",
          8440 => x"ff",
          8441 => x"fe",
          8442 => x"82",
          8443 => x"86",
          8444 => x"84",
          8445 => x"8a",
          8446 => x"e2",
          8447 => x"63",
          8448 => x"7b",
          8449 => x"38",
          8450 => x"7a",
          8451 => x"5c",
          8452 => x"26",
          8453 => x"e1",
          8454 => x"ff",
          8455 => x"ff",
          8456 => x"fe",
          8457 => x"82",
          8458 => x"80",
          8459 => x"38",
          8460 => x"fc",
          8461 => x"84",
          8462 => x"e9",
          8463 => x"93",
          8464 => x"2e",
          8465 => x"b4",
          8466 => x"11",
          8467 => x"05",
          8468 => x"cd",
          8469 => x"84",
          8470 => x"f9",
          8471 => x"8a",
          8472 => x"e1",
          8473 => x"5a",
          8474 => x"81",
          8475 => x"59",
          8476 => x"05",
          8477 => x"34",
          8478 => x"42",
          8479 => x"3d",
          8480 => x"53",
          8481 => x"51",
          8482 => x"3f",
          8483 => x"08",
          8484 => x"8f",
          8485 => x"fe",
          8486 => x"ff",
          8487 => x"fe",
          8488 => x"82",
          8489 => x"80",
          8490 => x"38",
          8491 => x"f8",
          8492 => x"84",
          8493 => x"e8",
          8494 => x"93",
          8495 => x"2e",
          8496 => x"82",
          8497 => x"fe",
          8498 => x"63",
          8499 => x"27",
          8500 => x"70",
          8501 => x"5e",
          8502 => x"7c",
          8503 => x"78",
          8504 => x"79",
          8505 => x"52",
          8506 => x"51",
          8507 => x"3f",
          8508 => x"81",
          8509 => x"d5",
          8510 => x"f8",
          8511 => x"39",
          8512 => x"80",
          8513 => x"84",
          8514 => x"e8",
          8515 => x"93",
          8516 => x"df",
          8517 => x"c8",
          8518 => x"80",
          8519 => x"82",
          8520 => x"44",
          8521 => x"82",
          8522 => x"59",
          8523 => x"88",
          8524 => x"88",
          8525 => x"39",
          8526 => x"33",
          8527 => x"2e",
          8528 => x"8e",
          8529 => x"ab",
          8530 => x"cb",
          8531 => x"80",
          8532 => x"82",
          8533 => x"44",
          8534 => x"8e",
          8535 => x"78",
          8536 => x"38",
          8537 => x"08",
          8538 => x"82",
          8539 => x"fc",
          8540 => x"b4",
          8541 => x"11",
          8542 => x"05",
          8543 => x"a1",
          8544 => x"84",
          8545 => x"38",
          8546 => x"33",
          8547 => x"2e",
          8548 => x"8e",
          8549 => x"80",
          8550 => x"8e",
          8551 => x"78",
          8552 => x"38",
          8553 => x"08",
          8554 => x"82",
          8555 => x"59",
          8556 => x"88",
          8557 => x"94",
          8558 => x"39",
          8559 => x"33",
          8560 => x"2e",
          8561 => x"8e",
          8562 => x"99",
          8563 => x"c6",
          8564 => x"80",
          8565 => x"82",
          8566 => x"43",
          8567 => x"8e",
          8568 => x"05",
          8569 => x"fe",
          8570 => x"ff",
          8571 => x"fe",
          8572 => x"82",
          8573 => x"80",
          8574 => x"80",
          8575 => x"7a",
          8576 => x"38",
          8577 => x"90",
          8578 => x"70",
          8579 => x"2a",
          8580 => x"51",
          8581 => x"78",
          8582 => x"38",
          8583 => x"83",
          8584 => x"82",
          8585 => x"fe",
          8586 => x"a0",
          8587 => x"61",
          8588 => x"63",
          8589 => x"3f",
          8590 => x"51",
          8591 => x"3f",
          8592 => x"b4",
          8593 => x"11",
          8594 => x"05",
          8595 => x"d1",
          8596 => x"84",
          8597 => x"f5",
          8598 => x"3d",
          8599 => x"53",
          8600 => x"51",
          8601 => x"3f",
          8602 => x"08",
          8603 => x"38",
          8604 => x"80",
          8605 => x"79",
          8606 => x"05",
          8607 => x"fe",
          8608 => x"ff",
          8609 => x"fe",
          8610 => x"82",
          8611 => x"e0",
          8612 => x"39",
          8613 => x"54",
          8614 => x"94",
          8615 => x"8c",
          8616 => x"52",
          8617 => x"e3",
          8618 => x"45",
          8619 => x"78",
          8620 => x"ef",
          8621 => x"27",
          8622 => x"3d",
          8623 => x"53",
          8624 => x"51",
          8625 => x"3f",
          8626 => x"08",
          8627 => x"38",
          8628 => x"80",
          8629 => x"79",
          8630 => x"05",
          8631 => x"39",
          8632 => x"51",
          8633 => x"3f",
          8634 => x"b4",
          8635 => x"11",
          8636 => x"05",
          8637 => x"9b",
          8638 => x"84",
          8639 => x"f4",
          8640 => x"3d",
          8641 => x"53",
          8642 => x"51",
          8643 => x"3f",
          8644 => x"08",
          8645 => x"38",
          8646 => x"be",
          8647 => x"70",
          8648 => x"23",
          8649 => x"3d",
          8650 => x"53",
          8651 => x"51",
          8652 => x"3f",
          8653 => x"08",
          8654 => x"e7",
          8655 => x"22",
          8656 => x"8b",
          8657 => x"e1",
          8658 => x"f8",
          8659 => x"fe",
          8660 => x"79",
          8661 => x"59",
          8662 => x"f3",
          8663 => x"9f",
          8664 => x"60",
          8665 => x"d5",
          8666 => x"fe",
          8667 => x"ff",
          8668 => x"fe",
          8669 => x"82",
          8670 => x"80",
          8671 => x"60",
          8672 => x"05",
          8673 => x"82",
          8674 => x"78",
          8675 => x"39",
          8676 => x"51",
          8677 => x"3f",
          8678 => x"b4",
          8679 => x"11",
          8680 => x"05",
          8681 => x"eb",
          8682 => x"84",
          8683 => x"f2",
          8684 => x"3d",
          8685 => x"53",
          8686 => x"51",
          8687 => x"3f",
          8688 => x"08",
          8689 => x"38",
          8690 => x"0c",
          8691 => x"05",
          8692 => x"fe",
          8693 => x"ff",
          8694 => x"fe",
          8695 => x"82",
          8696 => x"e4",
          8697 => x"39",
          8698 => x"54",
          8699 => x"b4",
          8700 => x"b8",
          8701 => x"52",
          8702 => x"e1",
          8703 => x"45",
          8704 => x"78",
          8705 => x"9b",
          8706 => x"27",
          8707 => x"3d",
          8708 => x"53",
          8709 => x"51",
          8710 => x"3f",
          8711 => x"08",
          8712 => x"38",
          8713 => x"0c",
          8714 => x"05",
          8715 => x"39",
          8716 => x"51",
          8717 => x"3f",
          8718 => x"82",
          8719 => x"fe",
          8720 => x"82",
          8721 => x"d7",
          8722 => x"39",
          8723 => x"51",
          8724 => x"3f",
          8725 => x"d4",
          8726 => x"c7",
          8727 => x"f0",
          8728 => x"e4",
          8729 => x"81",
          8730 => x"94",
          8731 => x"80",
          8732 => x"c0",
          8733 => x"f1",
          8734 => x"8c",
          8735 => x"d9",
          8736 => x"80",
          8737 => x"c0",
          8738 => x"8c",
          8739 => x"87",
          8740 => x"0c",
          8741 => x"b4",
          8742 => x"11",
          8743 => x"05",
          8744 => x"fd",
          8745 => x"84",
          8746 => x"f0",
          8747 => x"52",
          8748 => x"51",
          8749 => x"3f",
          8750 => x"04",
          8751 => x"80",
          8752 => x"84",
          8753 => x"e0",
          8754 => x"93",
          8755 => x"2e",
          8756 => x"63",
          8757 => x"b4",
          8758 => x"d0",
          8759 => x"78",
          8760 => x"84",
          8761 => x"f0",
          8762 => x"93",
          8763 => x"82",
          8764 => x"fe",
          8765 => x"f0",
          8766 => x"8c",
          8767 => x"d8",
          8768 => x"b8",
          8769 => x"9b",
          8770 => x"88",
          8771 => x"b8",
          8772 => x"ff",
          8773 => x"ce",
          8774 => x"87",
          8775 => x"79",
          8776 => x"80",
          8777 => x"38",
          8778 => x"59",
          8779 => x"81",
          8780 => x"3d",
          8781 => x"51",
          8782 => x"3f",
          8783 => x"08",
          8784 => x"7b",
          8785 => x"38",
          8786 => x"89",
          8787 => x"2e",
          8788 => x"cd",
          8789 => x"2e",
          8790 => x"c5",
          8791 => x"9c",
          8792 => x"82",
          8793 => x"80",
          8794 => x"a4",
          8795 => x"ff",
          8796 => x"fe",
          8797 => x"bb",
          8798 => x"c4",
          8799 => x"ff",
          8800 => x"fe",
          8801 => x"ab",
          8802 => x"82",
          8803 => x"80",
          8804 => x"b4",
          8805 => x"ff",
          8806 => x"fe",
          8807 => x"93",
          8808 => x"80",
          8809 => x"c0",
          8810 => x"ff",
          8811 => x"fe",
          8812 => x"82",
          8813 => x"82",
          8814 => x"80",
          8815 => x"80",
          8816 => x"80",
          8817 => x"80",
          8818 => x"ff",
          8819 => x"e6",
          8820 => x"93",
          8821 => x"93",
          8822 => x"70",
          8823 => x"07",
          8824 => x"5b",
          8825 => x"5a",
          8826 => x"83",
          8827 => x"78",
          8828 => x"78",
          8829 => x"38",
          8830 => x"81",
          8831 => x"59",
          8832 => x"38",
          8833 => x"7d",
          8834 => x"59",
          8835 => x"7e",
          8836 => x"81",
          8837 => x"38",
          8838 => x"51",
          8839 => x"3f",
          8840 => x"fc",
          8841 => x"0b",
          8842 => x"34",
          8843 => x"8c",
          8844 => x"55",
          8845 => x"52",
          8846 => x"b6",
          8847 => x"93",
          8848 => x"2b",
          8849 => x"53",
          8850 => x"52",
          8851 => x"b6",
          8852 => x"82",
          8853 => x"07",
          8854 => x"c0",
          8855 => x"08",
          8856 => x"84",
          8857 => x"51",
          8858 => x"3f",
          8859 => x"08",
          8860 => x"08",
          8861 => x"84",
          8862 => x"51",
          8863 => x"3f",
          8864 => x"84",
          8865 => x"0c",
          8866 => x"0b",
          8867 => x"84",
          8868 => x"83",
          8869 => x"94",
          8870 => x"ac",
          8871 => x"98",
          8872 => x"0b",
          8873 => x"0c",
          8874 => x"3f",
          8875 => x"3f",
          8876 => x"51",
          8877 => x"3f",
          8878 => x"51",
          8879 => x"3f",
          8880 => x"51",
          8881 => x"3f",
          8882 => x"fc",
          8883 => x"3f",
          8884 => x"00",
          8885 => x"55",
          8886 => x"5b",
          8887 => x"61",
          8888 => x"67",
          8889 => x"6d",
          8890 => x"19",
          8891 => x"f5",
          8892 => x"98",
          8893 => x"d8",
          8894 => x"fb",
          8895 => x"88",
          8896 => x"ee",
          8897 => x"ee",
          8898 => x"c5",
          8899 => x"3b",
          8900 => x"c6",
          8901 => x"ef",
          8902 => x"0d",
          8903 => x"91",
          8904 => x"98",
          8905 => x"9f",
          8906 => x"a6",
          8907 => x"ad",
          8908 => x"b4",
          8909 => x"bb",
          8910 => x"c2",
          8911 => x"c9",
          8912 => x"d0",
          8913 => x"d7",
          8914 => x"dd",
          8915 => x"e3",
          8916 => x"e9",
          8917 => x"ef",
          8918 => x"f5",
          8919 => x"fb",
          8920 => x"01",
          8921 => x"07",
          8922 => x"25",
          8923 => x"64",
          8924 => x"3a",
          8925 => x"25",
          8926 => x"64",
          8927 => x"00",
          8928 => x"20",
          8929 => x"66",
          8930 => x"72",
          8931 => x"6f",
          8932 => x"00",
          8933 => x"72",
          8934 => x"53",
          8935 => x"63",
          8936 => x"69",
          8937 => x"00",
          8938 => x"65",
          8939 => x"65",
          8940 => x"6d",
          8941 => x"6d",
          8942 => x"65",
          8943 => x"00",
          8944 => x"20",
          8945 => x"53",
          8946 => x"4d",
          8947 => x"25",
          8948 => x"3a",
          8949 => x"58",
          8950 => x"00",
          8951 => x"20",
          8952 => x"41",
          8953 => x"20",
          8954 => x"25",
          8955 => x"3a",
          8956 => x"58",
          8957 => x"00",
          8958 => x"20",
          8959 => x"4e",
          8960 => x"41",
          8961 => x"25",
          8962 => x"3a",
          8963 => x"58",
          8964 => x"00",
          8965 => x"20",
          8966 => x"4d",
          8967 => x"20",
          8968 => x"25",
          8969 => x"3a",
          8970 => x"58",
          8971 => x"00",
          8972 => x"20",
          8973 => x"20",
          8974 => x"20",
          8975 => x"25",
          8976 => x"3a",
          8977 => x"58",
          8978 => x"00",
          8979 => x"20",
          8980 => x"43",
          8981 => x"20",
          8982 => x"44",
          8983 => x"63",
          8984 => x"3d",
          8985 => x"64",
          8986 => x"00",
          8987 => x"20",
          8988 => x"45",
          8989 => x"20",
          8990 => x"54",
          8991 => x"72",
          8992 => x"3d",
          8993 => x"64",
          8994 => x"00",
          8995 => x"20",
          8996 => x"52",
          8997 => x"52",
          8998 => x"43",
          8999 => x"6e",
          9000 => x"3d",
          9001 => x"64",
          9002 => x"00",
          9003 => x"20",
          9004 => x"48",
          9005 => x"45",
          9006 => x"53",
          9007 => x"00",
          9008 => x"20",
          9009 => x"49",
          9010 => x"00",
          9011 => x"20",
          9012 => x"54",
          9013 => x"00",
          9014 => x"20",
          9015 => x"0a",
          9016 => x"00",
          9017 => x"20",
          9018 => x"0a",
          9019 => x"00",
          9020 => x"72",
          9021 => x"65",
          9022 => x"00",
          9023 => x"20",
          9024 => x"20",
          9025 => x"65",
          9026 => x"65",
          9027 => x"72",
          9028 => x"64",
          9029 => x"73",
          9030 => x"25",
          9031 => x"0a",
          9032 => x"00",
          9033 => x"20",
          9034 => x"20",
          9035 => x"6f",
          9036 => x"53",
          9037 => x"74",
          9038 => x"64",
          9039 => x"73",
          9040 => x"25",
          9041 => x"0a",
          9042 => x"00",
          9043 => x"20",
          9044 => x"63",
          9045 => x"74",
          9046 => x"20",
          9047 => x"72",
          9048 => x"20",
          9049 => x"20",
          9050 => x"25",
          9051 => x"0a",
          9052 => x"00",
          9053 => x"63",
          9054 => x"00",
          9055 => x"20",
          9056 => x"20",
          9057 => x"20",
          9058 => x"20",
          9059 => x"20",
          9060 => x"20",
          9061 => x"20",
          9062 => x"25",
          9063 => x"0a",
          9064 => x"00",
          9065 => x"20",
          9066 => x"74",
          9067 => x"43",
          9068 => x"6b",
          9069 => x"65",
          9070 => x"20",
          9071 => x"20",
          9072 => x"25",
          9073 => x"30",
          9074 => x"48",
          9075 => x"00",
          9076 => x"20",
          9077 => x"41",
          9078 => x"6c",
          9079 => x"20",
          9080 => x"71",
          9081 => x"20",
          9082 => x"20",
          9083 => x"25",
          9084 => x"30",
          9085 => x"48",
          9086 => x"00",
          9087 => x"20",
          9088 => x"68",
          9089 => x"65",
          9090 => x"52",
          9091 => x"43",
          9092 => x"6b",
          9093 => x"65",
          9094 => x"25",
          9095 => x"30",
          9096 => x"48",
          9097 => x"00",
          9098 => x"6c",
          9099 => x"00",
          9100 => x"69",
          9101 => x"00",
          9102 => x"78",
          9103 => x"00",
          9104 => x"00",
          9105 => x"6d",
          9106 => x"00",
          9107 => x"6e",
          9108 => x"00",
          9109 => x"74",
          9110 => x"2e",
          9111 => x"00",
          9112 => x"74",
          9113 => x"00",
          9114 => x"74",
          9115 => x"00",
          9116 => x"00",
          9117 => x"64",
          9118 => x"73",
          9119 => x"00",
          9120 => x"6c",
          9121 => x"74",
          9122 => x"65",
          9123 => x"20",
          9124 => x"20",
          9125 => x"74",
          9126 => x"20",
          9127 => x"65",
          9128 => x"20",
          9129 => x"2e",
          9130 => x"00",
          9131 => x"6e",
          9132 => x"6f",
          9133 => x"2f",
          9134 => x"61",
          9135 => x"68",
          9136 => x"6f",
          9137 => x"66",
          9138 => x"2c",
          9139 => x"73",
          9140 => x"69",
          9141 => x"0a",
          9142 => x"00",
          9143 => x"88",
          9144 => x"00",
          9145 => x"01",
          9146 => x"84",
          9147 => x"00",
          9148 => x"02",
          9149 => x"80",
          9150 => x"00",
          9151 => x"03",
          9152 => x"7c",
          9153 => x"00",
          9154 => x"04",
          9155 => x"78",
          9156 => x"00",
          9157 => x"05",
          9158 => x"74",
          9159 => x"00",
          9160 => x"06",
          9161 => x"70",
          9162 => x"00",
          9163 => x"07",
          9164 => x"6c",
          9165 => x"00",
          9166 => x"08",
          9167 => x"68",
          9168 => x"00",
          9169 => x"09",
          9170 => x"64",
          9171 => x"00",
          9172 => x"0a",
          9173 => x"60",
          9174 => x"00",
          9175 => x"0b",
          9176 => x"00",
          9177 => x"00",
          9178 => x"00",
          9179 => x"00",
          9180 => x"7e",
          9181 => x"7e",
          9182 => x"7e",
          9183 => x"7e",
          9184 => x"7e",
          9185 => x"00",
          9186 => x"00",
          9187 => x"00",
          9188 => x"2c",
          9189 => x"3d",
          9190 => x"5d",
          9191 => x"00",
          9192 => x"00",
          9193 => x"33",
          9194 => x"00",
          9195 => x"4d",
          9196 => x"53",
          9197 => x"00",
          9198 => x"4e",
          9199 => x"20",
          9200 => x"46",
          9201 => x"32",
          9202 => x"00",
          9203 => x"4e",
          9204 => x"20",
          9205 => x"46",
          9206 => x"20",
          9207 => x"00",
          9208 => x"8c",
          9209 => x"00",
          9210 => x"00",
          9211 => x"00",
          9212 => x"41",
          9213 => x"80",
          9214 => x"49",
          9215 => x"8f",
          9216 => x"4f",
          9217 => x"55",
          9218 => x"9b",
          9219 => x"9f",
          9220 => x"55",
          9221 => x"a7",
          9222 => x"ab",
          9223 => x"af",
          9224 => x"b3",
          9225 => x"b7",
          9226 => x"bb",
          9227 => x"bf",
          9228 => x"c3",
          9229 => x"c7",
          9230 => x"cb",
          9231 => x"cf",
          9232 => x"d3",
          9233 => x"d7",
          9234 => x"db",
          9235 => x"df",
          9236 => x"e3",
          9237 => x"e7",
          9238 => x"eb",
          9239 => x"ef",
          9240 => x"f3",
          9241 => x"f7",
          9242 => x"fb",
          9243 => x"ff",
          9244 => x"3b",
          9245 => x"2f",
          9246 => x"3a",
          9247 => x"7c",
          9248 => x"00",
          9249 => x"04",
          9250 => x"40",
          9251 => x"00",
          9252 => x"00",
          9253 => x"02",
          9254 => x"08",
          9255 => x"20",
          9256 => x"00",
          9257 => x"69",
          9258 => x"00",
          9259 => x"63",
          9260 => x"00",
          9261 => x"69",
          9262 => x"00",
          9263 => x"61",
          9264 => x"00",
          9265 => x"65",
          9266 => x"00",
          9267 => x"65",
          9268 => x"00",
          9269 => x"70",
          9270 => x"00",
          9271 => x"66",
          9272 => x"00",
          9273 => x"6d",
          9274 => x"00",
          9275 => x"00",
          9276 => x"00",
          9277 => x"00",
          9278 => x"00",
          9279 => x"00",
          9280 => x"00",
          9281 => x"00",
          9282 => x"6c",
          9283 => x"00",
          9284 => x"00",
          9285 => x"74",
          9286 => x"00",
          9287 => x"65",
          9288 => x"00",
          9289 => x"6f",
          9290 => x"00",
          9291 => x"74",
          9292 => x"00",
          9293 => x"73",
          9294 => x"00",
          9295 => x"73",
          9296 => x"00",
          9297 => x"6f",
          9298 => x"00",
          9299 => x"6b",
          9300 => x"72",
          9301 => x"00",
          9302 => x"65",
          9303 => x"6c",
          9304 => x"72",
          9305 => x"0a",
          9306 => x"00",
          9307 => x"6b",
          9308 => x"74",
          9309 => x"61",
          9310 => x"0a",
          9311 => x"00",
          9312 => x"66",
          9313 => x"20",
          9314 => x"6e",
          9315 => x"00",
          9316 => x"70",
          9317 => x"20",
          9318 => x"6e",
          9319 => x"00",
          9320 => x"61",
          9321 => x"20",
          9322 => x"65",
          9323 => x"65",
          9324 => x"00",
          9325 => x"65",
          9326 => x"64",
          9327 => x"65",
          9328 => x"00",
          9329 => x"65",
          9330 => x"72",
          9331 => x"79",
          9332 => x"69",
          9333 => x"2e",
          9334 => x"00",
          9335 => x"65",
          9336 => x"6e",
          9337 => x"20",
          9338 => x"61",
          9339 => x"2e",
          9340 => x"00",
          9341 => x"69",
          9342 => x"72",
          9343 => x"20",
          9344 => x"74",
          9345 => x"65",
          9346 => x"00",
          9347 => x"76",
          9348 => x"75",
          9349 => x"72",
          9350 => x"20",
          9351 => x"61",
          9352 => x"2e",
          9353 => x"00",
          9354 => x"6b",
          9355 => x"74",
          9356 => x"61",
          9357 => x"64",
          9358 => x"00",
          9359 => x"63",
          9360 => x"61",
          9361 => x"6c",
          9362 => x"69",
          9363 => x"79",
          9364 => x"6d",
          9365 => x"75",
          9366 => x"6f",
          9367 => x"69",
          9368 => x"0a",
          9369 => x"00",
          9370 => x"6d",
          9371 => x"61",
          9372 => x"74",
          9373 => x"0a",
          9374 => x"00",
          9375 => x"65",
          9376 => x"2c",
          9377 => x"65",
          9378 => x"69",
          9379 => x"63",
          9380 => x"65",
          9381 => x"64",
          9382 => x"00",
          9383 => x"65",
          9384 => x"20",
          9385 => x"6b",
          9386 => x"0a",
          9387 => x"00",
          9388 => x"75",
          9389 => x"63",
          9390 => x"74",
          9391 => x"6d",
          9392 => x"2e",
          9393 => x"00",
          9394 => x"20",
          9395 => x"79",
          9396 => x"65",
          9397 => x"69",
          9398 => x"2e",
          9399 => x"00",
          9400 => x"61",
          9401 => x"65",
          9402 => x"69",
          9403 => x"72",
          9404 => x"74",
          9405 => x"00",
          9406 => x"63",
          9407 => x"2e",
          9408 => x"00",
          9409 => x"6e",
          9410 => x"20",
          9411 => x"6f",
          9412 => x"00",
          9413 => x"75",
          9414 => x"74",
          9415 => x"25",
          9416 => x"74",
          9417 => x"75",
          9418 => x"74",
          9419 => x"73",
          9420 => x"0a",
          9421 => x"00",
          9422 => x"64",
          9423 => x"00",
          9424 => x"58",
          9425 => x"00",
          9426 => x"00",
          9427 => x"58",
          9428 => x"00",
          9429 => x"20",
          9430 => x"20",
          9431 => x"00",
          9432 => x"58",
          9433 => x"00",
          9434 => x"00",
          9435 => x"00",
          9436 => x"00",
          9437 => x"54",
          9438 => x"00",
          9439 => x"20",
          9440 => x"28",
          9441 => x"00",
          9442 => x"30",
          9443 => x"30",
          9444 => x"00",
          9445 => x"35",
          9446 => x"00",
          9447 => x"55",
          9448 => x"65",
          9449 => x"30",
          9450 => x"20",
          9451 => x"25",
          9452 => x"2a",
          9453 => x"00",
          9454 => x"54",
          9455 => x"6e",
          9456 => x"72",
          9457 => x"20",
          9458 => x"64",
          9459 => x"0a",
          9460 => x"00",
          9461 => x"65",
          9462 => x"6e",
          9463 => x"72",
          9464 => x"0a",
          9465 => x"00",
          9466 => x"20",
          9467 => x"65",
          9468 => x"70",
          9469 => x"00",
          9470 => x"54",
          9471 => x"44",
          9472 => x"74",
          9473 => x"75",
          9474 => x"00",
          9475 => x"54",
          9476 => x"52",
          9477 => x"74",
          9478 => x"75",
          9479 => x"00",
          9480 => x"54",
          9481 => x"58",
          9482 => x"74",
          9483 => x"75",
          9484 => x"00",
          9485 => x"54",
          9486 => x"58",
          9487 => x"74",
          9488 => x"75",
          9489 => x"00",
          9490 => x"54",
          9491 => x"58",
          9492 => x"74",
          9493 => x"75",
          9494 => x"00",
          9495 => x"54",
          9496 => x"58",
          9497 => x"74",
          9498 => x"75",
          9499 => x"00",
          9500 => x"74",
          9501 => x"20",
          9502 => x"74",
          9503 => x"72",
          9504 => x"0a",
          9505 => x"00",
          9506 => x"62",
          9507 => x"67",
          9508 => x"6d",
          9509 => x"2e",
          9510 => x"00",
          9511 => x"6f",
          9512 => x"63",
          9513 => x"74",
          9514 => x"00",
          9515 => x"00",
          9516 => x"6c",
          9517 => x"74",
          9518 => x"6e",
          9519 => x"61",
          9520 => x"65",
          9521 => x"20",
          9522 => x"64",
          9523 => x"20",
          9524 => x"61",
          9525 => x"69",
          9526 => x"20",
          9527 => x"75",
          9528 => x"79",
          9529 => x"00",
          9530 => x"00",
          9531 => x"20",
          9532 => x"6b",
          9533 => x"21",
          9534 => x"00",
          9535 => x"74",
          9536 => x"69",
          9537 => x"2e",
          9538 => x"00",
          9539 => x"6c",
          9540 => x"74",
          9541 => x"6e",
          9542 => x"61",
          9543 => x"65",
          9544 => x"00",
          9545 => x"25",
          9546 => x"00",
          9547 => x"00",
          9548 => x"61",
          9549 => x"67",
          9550 => x"2e",
          9551 => x"00",
          9552 => x"79",
          9553 => x"2e",
          9554 => x"00",
          9555 => x"70",
          9556 => x"6e",
          9557 => x"2e",
          9558 => x"00",
          9559 => x"6c",
          9560 => x"30",
          9561 => x"2d",
          9562 => x"38",
          9563 => x"25",
          9564 => x"29",
          9565 => x"00",
          9566 => x"70",
          9567 => x"6d",
          9568 => x"0a",
          9569 => x"00",
          9570 => x"6d",
          9571 => x"74",
          9572 => x"00",
          9573 => x"58",
          9574 => x"32",
          9575 => x"00",
          9576 => x"0a",
          9577 => x"00",
          9578 => x"58",
          9579 => x"34",
          9580 => x"00",
          9581 => x"58",
          9582 => x"38",
          9583 => x"00",
          9584 => x"61",
          9585 => x"6e",
          9586 => x"6e",
          9587 => x"72",
          9588 => x"73",
          9589 => x"00",
          9590 => x"62",
          9591 => x"67",
          9592 => x"74",
          9593 => x"75",
          9594 => x"0a",
          9595 => x"00",
          9596 => x"61",
          9597 => x"64",
          9598 => x"72",
          9599 => x"69",
          9600 => x"00",
          9601 => x"62",
          9602 => x"67",
          9603 => x"72",
          9604 => x"69",
          9605 => x"00",
          9606 => x"63",
          9607 => x"6e",
          9608 => x"6f",
          9609 => x"40",
          9610 => x"38",
          9611 => x"2e",
          9612 => x"00",
          9613 => x"6c",
          9614 => x"20",
          9615 => x"65",
          9616 => x"25",
          9617 => x"20",
          9618 => x"0a",
          9619 => x"00",
          9620 => x"6c",
          9621 => x"74",
          9622 => x"65",
          9623 => x"6f",
          9624 => x"28",
          9625 => x"2e",
          9626 => x"00",
          9627 => x"74",
          9628 => x"69",
          9629 => x"61",
          9630 => x"69",
          9631 => x"69",
          9632 => x"2e",
          9633 => x"00",
          9634 => x"64",
          9635 => x"62",
          9636 => x"69",
          9637 => x"2e",
          9638 => x"00",
          9639 => x"00",
          9640 => x"00",
          9641 => x"5c",
          9642 => x"25",
          9643 => x"73",
          9644 => x"00",
          9645 => x"5c",
          9646 => x"25",
          9647 => x"00",
          9648 => x"5c",
          9649 => x"00",
          9650 => x"20",
          9651 => x"6d",
          9652 => x"2e",
          9653 => x"00",
          9654 => x"6e",
          9655 => x"2e",
          9656 => x"00",
          9657 => x"62",
          9658 => x"67",
          9659 => x"74",
          9660 => x"75",
          9661 => x"2e",
          9662 => x"00",
          9663 => x"00",
          9664 => x"00",
          9665 => x"ff",
          9666 => x"00",
          9667 => x"ff",
          9668 => x"00",
          9669 => x"ff",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"ff",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"00",
          9679 => x"00",
          9680 => x"00",
          9681 => x"00",
          9682 => x"01",
          9683 => x"01",
          9684 => x"01",
          9685 => x"00",
          9686 => x"00",
          9687 => x"02",
          9688 => x"00",
          9689 => x"5c",
          9690 => x"5c",
          9691 => x"5c",
          9692 => x"5c",
          9693 => x"54",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"60",
          9718 => x"00",
          9719 => x"68",
          9720 => x"00",
          9721 => x"70",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"a4",
          9726 => x"00",
          9727 => x"00",
          9728 => x"00",
          9729 => x"ac",
          9730 => x"00",
          9731 => x"00",
          9732 => x"00",
          9733 => x"b4",
          9734 => x"00",
          9735 => x"00",
          9736 => x"00",
          9737 => x"bc",
          9738 => x"00",
          9739 => x"00",
          9740 => x"00",
          9741 => x"c4",
          9742 => x"00",
          9743 => x"00",
          9744 => x"00",
          9745 => x"cc",
          9746 => x"00",
          9747 => x"00",
          9748 => x"00",
          9749 => x"d4",
          9750 => x"00",
          9751 => x"00",
          9752 => x"00",
          9753 => x"dc",
          9754 => x"00",
          9755 => x"00",
          9756 => x"00",
          9757 => x"e4",
          9758 => x"00",
          9759 => x"00",
          9760 => x"00",
          9761 => x"ec",
          9762 => x"00",
          9763 => x"00",
          9764 => x"00",
          9765 => x"f0",
          9766 => x"00",
          9767 => x"00",
          9768 => x"00",
          9769 => x"f4",
          9770 => x"00",
          9771 => x"00",
          9772 => x"00",
          9773 => x"f8",
          9774 => x"00",
          9775 => x"00",
          9776 => x"00",
          9777 => x"fc",
          9778 => x"00",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"00",
          9783 => x"00",
          9784 => x"00",
          9785 => x"04",
          9786 => x"00",
          9787 => x"00",
          9788 => x"00",
          9789 => x"08",
          9790 => x"00",
          9791 => x"00",
          9792 => x"00",
          9793 => x"10",
          9794 => x"00",
          9795 => x"00",
          9796 => x"00",
          9797 => x"14",
          9798 => x"00",
          9799 => x"00",
          9800 => x"00",
          9801 => x"1c",
          9802 => x"00",
          9803 => x"00",
          9804 => x"00",
          9805 => x"24",
          9806 => x"00",
          9807 => x"00",
          9808 => x"00",
          9809 => x"2c",
          9810 => x"00",
          9811 => x"00",
          9812 => x"00",
          9813 => x"34",
          9814 => x"00",
          9815 => x"00",
          9816 => x"00",
          9817 => x"3c",
          9818 => x"00",
          9819 => x"00",
          9820 => x"00",
          9821 => x"44",
          9822 => x"00",
          9823 => x"00",
          9824 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"0b",
             1 => x"00",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"8c",
             9 => x"0b",
            10 => x"80",
            11 => x"0c",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"06",
            17 => x"06",
            18 => x"82",
            19 => x"2a",
            20 => x"06",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"06",
            25 => x"ff",
            26 => x"09",
            27 => x"05",
            28 => x"09",
            29 => x"ff",
            30 => x"0b",
            31 => x"04",
            32 => x"81",
            33 => x"73",
            34 => x"09",
            35 => x"73",
            36 => x"81",
            37 => x"04",
            38 => x"00",
            39 => x"00",
            40 => x"24",
            41 => x"07",
            42 => x"00",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"81",
            50 => x"05",
            51 => x"0a",
            52 => x"0a",
            53 => x"81",
            54 => x"53",
            55 => x"00",
            56 => x"26",
            57 => x"07",
            58 => x"00",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"00",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"51",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"9f",
            89 => x"05",
            90 => x"88",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"2a",
            97 => x"06",
            98 => x"09",
            99 => x"ff",
           100 => x"53",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"53",
           105 => x"73",
           106 => x"81",
           107 => x"83",
           108 => x"07",
           109 => x"0c",
           110 => x"00",
           111 => x"00",
           112 => x"81",
           113 => x"09",
           114 => x"09",
           115 => x"06",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"81",
           121 => x"09",
           122 => x"09",
           123 => x"81",
           124 => x"04",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"81",
           129 => x"00",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"09",
           137 => x"53",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"09",
           146 => x"51",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"06",
           153 => x"06",
           154 => x"83",
           155 => x"10",
           156 => x"06",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"06",
           161 => x"0b",
           162 => x"83",
           163 => x"05",
           164 => x"0b",
           165 => x"04",
           166 => x"00",
           167 => x"00",
           168 => x"8c",
           169 => x"75",
           170 => x"0b",
           171 => x"50",
           172 => x"56",
           173 => x"0c",
           174 => x"04",
           175 => x"00",
           176 => x"8c",
           177 => x"75",
           178 => x"0b",
           179 => x"50",
           180 => x"56",
           181 => x"0c",
           182 => x"04",
           183 => x"00",
           184 => x"70",
           185 => x"06",
           186 => x"ff",
           187 => x"71",
           188 => x"72",
           189 => x"05",
           190 => x"51",
           191 => x"00",
           192 => x"70",
           193 => x"06",
           194 => x"06",
           195 => x"54",
           196 => x"09",
           197 => x"ff",
           198 => x"51",
           199 => x"00",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"05",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"05",
           233 => x"05",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"05",
           249 => x"53",
           250 => x"04",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"04",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"00",
           267 => x"ff",
           268 => x"06",
           269 => x"83",
           270 => x"10",
           271 => x"fc",
           272 => x"51",
           273 => x"80",
           274 => x"ff",
           275 => x"06",
           276 => x"52",
           277 => x"0a",
           278 => x"38",
           279 => x"51",
           280 => x"70",
           281 => x"8e",
           282 => x"70",
           283 => x"0c",
           284 => x"88",
           285 => x"fe",
           286 => x"04",
           287 => x"00",
           288 => x"00",
           289 => x"08",
           290 => x"fd",
           291 => x"53",
           292 => x"05",
           293 => x"08",
           294 => x"51",
           295 => x"88",
           296 => x"0c",
           297 => x"0d",
           298 => x"94",
           299 => x"0c",
           300 => x"81",
           301 => x"8c",
           302 => x"94",
           303 => x"08",
           304 => x"3f",
           305 => x"88",
           306 => x"3d",
           307 => x"04",
           308 => x"94",
           309 => x"0d",
           310 => x"08",
           311 => x"94",
           312 => x"08",
           313 => x"38",
           314 => x"05",
           315 => x"08",
           316 => x"80",
           317 => x"f4",
           318 => x"08",
           319 => x"88",
           320 => x"94",
           321 => x"0c",
           322 => x"05",
           323 => x"fc",
           324 => x"08",
           325 => x"80",
           326 => x"94",
           327 => x"08",
           328 => x"8c",
           329 => x"0b",
           330 => x"05",
           331 => x"fc",
           332 => x"38",
           333 => x"08",
           334 => x"94",
           335 => x"08",
           336 => x"05",
           337 => x"94",
           338 => x"08",
           339 => x"88",
           340 => x"81",
           341 => x"08",
           342 => x"f8",
           343 => x"94",
           344 => x"08",
           345 => x"38",
           346 => x"05",
           347 => x"08",
           348 => x"94",
           349 => x"08",
           350 => x"54",
           351 => x"94",
           352 => x"08",
           353 => x"fb",
           354 => x"0b",
           355 => x"05",
           356 => x"88",
           357 => x"25",
           358 => x"08",
           359 => x"30",
           360 => x"05",
           361 => x"94",
           362 => x"0c",
           363 => x"05",
           364 => x"8c",
           365 => x"8c",
           366 => x"94",
           367 => x"0c",
           368 => x"08",
           369 => x"52",
           370 => x"05",
           371 => x"3f",
           372 => x"94",
           373 => x"0c",
           374 => x"fc",
           375 => x"2e",
           376 => x"08",
           377 => x"30",
           378 => x"05",
           379 => x"f8",
           380 => x"88",
           381 => x"3d",
           382 => x"04",
           383 => x"94",
           384 => x"0d",
           385 => x"08",
           386 => x"80",
           387 => x"f8",
           388 => x"08",
           389 => x"94",
           390 => x"08",
           391 => x"94",
           392 => x"08",
           393 => x"38",
           394 => x"08",
           395 => x"24",
           396 => x"08",
           397 => x"10",
           398 => x"05",
           399 => x"fc",
           400 => x"94",
           401 => x"0c",
           402 => x"08",
           403 => x"80",
           404 => x"38",
           405 => x"05",
           406 => x"88",
           407 => x"a1",
           408 => x"88",
           409 => x"08",
           410 => x"31",
           411 => x"05",
           412 => x"f8",
           413 => x"08",
           414 => x"07",
           415 => x"05",
           416 => x"fc",
           417 => x"2a",
           418 => x"05",
           419 => x"8c",
           420 => x"2a",
           421 => x"05",
           422 => x"39",
           423 => x"05",
           424 => x"8f",
           425 => x"88",
           426 => x"94",
           427 => x"0c",
           428 => x"94",
           429 => x"08",
           430 => x"f4",
           431 => x"94",
           432 => x"08",
           433 => x"3d",
           434 => x"04",
           435 => x"81",
           436 => x"c0",
           437 => x"81",
           438 => x"92",
           439 => x"0b",
           440 => x"8c",
           441 => x"92",
           442 => x"82",
           443 => x"70",
           444 => x"38",
           445 => x"8c",
           446 => x"e9",
           447 => x"92",
           448 => x"80",
           449 => x"71",
           450 => x"c0",
           451 => x"51",
           452 => x"88",
           453 => x"0b",
           454 => x"34",
           455 => x"9f",
           456 => x"0c",
           457 => x"04",
           458 => x"78",
           459 => x"58",
           460 => x"0b",
           461 => x"f0",
           462 => x"52",
           463 => x"70",
           464 => x"81",
           465 => x"38",
           466 => x"c0",
           467 => x"79",
           468 => x"80",
           469 => x"87",
           470 => x"0c",
           471 => x"8c",
           472 => x"2a",
           473 => x"51",
           474 => x"80",
           475 => x"87",
           476 => x"08",
           477 => x"06",
           478 => x"52",
           479 => x"80",
           480 => x"70",
           481 => x"38",
           482 => x"81",
           483 => x"ff",
           484 => x"15",
           485 => x"06",
           486 => x"2e",
           487 => x"c0",
           488 => x"51",
           489 => x"38",
           490 => x"8c",
           491 => x"95",
           492 => x"87",
           493 => x"0c",
           494 => x"8c",
           495 => x"06",
           496 => x"f4",
           497 => x"fc",
           498 => x"52",
           499 => x"2e",
           500 => x"8f",
           501 => x"98",
           502 => x"70",
           503 => x"81",
           504 => x"81",
           505 => x"0c",
           506 => x"04",
           507 => x"74",
           508 => x"71",
           509 => x"2b",
           510 => x"53",
           511 => x"0d",
           512 => x"0d",
           513 => x"33",
           514 => x"71",
           515 => x"88",
           516 => x"14",
           517 => x"07",
           518 => x"33",
           519 => x"0c",
           520 => x"56",
           521 => x"3d",
           522 => x"3d",
           523 => x"0b",
           524 => x"08",
           525 => x"77",
           526 => x"38",
           527 => x"08",
           528 => x"38",
           529 => x"74",
           530 => x"38",
           531 => x"ae",
           532 => x"39",
           533 => x"10",
           534 => x"53",
           535 => x"8c",
           536 => x"52",
           537 => x"52",
           538 => x"3f",
           539 => x"38",
           540 => x"f8",
           541 => x"83",
           542 => x"55",
           543 => x"54",
           544 => x"83",
           545 => x"76",
           546 => x"17",
           547 => x"88",
           548 => x"55",
           549 => x"88",
           550 => x"74",
           551 => x"3f",
           552 => x"0a",
           553 => x"39",
           554 => x"88",
           555 => x"0d",
           556 => x"0d",
           557 => x"9f",
           558 => x"19",
           559 => x"fe",
           560 => x"54",
           561 => x"73",
           562 => x"82",
           563 => x"71",
           564 => x"08",
           565 => x"75",
           566 => x"3d",
           567 => x"3d",
           568 => x"80",
           569 => x"0b",
           570 => x"70",
           571 => x"53",
           572 => x"09",
           573 => x"38",
           574 => x"fd",
           575 => x"08",
           576 => x"9a",
           577 => x"e4",
           578 => x"83",
           579 => x"73",
           580 => x"85",
           581 => x"fc",
           582 => x"0b",
           583 => x"f4",
           584 => x"80",
           585 => x"15",
           586 => x"81",
           587 => x"88",
           588 => x"26",
           589 => x"52",
           590 => x"90",
           591 => x"52",
           592 => x"09",
           593 => x"38",
           594 => x"53",
           595 => x"0c",
           596 => x"8b",
           597 => x"fe",
           598 => x"08",
           599 => x"90",
           600 => x"71",
           601 => x"80",
           602 => x"0c",
           603 => x"04",
           604 => x"78",
           605 => x"9f",
           606 => x"22",
           607 => x"83",
           608 => x"57",
           609 => x"73",
           610 => x"38",
           611 => x"53",
           612 => x"83",
           613 => x"39",
           614 => x"52",
           615 => x"38",
           616 => x"16",
           617 => x"08",
           618 => x"38",
           619 => x"17",
           620 => x"73",
           621 => x"38",
           622 => x"16",
           623 => x"74",
           624 => x"52",
           625 => x"72",
           626 => x"3f",
           627 => x"88",
           628 => x"38",
           629 => x"08",
           630 => x"27",
           631 => x"08",
           632 => x"88",
           633 => x"c9",
           634 => x"90",
           635 => x"75",
           636 => x"71",
           637 => x"3d",
           638 => x"3d",
           639 => x"64",
           640 => x"75",
           641 => x"a0",
           642 => x"06",
           643 => x"16",
           644 => x"ef",
           645 => x"33",
           646 => x"af",
           647 => x"06",
           648 => x"16",
           649 => x"88",
           650 => x"70",
           651 => x"74",
           652 => x"38",
           653 => x"df",
           654 => x"56",
           655 => x"82",
           656 => x"3d",
           657 => x"70",
           658 => x"8a",
           659 => x"70",
           660 => x"34",
           661 => x"74",
           662 => x"81",
           663 => x"80",
           664 => x"88",
           665 => x"5a",
           666 => x"70",
           667 => x"60",
           668 => x"70",
           669 => x"30",
           670 => x"71",
           671 => x"51",
           672 => x"53",
           673 => x"74",
           674 => x"76",
           675 => x"81",
           676 => x"81",
           677 => x"27",
           678 => x"74",
           679 => x"38",
           680 => x"70",
           681 => x"32",
           682 => x"73",
           683 => x"53",
           684 => x"56",
           685 => x"88",
           686 => x"ff",
           687 => x"81",
           688 => x"ff",
           689 => x"53",
           690 => x"76",
           691 => x"98",
           692 => x"7f",
           693 => x"76",
           694 => x"38",
           695 => x"8b",
           696 => x"51",
           697 => x"88",
           698 => x"38",
           699 => x"22",
           700 => x"83",
           701 => x"55",
           702 => x"52",
           703 => x"a8",
           704 => x"57",
           705 => x"fb",
           706 => x"55",
           707 => x"80",
           708 => x"1d",
           709 => x"2a",
           710 => x"51",
           711 => x"b2",
           712 => x"84",
           713 => x"08",
           714 => x"58",
           715 => x"77",
           716 => x"38",
           717 => x"05",
           718 => x"70",
           719 => x"33",
           720 => x"52",
           721 => x"80",
           722 => x"86",
           723 => x"2e",
           724 => x"51",
           725 => x"ff",
           726 => x"08",
           727 => x"b4",
           728 => x"76",
           729 => x"08",
           730 => x"51",
           731 => x"38",
           732 => x"70",
           733 => x"81",
           734 => x"56",
           735 => x"83",
           736 => x"81",
           737 => x"7c",
           738 => x"3f",
           739 => x"1d",
           740 => x"39",
           741 => x"90",
           742 => x"f9",
           743 => x"7b",
           744 => x"54",
           745 => x"77",
           746 => x"f6",
           747 => x"56",
           748 => x"e7",
           749 => x"f8",
           750 => x"08",
           751 => x"06",
           752 => x"74",
           753 => x"2e",
           754 => x"80",
           755 => x"54",
           756 => x"52",
           757 => x"d0",
           758 => x"56",
           759 => x"38",
           760 => x"88",
           761 => x"83",
           762 => x"55",
           763 => x"c6",
           764 => x"82",
           765 => x"53",
           766 => x"51",
           767 => x"88",
           768 => x"08",
           769 => x"51",
           770 => x"88",
           771 => x"ff",
           772 => x"81",
           773 => x"83",
           774 => x"75",
           775 => x"3d",
           776 => x"3d",
           777 => x"80",
           778 => x"0b",
           779 => x"f5",
           780 => x"08",
           781 => x"82",
           782 => x"f2",
           783 => x"53",
           784 => x"53",
           785 => x"d3",
           786 => x"81",
           787 => x"76",
           788 => x"81",
           789 => x"90",
           790 => x"53",
           791 => x"51",
           792 => x"88",
           793 => x"8d",
           794 => x"74",
           795 => x"38",
           796 => x"05",
           797 => x"3f",
           798 => x"08",
           799 => x"5a",
           800 => x"88",
           801 => x"06",
           802 => x"2e",
           803 => x"86",
           804 => x"82",
           805 => x"80",
           806 => x"86",
           807 => x"39",
           808 => x"53",
           809 => x"51",
           810 => x"81",
           811 => x"81",
           812 => x"3d",
           813 => x"f6",
           814 => x"08",
           815 => x"06",
           816 => x"38",
           817 => x"05",
           818 => x"3f",
           819 => x"02",
           820 => x"78",
           821 => x"88",
           822 => x"70",
           823 => x"5b",
           824 => x"88",
           825 => x"ff",
           826 => x"8c",
           827 => x"3d",
           828 => x"34",
           829 => x"05",
           830 => x"3f",
           831 => x"1a",
           832 => x"e2",
           833 => x"e4",
           834 => x"83",
           835 => x"56",
           836 => x"95",
           837 => x"51",
           838 => x"88",
           839 => x"51",
           840 => x"88",
           841 => x"ff",
           842 => x"31",
           843 => x"1b",
           844 => x"2a",
           845 => x"56",
           846 => x"55",
           847 => x"55",
           848 => x"88",
           849 => x"70",
           850 => x"88",
           851 => x"05",
           852 => x"83",
           853 => x"83",
           854 => x"83",
           855 => x"27",
           856 => x"57",
           857 => x"56",
           858 => x"80",
           859 => x"79",
           860 => x"2e",
           861 => x"90",
           862 => x"fb",
           863 => x"81",
           864 => x"90",
           865 => x"39",
           866 => x"18",
           867 => x"79",
           868 => x"06",
           869 => x"19",
           870 => x"05",
           871 => x"55",
           872 => x"1a",
           873 => x"0b",
           874 => x"0c",
           875 => x"88",
           876 => x"0d",
           877 => x"0d",
           878 => x"9f",
           879 => x"85",
           880 => x"2e",
           881 => x"80",
           882 => x"34",
           883 => x"11",
           884 => x"89",
           885 => x"57",
           886 => x"f8",
           887 => x"08",
           888 => x"80",
           889 => x"3d",
           890 => x"80",
           891 => x"02",
           892 => x"70",
           893 => x"81",
           894 => x"57",
           895 => x"85",
           896 => x"a1",
           897 => x"f5",
           898 => x"08",
           899 => x"98",
           900 => x"51",
           901 => x"88",
           902 => x"0c",
           903 => x"0c",
           904 => x"16",
           905 => x"0c",
           906 => x"04",
           907 => x"7d",
           908 => x"0b",
           909 => x"08",
           910 => x"58",
           911 => x"85",
           912 => x"2e",
           913 => x"81",
           914 => x"06",
           915 => x"74",
           916 => x"c3",
           917 => x"74",
           918 => x"86",
           919 => x"81",
           920 => x"57",
           921 => x"9c",
           922 => x"17",
           923 => x"74",
           924 => x"38",
           925 => x"80",
           926 => x"38",
           927 => x"70",
           928 => x"56",
           929 => x"c7",
           930 => x"33",
           931 => x"89",
           932 => x"81",
           933 => x"55",
           934 => x"76",
           935 => x"16",
           936 => x"39",
           937 => x"51",
           938 => x"88",
           939 => x"75",
           940 => x"38",
           941 => x"0c",
           942 => x"51",
           943 => x"88",
           944 => x"08",
           945 => x"8f",
           946 => x"1a",
           947 => x"98",
           948 => x"ff",
           949 => x"71",
           950 => x"77",
           951 => x"38",
           952 => x"54",
           953 => x"83",
           954 => x"a8",
           955 => x"78",
           956 => x"3f",
           957 => x"e5",
           958 => x"08",
           959 => x"0c",
           960 => x"7b",
           961 => x"0c",
           962 => x"2e",
           963 => x"74",
           964 => x"e2",
           965 => x"76",
           966 => x"3d",
           967 => x"3d",
           968 => x"94",
           969 => x"87",
           970 => x"73",
           971 => x"3f",
           972 => x"2b",
           973 => x"8c",
           974 => x"87",
           975 => x"74",
           976 => x"3f",
           977 => x"07",
           978 => x"8c",
           979 => x"94",
           980 => x"87",
           981 => x"73",
           982 => x"3f",
           983 => x"2b",
           984 => x"9c",
           985 => x"87",
           986 => x"74",
           987 => x"3f",
           988 => x"07",
           989 => x"9c",
           990 => x"83",
           991 => x"94",
           992 => x"80",
           993 => x"c0",
           994 => x"9f",
           995 => x"92",
           996 => x"b8",
           997 => x"51",
           998 => x"88",
           999 => x"a0",
          1000 => x"08",
          1001 => x"88",
          1002 => x"3d",
          1003 => x"84",
          1004 => x"51",
          1005 => x"88",
          1006 => x"75",
          1007 => x"2e",
          1008 => x"15",
          1009 => x"a0",
          1010 => x"04",
          1011 => x"39",
          1012 => x"ff",
          1013 => x"ff",
          1014 => x"00",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"4e",
          1018 => x"4f",
          1019 => x"00",
          1020 => x"00",
          2048 => x"0b",
          2049 => x"0b",
          2050 => x"bb",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"0b",
          2058 => x"84",
          2059 => x"0b",
          2060 => x"0b",
          2061 => x"a3",
          2062 => x"0b",
          2063 => x"0b",
          2064 => x"c3",
          2065 => x"0b",
          2066 => x"0b",
          2067 => x"e3",
          2068 => x"0b",
          2069 => x"0b",
          2070 => x"83",
          2071 => x"0b",
          2072 => x"0b",
          2073 => x"a3",
          2074 => x"0b",
          2075 => x"0b",
          2076 => x"c3",
          2077 => x"0b",
          2078 => x"0b",
          2079 => x"e2",
          2080 => x"0b",
          2081 => x"0b",
          2082 => x"80",
          2083 => x"0b",
          2084 => x"0b",
          2085 => x"9e",
          2086 => x"0b",
          2087 => x"0b",
          2088 => x"be",
          2089 => x"0b",
          2090 => x"0b",
          2091 => x"de",
          2092 => x"0b",
          2093 => x"0b",
          2094 => x"fe",
          2095 => x"0b",
          2096 => x"0b",
          2097 => x"9e",
          2098 => x"0b",
          2099 => x"0b",
          2100 => x"be",
          2101 => x"0b",
          2102 => x"0b",
          2103 => x"de",
          2104 => x"0b",
          2105 => x"0b",
          2106 => x"fe",
          2107 => x"0b",
          2108 => x"0b",
          2109 => x"9e",
          2110 => x"0b",
          2111 => x"0b",
          2112 => x"be",
          2113 => x"0b",
          2114 => x"0b",
          2115 => x"de",
          2116 => x"0b",
          2117 => x"0b",
          2118 => x"fe",
          2119 => x"0b",
          2120 => x"0b",
          2121 => x"9e",
          2122 => x"0b",
          2123 => x"0b",
          2124 => x"be",
          2125 => x"0b",
          2126 => x"0b",
          2127 => x"de",
          2128 => x"0b",
          2129 => x"0b",
          2130 => x"fe",
          2131 => x"0b",
          2132 => x"0b",
          2133 => x"9c",
          2134 => x"0b",
          2135 => x"00",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"80",
          2177 => x"90",
          2178 => x"2d",
          2179 => x"08",
          2180 => x"04",
          2181 => x"0c",
          2182 => x"2d",
          2183 => x"08",
          2184 => x"04",
          2185 => x"0c",
          2186 => x"2d",
          2187 => x"08",
          2188 => x"04",
          2189 => x"0c",
          2190 => x"2d",
          2191 => x"08",
          2192 => x"04",
          2193 => x"0c",
          2194 => x"2d",
          2195 => x"08",
          2196 => x"04",
          2197 => x"0c",
          2198 => x"2d",
          2199 => x"08",
          2200 => x"04",
          2201 => x"0c",
          2202 => x"2d",
          2203 => x"08",
          2204 => x"04",
          2205 => x"0c",
          2206 => x"2d",
          2207 => x"08",
          2208 => x"04",
          2209 => x"0c",
          2210 => x"2d",
          2211 => x"08",
          2212 => x"04",
          2213 => x"0c",
          2214 => x"2d",
          2215 => x"08",
          2216 => x"04",
          2217 => x"0c",
          2218 => x"2d",
          2219 => x"08",
          2220 => x"04",
          2221 => x"0c",
          2222 => x"2d",
          2223 => x"08",
          2224 => x"04",
          2225 => x"0c",
          2226 => x"2d",
          2227 => x"08",
          2228 => x"04",
          2229 => x"0c",
          2230 => x"82",
          2231 => x"83",
          2232 => x"82",
          2233 => x"ba",
          2234 => x"93",
          2235 => x"80",
          2236 => x"93",
          2237 => x"9a",
          2238 => x"90",
          2239 => x"90",
          2240 => x"90",
          2241 => x"2d",
          2242 => x"08",
          2243 => x"04",
          2244 => x"0c",
          2245 => x"82",
          2246 => x"83",
          2247 => x"82",
          2248 => x"81",
          2249 => x"82",
          2250 => x"83",
          2251 => x"82",
          2252 => x"81",
          2253 => x"82",
          2254 => x"83",
          2255 => x"82",
          2256 => x"81",
          2257 => x"82",
          2258 => x"83",
          2259 => x"82",
          2260 => x"81",
          2261 => x"82",
          2262 => x"83",
          2263 => x"82",
          2264 => x"81",
          2265 => x"82",
          2266 => x"83",
          2267 => x"82",
          2268 => x"81",
          2269 => x"82",
          2270 => x"83",
          2271 => x"82",
          2272 => x"81",
          2273 => x"82",
          2274 => x"83",
          2275 => x"82",
          2276 => x"81",
          2277 => x"82",
          2278 => x"83",
          2279 => x"82",
          2280 => x"81",
          2281 => x"82",
          2282 => x"83",
          2283 => x"82",
          2284 => x"81",
          2285 => x"82",
          2286 => x"83",
          2287 => x"82",
          2288 => x"81",
          2289 => x"82",
          2290 => x"83",
          2291 => x"82",
          2292 => x"81",
          2293 => x"82",
          2294 => x"83",
          2295 => x"82",
          2296 => x"81",
          2297 => x"82",
          2298 => x"83",
          2299 => x"82",
          2300 => x"81",
          2301 => x"82",
          2302 => x"83",
          2303 => x"82",
          2304 => x"81",
          2305 => x"82",
          2306 => x"83",
          2307 => x"82",
          2308 => x"81",
          2309 => x"82",
          2310 => x"83",
          2311 => x"82",
          2312 => x"81",
          2313 => x"82",
          2314 => x"83",
          2315 => x"82",
          2316 => x"81",
          2317 => x"82",
          2318 => x"83",
          2319 => x"82",
          2320 => x"81",
          2321 => x"82",
          2322 => x"83",
          2323 => x"82",
          2324 => x"81",
          2325 => x"82",
          2326 => x"83",
          2327 => x"82",
          2328 => x"81",
          2329 => x"82",
          2330 => x"83",
          2331 => x"82",
          2332 => x"81",
          2333 => x"82",
          2334 => x"83",
          2335 => x"82",
          2336 => x"81",
          2337 => x"82",
          2338 => x"83",
          2339 => x"82",
          2340 => x"81",
          2341 => x"82",
          2342 => x"83",
          2343 => x"82",
          2344 => x"81",
          2345 => x"82",
          2346 => x"83",
          2347 => x"82",
          2348 => x"81",
          2349 => x"82",
          2350 => x"83",
          2351 => x"82",
          2352 => x"81",
          2353 => x"82",
          2354 => x"83",
          2355 => x"82",
          2356 => x"80",
          2357 => x"82",
          2358 => x"83",
          2359 => x"82",
          2360 => x"80",
          2361 => x"82",
          2362 => x"83",
          2363 => x"82",
          2364 => x"80",
          2365 => x"82",
          2366 => x"83",
          2367 => x"82",
          2368 => x"b3",
          2369 => x"93",
          2370 => x"80",
          2371 => x"93",
          2372 => x"a5",
          2373 => x"90",
          2374 => x"90",
          2375 => x"90",
          2376 => x"2d",
          2377 => x"08",
          2378 => x"04",
          2379 => x"0c",
          2380 => x"2d",
          2381 => x"08",
          2382 => x"04",
          2383 => x"70",
          2384 => x"27",
          2385 => x"71",
          2386 => x"53",
          2387 => x"0b",
          2388 => x"a4",
          2389 => x"f4",
          2390 => x"04",
          2391 => x"08",
          2392 => x"90",
          2393 => x"0d",
          2394 => x"93",
          2395 => x"05",
          2396 => x"93",
          2397 => x"05",
          2398 => x"c5",
          2399 => x"84",
          2400 => x"93",
          2401 => x"85",
          2402 => x"93",
          2403 => x"82",
          2404 => x"02",
          2405 => x"0c",
          2406 => x"81",
          2407 => x"90",
          2408 => x"08",
          2409 => x"90",
          2410 => x"08",
          2411 => x"82",
          2412 => x"70",
          2413 => x"0c",
          2414 => x"0d",
          2415 => x"0c",
          2416 => x"90",
          2417 => x"93",
          2418 => x"3d",
          2419 => x"82",
          2420 => x"fc",
          2421 => x"0b",
          2422 => x"08",
          2423 => x"82",
          2424 => x"8c",
          2425 => x"93",
          2426 => x"05",
          2427 => x"38",
          2428 => x"08",
          2429 => x"80",
          2430 => x"80",
          2431 => x"90",
          2432 => x"08",
          2433 => x"82",
          2434 => x"8c",
          2435 => x"82",
          2436 => x"8c",
          2437 => x"93",
          2438 => x"05",
          2439 => x"93",
          2440 => x"05",
          2441 => x"39",
          2442 => x"08",
          2443 => x"80",
          2444 => x"38",
          2445 => x"08",
          2446 => x"82",
          2447 => x"88",
          2448 => x"ad",
          2449 => x"90",
          2450 => x"08",
          2451 => x"08",
          2452 => x"31",
          2453 => x"08",
          2454 => x"82",
          2455 => x"f8",
          2456 => x"93",
          2457 => x"05",
          2458 => x"93",
          2459 => x"05",
          2460 => x"90",
          2461 => x"08",
          2462 => x"93",
          2463 => x"05",
          2464 => x"90",
          2465 => x"08",
          2466 => x"93",
          2467 => x"05",
          2468 => x"39",
          2469 => x"08",
          2470 => x"80",
          2471 => x"82",
          2472 => x"88",
          2473 => x"82",
          2474 => x"f4",
          2475 => x"91",
          2476 => x"90",
          2477 => x"08",
          2478 => x"90",
          2479 => x"0c",
          2480 => x"90",
          2481 => x"08",
          2482 => x"0c",
          2483 => x"82",
          2484 => x"04",
          2485 => x"76",
          2486 => x"55",
          2487 => x"8f",
          2488 => x"38",
          2489 => x"83",
          2490 => x"80",
          2491 => x"ff",
          2492 => x"ff",
          2493 => x"72",
          2494 => x"54",
          2495 => x"81",
          2496 => x"ff",
          2497 => x"ff",
          2498 => x"06",
          2499 => x"82",
          2500 => x"86",
          2501 => x"74",
          2502 => x"84",
          2503 => x"71",
          2504 => x"53",
          2505 => x"84",
          2506 => x"71",
          2507 => x"53",
          2508 => x"84",
          2509 => x"71",
          2510 => x"53",
          2511 => x"84",
          2512 => x"71",
          2513 => x"53",
          2514 => x"52",
          2515 => x"c9",
          2516 => x"27",
          2517 => x"70",
          2518 => x"08",
          2519 => x"05",
          2520 => x"12",
          2521 => x"26",
          2522 => x"54",
          2523 => x"fc",
          2524 => x"79",
          2525 => x"05",
          2526 => x"57",
          2527 => x"83",
          2528 => x"38",
          2529 => x"51",
          2530 => x"a4",
          2531 => x"52",
          2532 => x"93",
          2533 => x"70",
          2534 => x"34",
          2535 => x"71",
          2536 => x"81",
          2537 => x"74",
          2538 => x"0c",
          2539 => x"04",
          2540 => x"2b",
          2541 => x"71",
          2542 => x"51",
          2543 => x"72",
          2544 => x"72",
          2545 => x"05",
          2546 => x"71",
          2547 => x"53",
          2548 => x"70",
          2549 => x"0c",
          2550 => x"84",
          2551 => x"f0",
          2552 => x"8f",
          2553 => x"83",
          2554 => x"38",
          2555 => x"84",
          2556 => x"fc",
          2557 => x"83",
          2558 => x"70",
          2559 => x"39",
          2560 => x"76",
          2561 => x"73",
          2562 => x"54",
          2563 => x"70",
          2564 => x"71",
          2565 => x"09",
          2566 => x"fd",
          2567 => x"70",
          2568 => x"81",
          2569 => x"51",
          2570 => x"70",
          2571 => x"14",
          2572 => x"84",
          2573 => x"70",
          2574 => x"70",
          2575 => x"ff",
          2576 => x"f8",
          2577 => x"80",
          2578 => x"53",
          2579 => x"80",
          2580 => x"73",
          2581 => x"81",
          2582 => x"51",
          2583 => x"81",
          2584 => x"70",
          2585 => x"82",
          2586 => x"86",
          2587 => x"fd",
          2588 => x"70",
          2589 => x"53",
          2590 => x"b8",
          2591 => x"08",
          2592 => x"fb",
          2593 => x"06",
          2594 => x"82",
          2595 => x"51",
          2596 => x"70",
          2597 => x"13",
          2598 => x"09",
          2599 => x"ff",
          2600 => x"f8",
          2601 => x"80",
          2602 => x"52",
          2603 => x"2e",
          2604 => x"52",
          2605 => x"70",
          2606 => x"38",
          2607 => x"33",
          2608 => x"f8",
          2609 => x"31",
          2610 => x"0c",
          2611 => x"04",
          2612 => x"78",
          2613 => x"54",
          2614 => x"72",
          2615 => x"d9",
          2616 => x"07",
          2617 => x"70",
          2618 => x"d6",
          2619 => x"53",
          2620 => x"b1",
          2621 => x"74",
          2622 => x"74",
          2623 => x"81",
          2624 => x"72",
          2625 => x"89",
          2626 => x"ff",
          2627 => x"80",
          2628 => x"38",
          2629 => x"15",
          2630 => x"55",
          2631 => x"2e",
          2632 => x"d1",
          2633 => x"74",
          2634 => x"70",
          2635 => x"75",
          2636 => x"71",
          2637 => x"52",
          2638 => x"93",
          2639 => x"3d",
          2640 => x"74",
          2641 => x"73",
          2642 => x"71",
          2643 => x"2e",
          2644 => x"76",
          2645 => x"95",
          2646 => x"53",
          2647 => x"b1",
          2648 => x"70",
          2649 => x"fd",
          2650 => x"70",
          2651 => x"81",
          2652 => x"51",
          2653 => x"38",
          2654 => x"17",
          2655 => x"73",
          2656 => x"74",
          2657 => x"2e",
          2658 => x"76",
          2659 => x"dd",
          2660 => x"82",
          2661 => x"88",
          2662 => x"fe",
          2663 => x"52",
          2664 => x"88",
          2665 => x"86",
          2666 => x"84",
          2667 => x"06",
          2668 => x"14",
          2669 => x"80",
          2670 => x"71",
          2671 => x"0c",
          2672 => x"04",
          2673 => x"77",
          2674 => x"53",
          2675 => x"80",
          2676 => x"38",
          2677 => x"70",
          2678 => x"81",
          2679 => x"81",
          2680 => x"39",
          2681 => x"39",
          2682 => x"80",
          2683 => x"81",
          2684 => x"55",
          2685 => x"2e",
          2686 => x"55",
          2687 => x"84",
          2688 => x"38",
          2689 => x"06",
          2690 => x"2e",
          2691 => x"88",
          2692 => x"70",
          2693 => x"34",
          2694 => x"71",
          2695 => x"93",
          2696 => x"3d",
          2697 => x"3d",
          2698 => x"72",
          2699 => x"91",
          2700 => x"fc",
          2701 => x"51",
          2702 => x"82",
          2703 => x"85",
          2704 => x"83",
          2705 => x"72",
          2706 => x"0c",
          2707 => x"04",
          2708 => x"76",
          2709 => x"ff",
          2710 => x"81",
          2711 => x"26",
          2712 => x"83",
          2713 => x"05",
          2714 => x"70",
          2715 => x"8a",
          2716 => x"33",
          2717 => x"70",
          2718 => x"fe",
          2719 => x"33",
          2720 => x"70",
          2721 => x"f2",
          2722 => x"33",
          2723 => x"70",
          2724 => x"e6",
          2725 => x"22",
          2726 => x"74",
          2727 => x"80",
          2728 => x"13",
          2729 => x"52",
          2730 => x"26",
          2731 => x"81",
          2732 => x"98",
          2733 => x"22",
          2734 => x"bc",
          2735 => x"33",
          2736 => x"b8",
          2737 => x"33",
          2738 => x"b4",
          2739 => x"33",
          2740 => x"b0",
          2741 => x"33",
          2742 => x"ac",
          2743 => x"33",
          2744 => x"a8",
          2745 => x"c0",
          2746 => x"73",
          2747 => x"a0",
          2748 => x"87",
          2749 => x"0c",
          2750 => x"82",
          2751 => x"86",
          2752 => x"f3",
          2753 => x"5b",
          2754 => x"9c",
          2755 => x"0c",
          2756 => x"bc",
          2757 => x"7b",
          2758 => x"98",
          2759 => x"79",
          2760 => x"87",
          2761 => x"08",
          2762 => x"1c",
          2763 => x"98",
          2764 => x"79",
          2765 => x"87",
          2766 => x"08",
          2767 => x"1c",
          2768 => x"98",
          2769 => x"79",
          2770 => x"87",
          2771 => x"08",
          2772 => x"1c",
          2773 => x"98",
          2774 => x"79",
          2775 => x"80",
          2776 => x"83",
          2777 => x"59",
          2778 => x"ff",
          2779 => x"1b",
          2780 => x"1b",
          2781 => x"1b",
          2782 => x"1b",
          2783 => x"1b",
          2784 => x"83",
          2785 => x"52",
          2786 => x"51",
          2787 => x"8f",
          2788 => x"ff",
          2789 => x"8f",
          2790 => x"30",
          2791 => x"51",
          2792 => x"0b",
          2793 => x"fc",
          2794 => x"0d",
          2795 => x"0d",
          2796 => x"82",
          2797 => x"70",
          2798 => x"57",
          2799 => x"c0",
          2800 => x"74",
          2801 => x"38",
          2802 => x"94",
          2803 => x"70",
          2804 => x"81",
          2805 => x"52",
          2806 => x"8c",
          2807 => x"2a",
          2808 => x"51",
          2809 => x"38",
          2810 => x"70",
          2811 => x"51",
          2812 => x"8d",
          2813 => x"2a",
          2814 => x"51",
          2815 => x"be",
          2816 => x"ff",
          2817 => x"c0",
          2818 => x"70",
          2819 => x"38",
          2820 => x"90",
          2821 => x"0c",
          2822 => x"84",
          2823 => x"0d",
          2824 => x"0d",
          2825 => x"33",
          2826 => x"8d",
          2827 => x"81",
          2828 => x"55",
          2829 => x"94",
          2830 => x"80",
          2831 => x"87",
          2832 => x"51",
          2833 => x"96",
          2834 => x"06",
          2835 => x"70",
          2836 => x"38",
          2837 => x"70",
          2838 => x"51",
          2839 => x"72",
          2840 => x"81",
          2841 => x"70",
          2842 => x"38",
          2843 => x"70",
          2844 => x"51",
          2845 => x"38",
          2846 => x"06",
          2847 => x"94",
          2848 => x"80",
          2849 => x"87",
          2850 => x"52",
          2851 => x"87",
          2852 => x"f9",
          2853 => x"54",
          2854 => x"70",
          2855 => x"53",
          2856 => x"77",
          2857 => x"38",
          2858 => x"06",
          2859 => x"0b",
          2860 => x"33",
          2861 => x"06",
          2862 => x"58",
          2863 => x"84",
          2864 => x"2e",
          2865 => x"c0",
          2866 => x"70",
          2867 => x"2a",
          2868 => x"53",
          2869 => x"80",
          2870 => x"71",
          2871 => x"81",
          2872 => x"70",
          2873 => x"81",
          2874 => x"06",
          2875 => x"80",
          2876 => x"71",
          2877 => x"81",
          2878 => x"70",
          2879 => x"74",
          2880 => x"51",
          2881 => x"80",
          2882 => x"2e",
          2883 => x"c0",
          2884 => x"77",
          2885 => x"17",
          2886 => x"81",
          2887 => x"53",
          2888 => x"84",
          2889 => x"93",
          2890 => x"3d",
          2891 => x"3d",
          2892 => x"82",
          2893 => x"70",
          2894 => x"54",
          2895 => x"94",
          2896 => x"80",
          2897 => x"87",
          2898 => x"51",
          2899 => x"82",
          2900 => x"06",
          2901 => x"70",
          2902 => x"38",
          2903 => x"06",
          2904 => x"94",
          2905 => x"80",
          2906 => x"87",
          2907 => x"52",
          2908 => x"81",
          2909 => x"93",
          2910 => x"84",
          2911 => x"fe",
          2912 => x"0b",
          2913 => x"33",
          2914 => x"06",
          2915 => x"c0",
          2916 => x"70",
          2917 => x"38",
          2918 => x"94",
          2919 => x"70",
          2920 => x"81",
          2921 => x"51",
          2922 => x"80",
          2923 => x"72",
          2924 => x"51",
          2925 => x"80",
          2926 => x"2e",
          2927 => x"c0",
          2928 => x"71",
          2929 => x"2b",
          2930 => x"51",
          2931 => x"82",
          2932 => x"84",
          2933 => x"ff",
          2934 => x"c0",
          2935 => x"70",
          2936 => x"06",
          2937 => x"80",
          2938 => x"38",
          2939 => x"a4",
          2940 => x"80",
          2941 => x"9e",
          2942 => x"8e",
          2943 => x"c0",
          2944 => x"82",
          2945 => x"87",
          2946 => x"08",
          2947 => x"0c",
          2948 => x"9c",
          2949 => x"90",
          2950 => x"9e",
          2951 => x"8e",
          2952 => x"c0",
          2953 => x"82",
          2954 => x"87",
          2955 => x"08",
          2956 => x"0c",
          2957 => x"b4",
          2958 => x"a0",
          2959 => x"9e",
          2960 => x"8e",
          2961 => x"c0",
          2962 => x"82",
          2963 => x"87",
          2964 => x"08",
          2965 => x"0c",
          2966 => x"c4",
          2967 => x"b0",
          2968 => x"9e",
          2969 => x"70",
          2970 => x"23",
          2971 => x"84",
          2972 => x"b8",
          2973 => x"9e",
          2974 => x"8e",
          2975 => x"c0",
          2976 => x"82",
          2977 => x"81",
          2978 => x"c4",
          2979 => x"87",
          2980 => x"08",
          2981 => x"0a",
          2982 => x"52",
          2983 => x"83",
          2984 => x"71",
          2985 => x"34",
          2986 => x"c0",
          2987 => x"70",
          2988 => x"06",
          2989 => x"70",
          2990 => x"38",
          2991 => x"82",
          2992 => x"80",
          2993 => x"9e",
          2994 => x"90",
          2995 => x"51",
          2996 => x"80",
          2997 => x"81",
          2998 => x"8e",
          2999 => x"0b",
          3000 => x"90",
          3001 => x"80",
          3002 => x"52",
          3003 => x"2e",
          3004 => x"52",
          3005 => x"c8",
          3006 => x"87",
          3007 => x"08",
          3008 => x"80",
          3009 => x"52",
          3010 => x"83",
          3011 => x"71",
          3012 => x"34",
          3013 => x"c0",
          3014 => x"70",
          3015 => x"06",
          3016 => x"70",
          3017 => x"38",
          3018 => x"82",
          3019 => x"80",
          3020 => x"9e",
          3021 => x"84",
          3022 => x"51",
          3023 => x"80",
          3024 => x"81",
          3025 => x"8e",
          3026 => x"0b",
          3027 => x"90",
          3028 => x"80",
          3029 => x"52",
          3030 => x"2e",
          3031 => x"52",
          3032 => x"cc",
          3033 => x"87",
          3034 => x"08",
          3035 => x"80",
          3036 => x"52",
          3037 => x"83",
          3038 => x"71",
          3039 => x"34",
          3040 => x"c0",
          3041 => x"70",
          3042 => x"06",
          3043 => x"70",
          3044 => x"38",
          3045 => x"82",
          3046 => x"80",
          3047 => x"9e",
          3048 => x"a0",
          3049 => x"52",
          3050 => x"2e",
          3051 => x"52",
          3052 => x"cf",
          3053 => x"9e",
          3054 => x"98",
          3055 => x"8a",
          3056 => x"51",
          3057 => x"d0",
          3058 => x"87",
          3059 => x"08",
          3060 => x"06",
          3061 => x"70",
          3062 => x"38",
          3063 => x"82",
          3064 => x"87",
          3065 => x"08",
          3066 => x"06",
          3067 => x"51",
          3068 => x"82",
          3069 => x"80",
          3070 => x"9e",
          3071 => x"88",
          3072 => x"52",
          3073 => x"83",
          3074 => x"71",
          3075 => x"34",
          3076 => x"90",
          3077 => x"06",
          3078 => x"82",
          3079 => x"83",
          3080 => x"fb",
          3081 => x"f7",
          3082 => x"9d",
          3083 => x"c4",
          3084 => x"80",
          3085 => x"81",
          3086 => x"8a",
          3087 => x"f7",
          3088 => x"85",
          3089 => x"c6",
          3090 => x"80",
          3091 => x"82",
          3092 => x"82",
          3093 => x"11",
          3094 => x"f7",
          3095 => x"cd",
          3096 => x"cb",
          3097 => x"80",
          3098 => x"82",
          3099 => x"82",
          3100 => x"11",
          3101 => x"f7",
          3102 => x"b1",
          3103 => x"c8",
          3104 => x"80",
          3105 => x"82",
          3106 => x"82",
          3107 => x"11",
          3108 => x"f7",
          3109 => x"95",
          3110 => x"c9",
          3111 => x"80",
          3112 => x"82",
          3113 => x"82",
          3114 => x"11",
          3115 => x"f8",
          3116 => x"f9",
          3117 => x"ca",
          3118 => x"80",
          3119 => x"82",
          3120 => x"82",
          3121 => x"11",
          3122 => x"f8",
          3123 => x"dd",
          3124 => x"cf",
          3125 => x"80",
          3126 => x"82",
          3127 => x"52",
          3128 => x"51",
          3129 => x"82",
          3130 => x"54",
          3131 => x"8d",
          3132 => x"d4",
          3133 => x"f8",
          3134 => x"b1",
          3135 => x"d1",
          3136 => x"80",
          3137 => x"82",
          3138 => x"52",
          3139 => x"51",
          3140 => x"82",
          3141 => x"54",
          3142 => x"88",
          3143 => x"ac",
          3144 => x"3f",
          3145 => x"33",
          3146 => x"2e",
          3147 => x"f9",
          3148 => x"95",
          3149 => x"cc",
          3150 => x"80",
          3151 => x"81",
          3152 => x"88",
          3153 => x"8e",
          3154 => x"73",
          3155 => x"38",
          3156 => x"51",
          3157 => x"82",
          3158 => x"54",
          3159 => x"88",
          3160 => x"e4",
          3161 => x"3f",
          3162 => x"51",
          3163 => x"82",
          3164 => x"52",
          3165 => x"51",
          3166 => x"82",
          3167 => x"52",
          3168 => x"51",
          3169 => x"82",
          3170 => x"52",
          3171 => x"51",
          3172 => x"81",
          3173 => x"87",
          3174 => x"8e",
          3175 => x"81",
          3176 => x"8d",
          3177 => x"8e",
          3178 => x"bd",
          3179 => x"75",
          3180 => x"3f",
          3181 => x"08",
          3182 => x"29",
          3183 => x"54",
          3184 => x"84",
          3185 => x"fb",
          3186 => x"e1",
          3187 => x"cb",
          3188 => x"80",
          3189 => x"82",
          3190 => x"56",
          3191 => x"52",
          3192 => x"f8",
          3193 => x"84",
          3194 => x"c0",
          3195 => x"31",
          3196 => x"93",
          3197 => x"81",
          3198 => x"8c",
          3199 => x"8e",
          3200 => x"73",
          3201 => x"38",
          3202 => x"08",
          3203 => x"c0",
          3204 => x"e6",
          3205 => x"93",
          3206 => x"84",
          3207 => x"71",
          3208 => x"82",
          3209 => x"52",
          3210 => x"51",
          3211 => x"82",
          3212 => x"86",
          3213 => x"3d",
          3214 => x"3d",
          3215 => x"05",
          3216 => x"52",
          3217 => x"ac",
          3218 => x"29",
          3219 => x"f5",
          3220 => x"71",
          3221 => x"fc",
          3222 => x"39",
          3223 => x"51",
          3224 => x"fc",
          3225 => x"39",
          3226 => x"51",
          3227 => x"fc",
          3228 => x"39",
          3229 => x"51",
          3230 => x"84",
          3231 => x"71",
          3232 => x"04",
          3233 => x"87",
          3234 => x"70",
          3235 => x"80",
          3236 => x"74",
          3237 => x"8e",
          3238 => x"0c",
          3239 => x"04",
          3240 => x"87",
          3241 => x"70",
          3242 => x"d8",
          3243 => x"72",
          3244 => x"70",
          3245 => x"08",
          3246 => x"8e",
          3247 => x"0c",
          3248 => x"0d",
          3249 => x"87",
          3250 => x"0c",
          3251 => x"d8",
          3252 => x"96",
          3253 => x"fe",
          3254 => x"93",
          3255 => x"38",
          3256 => x"0b",
          3257 => x"0c",
          3258 => x"08",
          3259 => x"52",
          3260 => x"83",
          3261 => x"88",
          3262 => x"93",
          3263 => x"53",
          3264 => x"84",
          3265 => x"0d",
          3266 => x"0d",
          3267 => x"12",
          3268 => x"90",
          3269 => x"15",
          3270 => x"5e",
          3271 => x"59",
          3272 => x"77",
          3273 => x"75",
          3274 => x"08",
          3275 => x"71",
          3276 => x"31",
          3277 => x"80",
          3278 => x"84",
          3279 => x"8c",
          3280 => x"88",
          3281 => x"8c",
          3282 => x"88",
          3283 => x"90",
          3284 => x"94",
          3285 => x"94",
          3286 => x"90",
          3287 => x"39",
          3288 => x"73",
          3289 => x"74",
          3290 => x"77",
          3291 => x"0c",
          3292 => x"04",
          3293 => x"76",
          3294 => x"88",
          3295 => x"53",
          3296 => x"81",
          3297 => x"06",
          3298 => x"12",
          3299 => x"52",
          3300 => x"2e",
          3301 => x"94",
          3302 => x"08",
          3303 => x"0c",
          3304 => x"0c",
          3305 => x"0c",
          3306 => x"39",
          3307 => x"82",
          3308 => x"90",
          3309 => x"8e",
          3310 => x"14",
          3311 => x"8e",
          3312 => x"13",
          3313 => x"12",
          3314 => x"08",
          3315 => x"81",
          3316 => x"84",
          3317 => x"14",
          3318 => x"74",
          3319 => x"06",
          3320 => x"14",
          3321 => x"14",
          3322 => x"08",
          3323 => x"70",
          3324 => x"52",
          3325 => x"8c",
          3326 => x"15",
          3327 => x"13",
          3328 => x"12",
          3329 => x"93",
          3330 => x"3d",
          3331 => x"3d",
          3332 => x"55",
          3333 => x"2e",
          3334 => x"9f",
          3335 => x"82",
          3336 => x"57",
          3337 => x"82",
          3338 => x"84",
          3339 => x"27",
          3340 => x"90",
          3341 => x"ed",
          3342 => x"ff",
          3343 => x"80",
          3344 => x"58",
          3345 => x"82",
          3346 => x"82",
          3347 => x"30",
          3348 => x"84",
          3349 => x"25",
          3350 => x"08",
          3351 => x"70",
          3352 => x"25",
          3353 => x"58",
          3354 => x"56",
          3355 => x"74",
          3356 => x"06",
          3357 => x"88",
          3358 => x"75",
          3359 => x"39",
          3360 => x"93",
          3361 => x"77",
          3362 => x"08",
          3363 => x"82",
          3364 => x"53",
          3365 => x"2e",
          3366 => x"73",
          3367 => x"8c",
          3368 => x"f0",
          3369 => x"08",
          3370 => x"72",
          3371 => x"75",
          3372 => x"88",
          3373 => x"8c",
          3374 => x"75",
          3375 => x"3f",
          3376 => x"93",
          3377 => x"fc",
          3378 => x"93",
          3379 => x"73",
          3380 => x"0c",
          3381 => x"04",
          3382 => x"73",
          3383 => x"2e",
          3384 => x"12",
          3385 => x"3f",
          3386 => x"04",
          3387 => x"02",
          3388 => x"53",
          3389 => x"09",
          3390 => x"38",
          3391 => x"3f",
          3392 => x"08",
          3393 => x"2e",
          3394 => x"72",
          3395 => x"a0",
          3396 => x"82",
          3397 => x"8f",
          3398 => x"98",
          3399 => x"80",
          3400 => x"72",
          3401 => x"84",
          3402 => x"fe",
          3403 => x"97",
          3404 => x"93",
          3405 => x"82",
          3406 => x"54",
          3407 => x"3f",
          3408 => x"98",
          3409 => x"0d",
          3410 => x"0d",
          3411 => x"33",
          3412 => x"06",
          3413 => x"80",
          3414 => x"72",
          3415 => x"51",
          3416 => x"ff",
          3417 => x"39",
          3418 => x"04",
          3419 => x"77",
          3420 => x"08",
          3421 => x"98",
          3422 => x"73",
          3423 => x"ff",
          3424 => x"71",
          3425 => x"38",
          3426 => x"06",
          3427 => x"54",
          3428 => x"e7",
          3429 => x"93",
          3430 => x"3d",
          3431 => x"3d",
          3432 => x"59",
          3433 => x"81",
          3434 => x"56",
          3435 => x"84",
          3436 => x"a5",
          3437 => x"06",
          3438 => x"80",
          3439 => x"81",
          3440 => x"58",
          3441 => x"b0",
          3442 => x"06",
          3443 => x"5a",
          3444 => x"ad",
          3445 => x"06",
          3446 => x"5a",
          3447 => x"05",
          3448 => x"75",
          3449 => x"81",
          3450 => x"77",
          3451 => x"08",
          3452 => x"05",
          3453 => x"5d",
          3454 => x"39",
          3455 => x"72",
          3456 => x"38",
          3457 => x"7b",
          3458 => x"05",
          3459 => x"70",
          3460 => x"33",
          3461 => x"39",
          3462 => x"32",
          3463 => x"72",
          3464 => x"78",
          3465 => x"70",
          3466 => x"07",
          3467 => x"07",
          3468 => x"51",
          3469 => x"80",
          3470 => x"79",
          3471 => x"70",
          3472 => x"33",
          3473 => x"80",
          3474 => x"38",
          3475 => x"e0",
          3476 => x"38",
          3477 => x"81",
          3478 => x"53",
          3479 => x"2e",
          3480 => x"73",
          3481 => x"a2",
          3482 => x"c3",
          3483 => x"38",
          3484 => x"24",
          3485 => x"80",
          3486 => x"8c",
          3487 => x"39",
          3488 => x"2e",
          3489 => x"81",
          3490 => x"80",
          3491 => x"80",
          3492 => x"d5",
          3493 => x"73",
          3494 => x"8e",
          3495 => x"39",
          3496 => x"2e",
          3497 => x"80",
          3498 => x"84",
          3499 => x"56",
          3500 => x"74",
          3501 => x"72",
          3502 => x"38",
          3503 => x"15",
          3504 => x"54",
          3505 => x"38",
          3506 => x"56",
          3507 => x"81",
          3508 => x"72",
          3509 => x"38",
          3510 => x"90",
          3511 => x"06",
          3512 => x"2e",
          3513 => x"51",
          3514 => x"74",
          3515 => x"53",
          3516 => x"fd",
          3517 => x"51",
          3518 => x"ef",
          3519 => x"19",
          3520 => x"53",
          3521 => x"39",
          3522 => x"39",
          3523 => x"39",
          3524 => x"39",
          3525 => x"39",
          3526 => x"d0",
          3527 => x"39",
          3528 => x"70",
          3529 => x"53",
          3530 => x"88",
          3531 => x"19",
          3532 => x"39",
          3533 => x"54",
          3534 => x"74",
          3535 => x"70",
          3536 => x"07",
          3537 => x"55",
          3538 => x"80",
          3539 => x"72",
          3540 => x"38",
          3541 => x"90",
          3542 => x"80",
          3543 => x"5e",
          3544 => x"74",
          3545 => x"3f",
          3546 => x"08",
          3547 => x"7c",
          3548 => x"54",
          3549 => x"82",
          3550 => x"55",
          3551 => x"92",
          3552 => x"53",
          3553 => x"2e",
          3554 => x"14",
          3555 => x"ff",
          3556 => x"14",
          3557 => x"70",
          3558 => x"34",
          3559 => x"30",
          3560 => x"9f",
          3561 => x"57",
          3562 => x"85",
          3563 => x"b1",
          3564 => x"2a",
          3565 => x"51",
          3566 => x"2e",
          3567 => x"3d",
          3568 => x"05",
          3569 => x"34",
          3570 => x"76",
          3571 => x"54",
          3572 => x"72",
          3573 => x"54",
          3574 => x"70",
          3575 => x"56",
          3576 => x"81",
          3577 => x"7b",
          3578 => x"73",
          3579 => x"3f",
          3580 => x"53",
          3581 => x"74",
          3582 => x"53",
          3583 => x"eb",
          3584 => x"77",
          3585 => x"53",
          3586 => x"14",
          3587 => x"54",
          3588 => x"3f",
          3589 => x"74",
          3590 => x"53",
          3591 => x"fb",
          3592 => x"51",
          3593 => x"ef",
          3594 => x"0d",
          3595 => x"0d",
          3596 => x"70",
          3597 => x"08",
          3598 => x"51",
          3599 => x"85",
          3600 => x"fe",
          3601 => x"82",
          3602 => x"85",
          3603 => x"52",
          3604 => x"ca",
          3605 => x"a0",
          3606 => x"73",
          3607 => x"82",
          3608 => x"84",
          3609 => x"fd",
          3610 => x"93",
          3611 => x"82",
          3612 => x"87",
          3613 => x"53",
          3614 => x"fa",
          3615 => x"82",
          3616 => x"85",
          3617 => x"fb",
          3618 => x"79",
          3619 => x"08",
          3620 => x"57",
          3621 => x"71",
          3622 => x"e0",
          3623 => x"9c",
          3624 => x"2d",
          3625 => x"08",
          3626 => x"53",
          3627 => x"80",
          3628 => x"8d",
          3629 => x"72",
          3630 => x"30",
          3631 => x"51",
          3632 => x"80",
          3633 => x"71",
          3634 => x"38",
          3635 => x"97",
          3636 => x"25",
          3637 => x"16",
          3638 => x"25",
          3639 => x"14",
          3640 => x"34",
          3641 => x"72",
          3642 => x"3f",
          3643 => x"73",
          3644 => x"72",
          3645 => x"f7",
          3646 => x"53",
          3647 => x"84",
          3648 => x"0d",
          3649 => x"0d",
          3650 => x"08",
          3651 => x"9c",
          3652 => x"76",
          3653 => x"ef",
          3654 => x"93",
          3655 => x"3d",
          3656 => x"3d",
          3657 => x"5a",
          3658 => x"7a",
          3659 => x"08",
          3660 => x"53",
          3661 => x"09",
          3662 => x"38",
          3663 => x"0c",
          3664 => x"ad",
          3665 => x"06",
          3666 => x"76",
          3667 => x"0c",
          3668 => x"33",
          3669 => x"73",
          3670 => x"81",
          3671 => x"38",
          3672 => x"05",
          3673 => x"08",
          3674 => x"53",
          3675 => x"2e",
          3676 => x"57",
          3677 => x"2e",
          3678 => x"39",
          3679 => x"13",
          3680 => x"08",
          3681 => x"53",
          3682 => x"55",
          3683 => x"80",
          3684 => x"14",
          3685 => x"88",
          3686 => x"27",
          3687 => x"eb",
          3688 => x"53",
          3689 => x"89",
          3690 => x"38",
          3691 => x"55",
          3692 => x"8a",
          3693 => x"a0",
          3694 => x"c2",
          3695 => x"74",
          3696 => x"e0",
          3697 => x"ff",
          3698 => x"d0",
          3699 => x"ff",
          3700 => x"90",
          3701 => x"38",
          3702 => x"81",
          3703 => x"53",
          3704 => x"ca",
          3705 => x"27",
          3706 => x"77",
          3707 => x"08",
          3708 => x"0c",
          3709 => x"33",
          3710 => x"ff",
          3711 => x"80",
          3712 => x"74",
          3713 => x"79",
          3714 => x"74",
          3715 => x"0c",
          3716 => x"04",
          3717 => x"7a",
          3718 => x"80",
          3719 => x"58",
          3720 => x"33",
          3721 => x"a0",
          3722 => x"06",
          3723 => x"13",
          3724 => x"39",
          3725 => x"09",
          3726 => x"38",
          3727 => x"11",
          3728 => x"08",
          3729 => x"54",
          3730 => x"2e",
          3731 => x"80",
          3732 => x"08",
          3733 => x"0c",
          3734 => x"33",
          3735 => x"80",
          3736 => x"38",
          3737 => x"80",
          3738 => x"38",
          3739 => x"57",
          3740 => x"0c",
          3741 => x"33",
          3742 => x"39",
          3743 => x"74",
          3744 => x"38",
          3745 => x"80",
          3746 => x"89",
          3747 => x"38",
          3748 => x"d0",
          3749 => x"55",
          3750 => x"80",
          3751 => x"39",
          3752 => x"d9",
          3753 => x"80",
          3754 => x"27",
          3755 => x"80",
          3756 => x"89",
          3757 => x"70",
          3758 => x"55",
          3759 => x"70",
          3760 => x"55",
          3761 => x"27",
          3762 => x"14",
          3763 => x"06",
          3764 => x"74",
          3765 => x"73",
          3766 => x"38",
          3767 => x"14",
          3768 => x"05",
          3769 => x"08",
          3770 => x"54",
          3771 => x"39",
          3772 => x"84",
          3773 => x"55",
          3774 => x"81",
          3775 => x"93",
          3776 => x"3d",
          3777 => x"3d",
          3778 => x"2b",
          3779 => x"79",
          3780 => x"98",
          3781 => x"13",
          3782 => x"51",
          3783 => x"51",
          3784 => x"81",
          3785 => x"33",
          3786 => x"74",
          3787 => x"81",
          3788 => x"08",
          3789 => x"05",
          3790 => x"71",
          3791 => x"52",
          3792 => x"09",
          3793 => x"38",
          3794 => x"82",
          3795 => x"85",
          3796 => x"fc",
          3797 => x"02",
          3798 => x"05",
          3799 => x"54",
          3800 => x"80",
          3801 => x"88",
          3802 => x"3f",
          3803 => x"fc",
          3804 => x"f2",
          3805 => x"33",
          3806 => x"71",
          3807 => x"81",
          3808 => x"de",
          3809 => x"f3",
          3810 => x"73",
          3811 => x"0d",
          3812 => x"0d",
          3813 => x"05",
          3814 => x"02",
          3815 => x"05",
          3816 => x"d0",
          3817 => x"29",
          3818 => x"05",
          3819 => x"59",
          3820 => x"59",
          3821 => x"86",
          3822 => x"f2",
          3823 => x"8f",
          3824 => x"84",
          3825 => x"f8",
          3826 => x"70",
          3827 => x"5a",
          3828 => x"82",
          3829 => x"75",
          3830 => x"d0",
          3831 => x"29",
          3832 => x"05",
          3833 => x"56",
          3834 => x"2e",
          3835 => x"53",
          3836 => x"51",
          3837 => x"82",
          3838 => x"81",
          3839 => x"82",
          3840 => x"74",
          3841 => x"55",
          3842 => x"87",
          3843 => x"82",
          3844 => x"77",
          3845 => x"38",
          3846 => x"08",
          3847 => x"2e",
          3848 => x"8f",
          3849 => x"74",
          3850 => x"3d",
          3851 => x"76",
          3852 => x"75",
          3853 => x"91",
          3854 => x"cc",
          3855 => x"51",
          3856 => x"3f",
          3857 => x"08",
          3858 => x"ee",
          3859 => x"0d",
          3860 => x"0d",
          3861 => x"52",
          3862 => x"08",
          3863 => x"87",
          3864 => x"84",
          3865 => x"38",
          3866 => x"08",
          3867 => x"52",
          3868 => x"52",
          3869 => x"d5",
          3870 => x"84",
          3871 => x"b8",
          3872 => x"d7",
          3873 => x"93",
          3874 => x"80",
          3875 => x"84",
          3876 => x"38",
          3877 => x"08",
          3878 => x"17",
          3879 => x"74",
          3880 => x"76",
          3881 => x"81",
          3882 => x"57",
          3883 => x"74",
          3884 => x"81",
          3885 => x"38",
          3886 => x"04",
          3887 => x"aa",
          3888 => x"3d",
          3889 => x"81",
          3890 => x"80",
          3891 => x"cc",
          3892 => x"d1",
          3893 => x"93",
          3894 => x"91",
          3895 => x"82",
          3896 => x"54",
          3897 => x"52",
          3898 => x"52",
          3899 => x"dd",
          3900 => x"84",
          3901 => x"a4",
          3902 => x"d6",
          3903 => x"93",
          3904 => x"18",
          3905 => x"0b",
          3906 => x"08",
          3907 => x"82",
          3908 => x"ff",
          3909 => x"55",
          3910 => x"34",
          3911 => x"30",
          3912 => x"9f",
          3913 => x"55",
          3914 => x"85",
          3915 => x"ad",
          3916 => x"cc",
          3917 => x"08",
          3918 => x"d0",
          3919 => x"93",
          3920 => x"2e",
          3921 => x"fd",
          3922 => x"fd",
          3923 => x"2e",
          3924 => x"99",
          3925 => x"79",
          3926 => x"3f",
          3927 => x"8f",
          3928 => x"08",
          3929 => x"84",
          3930 => x"80",
          3931 => x"93",
          3932 => x"3d",
          3933 => x"3d",
          3934 => x"71",
          3935 => x"33",
          3936 => x"58",
          3937 => x"09",
          3938 => x"38",
          3939 => x"05",
          3940 => x"27",
          3941 => x"17",
          3942 => x"71",
          3943 => x"55",
          3944 => x"09",
          3945 => x"38",
          3946 => x"ea",
          3947 => x"73",
          3948 => x"8f",
          3949 => x"08",
          3950 => x"b3",
          3951 => x"84",
          3952 => x"52",
          3953 => x"d6",
          3954 => x"93",
          3955 => x"c4",
          3956 => x"33",
          3957 => x"2e",
          3958 => x"82",
          3959 => x"b4",
          3960 => x"3f",
          3961 => x"1a",
          3962 => x"fc",
          3963 => x"05",
          3964 => x"3f",
          3965 => x"08",
          3966 => x"38",
          3967 => x"52",
          3968 => x"b8",
          3969 => x"84",
          3970 => x"06",
          3971 => x"38",
          3972 => x"39",
          3973 => x"81",
          3974 => x"54",
          3975 => x"ff",
          3976 => x"54",
          3977 => x"84",
          3978 => x"0d",
          3979 => x"0d",
          3980 => x"02",
          3981 => x"c3",
          3982 => x"5a",
          3983 => x"3d",
          3984 => x"d0",
          3985 => x"8f",
          3986 => x"a3",
          3987 => x"c8",
          3988 => x"81",
          3989 => x"51",
          3990 => x"82",
          3991 => x"82",
          3992 => x"82",
          3993 => x"80",
          3994 => x"38",
          3995 => x"8e",
          3996 => x"82",
          3997 => x"51",
          3998 => x"82",
          3999 => x"80",
          4000 => x"81",
          4001 => x"f3",
          4002 => x"e3",
          4003 => x"cc",
          4004 => x"f8",
          4005 => x"70",
          4006 => x"f6",
          4007 => x"93",
          4008 => x"82",
          4009 => x"74",
          4010 => x"06",
          4011 => x"82",
          4012 => x"51",
          4013 => x"82",
          4014 => x"55",
          4015 => x"93",
          4016 => x"9a",
          4017 => x"84",
          4018 => x"70",
          4019 => x"80",
          4020 => x"53",
          4021 => x"06",
          4022 => x"f9",
          4023 => x"ff",
          4024 => x"06",
          4025 => x"87",
          4026 => x"82",
          4027 => x"8f",
          4028 => x"8b",
          4029 => x"84",
          4030 => x"70",
          4031 => x"59",
          4032 => x"ee",
          4033 => x"ff",
          4034 => x"a8",
          4035 => x"2b",
          4036 => x"82",
          4037 => x"70",
          4038 => x"97",
          4039 => x"2c",
          4040 => x"29",
          4041 => x"05",
          4042 => x"70",
          4043 => x"51",
          4044 => x"51",
          4045 => x"81",
          4046 => x"2e",
          4047 => x"77",
          4048 => x"38",
          4049 => x"0a",
          4050 => x"0a",
          4051 => x"2c",
          4052 => x"75",
          4053 => x"38",
          4054 => x"52",
          4055 => x"a6",
          4056 => x"84",
          4057 => x"06",
          4058 => x"2e",
          4059 => x"82",
          4060 => x"81",
          4061 => x"74",
          4062 => x"29",
          4063 => x"05",
          4064 => x"70",
          4065 => x"56",
          4066 => x"8a",
          4067 => x"76",
          4068 => x"77",
          4069 => x"3f",
          4070 => x"08",
          4071 => x"54",
          4072 => x"d3",
          4073 => x"75",
          4074 => x"ca",
          4075 => x"55",
          4076 => x"a8",
          4077 => x"2b",
          4078 => x"82",
          4079 => x"70",
          4080 => x"98",
          4081 => x"11",
          4082 => x"81",
          4083 => x"33",
          4084 => x"51",
          4085 => x"55",
          4086 => x"09",
          4087 => x"92",
          4088 => x"e4",
          4089 => x"0c",
          4090 => x"93",
          4091 => x"0b",
          4092 => x"34",
          4093 => x"82",
          4094 => x"75",
          4095 => x"34",
          4096 => x"34",
          4097 => x"7e",
          4098 => x"26",
          4099 => x"73",
          4100 => x"f5",
          4101 => x"73",
          4102 => x"93",
          4103 => x"73",
          4104 => x"cb",
          4105 => x"ac",
          4106 => x"75",
          4107 => x"74",
          4108 => x"98",
          4109 => x"73",
          4110 => x"38",
          4111 => x"73",
          4112 => x"34",
          4113 => x"0a",
          4114 => x"0a",
          4115 => x"2c",
          4116 => x"33",
          4117 => x"df",
          4118 => x"b0",
          4119 => x"56",
          4120 => x"93",
          4121 => x"1a",
          4122 => x"33",
          4123 => x"93",
          4124 => x"73",
          4125 => x"38",
          4126 => x"73",
          4127 => x"34",
          4128 => x"33",
          4129 => x"0a",
          4130 => x"0a",
          4131 => x"2c",
          4132 => x"33",
          4133 => x"56",
          4134 => x"a2",
          4135 => x"70",
          4136 => x"e8",
          4137 => x"81",
          4138 => x"81",
          4139 => x"70",
          4140 => x"93",
          4141 => x"51",
          4142 => x"24",
          4143 => x"93",
          4144 => x"98",
          4145 => x"2c",
          4146 => x"33",
          4147 => x"56",
          4148 => x"fc",
          4149 => x"51",
          4150 => x"74",
          4151 => x"29",
          4152 => x"05",
          4153 => x"82",
          4154 => x"56",
          4155 => x"75",
          4156 => x"fb",
          4157 => x"93",
          4158 => x"81",
          4159 => x"55",
          4160 => x"fb",
          4161 => x"93",
          4162 => x"05",
          4163 => x"93",
          4164 => x"15",
          4165 => x"93",
          4166 => x"51",
          4167 => x"82",
          4168 => x"70",
          4169 => x"98",
          4170 => x"ac",
          4171 => x"56",
          4172 => x"25",
          4173 => x"1a",
          4174 => x"33",
          4175 => x"33",
          4176 => x"3f",
          4177 => x"0a",
          4178 => x"0a",
          4179 => x"2c",
          4180 => x"33",
          4181 => x"75",
          4182 => x"38",
          4183 => x"8c",
          4184 => x"b0",
          4185 => x"2b",
          4186 => x"82",
          4187 => x"57",
          4188 => x"74",
          4189 => x"f7",
          4190 => x"e6",
          4191 => x"81",
          4192 => x"81",
          4193 => x"70",
          4194 => x"93",
          4195 => x"51",
          4196 => x"25",
          4197 => x"d7",
          4198 => x"ac",
          4199 => x"54",
          4200 => x"8a",
          4201 => x"3f",
          4202 => x"52",
          4203 => x"c6",
          4204 => x"84",
          4205 => x"06",
          4206 => x"38",
          4207 => x"33",
          4208 => x"2e",
          4209 => x"81",
          4210 => x"79",
          4211 => x"3f",
          4212 => x"80",
          4213 => x"b7",
          4214 => x"b0",
          4215 => x"80",
          4216 => x"38",
          4217 => x"84",
          4218 => x"b0",
          4219 => x"54",
          4220 => x"b0",
          4221 => x"ff",
          4222 => x"39",
          4223 => x"33",
          4224 => x"33",
          4225 => x"75",
          4226 => x"38",
          4227 => x"73",
          4228 => x"34",
          4229 => x"70",
          4230 => x"81",
          4231 => x"51",
          4232 => x"25",
          4233 => x"1a",
          4234 => x"33",
          4235 => x"33",
          4236 => x"3f",
          4237 => x"0a",
          4238 => x"0a",
          4239 => x"2c",
          4240 => x"33",
          4241 => x"75",
          4242 => x"38",
          4243 => x"9c",
          4244 => x"b0",
          4245 => x"2b",
          4246 => x"82",
          4247 => x"57",
          4248 => x"74",
          4249 => x"87",
          4250 => x"e4",
          4251 => x"81",
          4252 => x"81",
          4253 => x"70",
          4254 => x"93",
          4255 => x"51",
          4256 => x"25",
          4257 => x"e7",
          4258 => x"b0",
          4259 => x"ff",
          4260 => x"ac",
          4261 => x"54",
          4262 => x"f8",
          4263 => x"14",
          4264 => x"93",
          4265 => x"1a",
          4266 => x"54",
          4267 => x"82",
          4268 => x"70",
          4269 => x"82",
          4270 => x"58",
          4271 => x"75",
          4272 => x"f8",
          4273 => x"ae",
          4274 => x"c4",
          4275 => x"80",
          4276 => x"74",
          4277 => x"3f",
          4278 => x"08",
          4279 => x"34",
          4280 => x"08",
          4281 => x"81",
          4282 => x"52",
          4283 => x"e4",
          4284 => x"81",
          4285 => x"84",
          4286 => x"f8",
          4287 => x"08",
          4288 => x"80",
          4289 => x"74",
          4290 => x"3f",
          4291 => x"08",
          4292 => x"34",
          4293 => x"08",
          4294 => x"81",
          4295 => x"52",
          4296 => x"b0",
          4297 => x"54",
          4298 => x"73",
          4299 => x"80",
          4300 => x"38",
          4301 => x"b7",
          4302 => x"39",
          4303 => x"09",
          4304 => x"38",
          4305 => x"08",
          4306 => x"2e",
          4307 => x"51",
          4308 => x"80",
          4309 => x"84",
          4310 => x"f8",
          4311 => x"08",
          4312 => x"80",
          4313 => x"74",
          4314 => x"3f",
          4315 => x"08",
          4316 => x"34",
          4317 => x"08",
          4318 => x"81",
          4319 => x"52",
          4320 => x"d0",
          4321 => x"54",
          4322 => x"06",
          4323 => x"73",
          4324 => x"80",
          4325 => x"38",
          4326 => x"d3",
          4327 => x"84",
          4328 => x"ac",
          4329 => x"84",
          4330 => x"06",
          4331 => x"74",
          4332 => x"c6",
          4333 => x"93",
          4334 => x"93",
          4335 => x"79",
          4336 => x"3f",
          4337 => x"82",
          4338 => x"70",
          4339 => x"82",
          4340 => x"59",
          4341 => x"77",
          4342 => x"38",
          4343 => x"73",
          4344 => x"34",
          4345 => x"33",
          4346 => x"80",
          4347 => x"39",
          4348 => x"33",
          4349 => x"2e",
          4350 => x"88",
          4351 => x"3f",
          4352 => x"33",
          4353 => x"73",
          4354 => x"34",
          4355 => x"80",
          4356 => x"b0",
          4357 => x"82",
          4358 => x"79",
          4359 => x"0c",
          4360 => x"04",
          4361 => x"02",
          4362 => x"51",
          4363 => x"72",
          4364 => x"82",
          4365 => x"33",
          4366 => x"93",
          4367 => x"3d",
          4368 => x"3d",
          4369 => x"05",
          4370 => x"05",
          4371 => x"56",
          4372 => x"72",
          4373 => x"e0",
          4374 => x"2b",
          4375 => x"8c",
          4376 => x"88",
          4377 => x"2e",
          4378 => x"88",
          4379 => x"0c",
          4380 => x"8c",
          4381 => x"71",
          4382 => x"87",
          4383 => x"0c",
          4384 => x"08",
          4385 => x"51",
          4386 => x"2e",
          4387 => x"c0",
          4388 => x"51",
          4389 => x"71",
          4390 => x"80",
          4391 => x"92",
          4392 => x"98",
          4393 => x"70",
          4394 => x"38",
          4395 => x"ec",
          4396 => x"8f",
          4397 => x"51",
          4398 => x"84",
          4399 => x"0d",
          4400 => x"0d",
          4401 => x"02",
          4402 => x"05",
          4403 => x"58",
          4404 => x"52",
          4405 => x"3f",
          4406 => x"08",
          4407 => x"54",
          4408 => x"be",
          4409 => x"75",
          4410 => x"c0",
          4411 => x"87",
          4412 => x"12",
          4413 => x"84",
          4414 => x"40",
          4415 => x"85",
          4416 => x"98",
          4417 => x"7d",
          4418 => x"0c",
          4419 => x"85",
          4420 => x"06",
          4421 => x"71",
          4422 => x"38",
          4423 => x"71",
          4424 => x"05",
          4425 => x"19",
          4426 => x"a2",
          4427 => x"71",
          4428 => x"38",
          4429 => x"83",
          4430 => x"38",
          4431 => x"8a",
          4432 => x"98",
          4433 => x"71",
          4434 => x"c0",
          4435 => x"52",
          4436 => x"87",
          4437 => x"80",
          4438 => x"81",
          4439 => x"c0",
          4440 => x"53",
          4441 => x"82",
          4442 => x"71",
          4443 => x"1a",
          4444 => x"84",
          4445 => x"19",
          4446 => x"06",
          4447 => x"79",
          4448 => x"38",
          4449 => x"80",
          4450 => x"87",
          4451 => x"26",
          4452 => x"73",
          4453 => x"06",
          4454 => x"2e",
          4455 => x"52",
          4456 => x"82",
          4457 => x"8f",
          4458 => x"f3",
          4459 => x"62",
          4460 => x"05",
          4461 => x"57",
          4462 => x"83",
          4463 => x"52",
          4464 => x"3f",
          4465 => x"08",
          4466 => x"54",
          4467 => x"2e",
          4468 => x"81",
          4469 => x"74",
          4470 => x"c0",
          4471 => x"87",
          4472 => x"12",
          4473 => x"84",
          4474 => x"5f",
          4475 => x"0b",
          4476 => x"8c",
          4477 => x"0c",
          4478 => x"80",
          4479 => x"70",
          4480 => x"81",
          4481 => x"54",
          4482 => x"8c",
          4483 => x"81",
          4484 => x"7c",
          4485 => x"58",
          4486 => x"70",
          4487 => x"52",
          4488 => x"8a",
          4489 => x"98",
          4490 => x"71",
          4491 => x"c0",
          4492 => x"52",
          4493 => x"87",
          4494 => x"80",
          4495 => x"81",
          4496 => x"c0",
          4497 => x"53",
          4498 => x"82",
          4499 => x"71",
          4500 => x"19",
          4501 => x"81",
          4502 => x"ff",
          4503 => x"19",
          4504 => x"78",
          4505 => x"38",
          4506 => x"80",
          4507 => x"87",
          4508 => x"26",
          4509 => x"73",
          4510 => x"06",
          4511 => x"2e",
          4512 => x"52",
          4513 => x"82",
          4514 => x"8f",
          4515 => x"fa",
          4516 => x"02",
          4517 => x"05",
          4518 => x"05",
          4519 => x"71",
          4520 => x"57",
          4521 => x"82",
          4522 => x"81",
          4523 => x"54",
          4524 => x"38",
          4525 => x"c0",
          4526 => x"81",
          4527 => x"2e",
          4528 => x"71",
          4529 => x"38",
          4530 => x"87",
          4531 => x"11",
          4532 => x"80",
          4533 => x"80",
          4534 => x"83",
          4535 => x"38",
          4536 => x"72",
          4537 => x"2a",
          4538 => x"51",
          4539 => x"80",
          4540 => x"87",
          4541 => x"08",
          4542 => x"38",
          4543 => x"8c",
          4544 => x"96",
          4545 => x"0c",
          4546 => x"8c",
          4547 => x"08",
          4548 => x"51",
          4549 => x"38",
          4550 => x"56",
          4551 => x"80",
          4552 => x"85",
          4553 => x"77",
          4554 => x"83",
          4555 => x"75",
          4556 => x"93",
          4557 => x"3d",
          4558 => x"3d",
          4559 => x"11",
          4560 => x"71",
          4561 => x"82",
          4562 => x"53",
          4563 => x"0d",
          4564 => x"0d",
          4565 => x"33",
          4566 => x"71",
          4567 => x"88",
          4568 => x"14",
          4569 => x"07",
          4570 => x"33",
          4571 => x"93",
          4572 => x"53",
          4573 => x"52",
          4574 => x"04",
          4575 => x"73",
          4576 => x"92",
          4577 => x"52",
          4578 => x"81",
          4579 => x"70",
          4580 => x"70",
          4581 => x"3d",
          4582 => x"3d",
          4583 => x"52",
          4584 => x"70",
          4585 => x"34",
          4586 => x"51",
          4587 => x"81",
          4588 => x"70",
          4589 => x"70",
          4590 => x"05",
          4591 => x"88",
          4592 => x"72",
          4593 => x"0d",
          4594 => x"0d",
          4595 => x"54",
          4596 => x"80",
          4597 => x"71",
          4598 => x"53",
          4599 => x"81",
          4600 => x"ff",
          4601 => x"39",
          4602 => x"04",
          4603 => x"75",
          4604 => x"52",
          4605 => x"70",
          4606 => x"34",
          4607 => x"70",
          4608 => x"3d",
          4609 => x"3d",
          4610 => x"79",
          4611 => x"74",
          4612 => x"56",
          4613 => x"81",
          4614 => x"71",
          4615 => x"16",
          4616 => x"52",
          4617 => x"86",
          4618 => x"2e",
          4619 => x"82",
          4620 => x"86",
          4621 => x"fe",
          4622 => x"76",
          4623 => x"39",
          4624 => x"8a",
          4625 => x"51",
          4626 => x"71",
          4627 => x"33",
          4628 => x"0c",
          4629 => x"04",
          4630 => x"93",
          4631 => x"80",
          4632 => x"84",
          4633 => x"3d",
          4634 => x"80",
          4635 => x"33",
          4636 => x"7a",
          4637 => x"38",
          4638 => x"16",
          4639 => x"16",
          4640 => x"17",
          4641 => x"fa",
          4642 => x"93",
          4643 => x"2e",
          4644 => x"b7",
          4645 => x"84",
          4646 => x"34",
          4647 => x"70",
          4648 => x"31",
          4649 => x"59",
          4650 => x"77",
          4651 => x"82",
          4652 => x"74",
          4653 => x"81",
          4654 => x"81",
          4655 => x"53",
          4656 => x"16",
          4657 => x"e3",
          4658 => x"81",
          4659 => x"93",
          4660 => x"3d",
          4661 => x"3d",
          4662 => x"56",
          4663 => x"74",
          4664 => x"2e",
          4665 => x"51",
          4666 => x"82",
          4667 => x"57",
          4668 => x"08",
          4669 => x"54",
          4670 => x"16",
          4671 => x"33",
          4672 => x"3f",
          4673 => x"08",
          4674 => x"38",
          4675 => x"57",
          4676 => x"0c",
          4677 => x"84",
          4678 => x"0d",
          4679 => x"0d",
          4680 => x"57",
          4681 => x"82",
          4682 => x"58",
          4683 => x"08",
          4684 => x"76",
          4685 => x"83",
          4686 => x"06",
          4687 => x"84",
          4688 => x"78",
          4689 => x"81",
          4690 => x"38",
          4691 => x"82",
          4692 => x"52",
          4693 => x"52",
          4694 => x"3f",
          4695 => x"52",
          4696 => x"51",
          4697 => x"84",
          4698 => x"d2",
          4699 => x"fc",
          4700 => x"8a",
          4701 => x"52",
          4702 => x"51",
          4703 => x"90",
          4704 => x"84",
          4705 => x"fc",
          4706 => x"17",
          4707 => x"a0",
          4708 => x"86",
          4709 => x"08",
          4710 => x"b0",
          4711 => x"55",
          4712 => x"81",
          4713 => x"f8",
          4714 => x"84",
          4715 => x"53",
          4716 => x"17",
          4717 => x"d7",
          4718 => x"84",
          4719 => x"83",
          4720 => x"77",
          4721 => x"0c",
          4722 => x"04",
          4723 => x"77",
          4724 => x"12",
          4725 => x"55",
          4726 => x"56",
          4727 => x"8d",
          4728 => x"22",
          4729 => x"ac",
          4730 => x"57",
          4731 => x"93",
          4732 => x"3d",
          4733 => x"3d",
          4734 => x"70",
          4735 => x"57",
          4736 => x"81",
          4737 => x"98",
          4738 => x"81",
          4739 => x"74",
          4740 => x"72",
          4741 => x"f5",
          4742 => x"24",
          4743 => x"81",
          4744 => x"81",
          4745 => x"83",
          4746 => x"38",
          4747 => x"76",
          4748 => x"70",
          4749 => x"16",
          4750 => x"74",
          4751 => x"96",
          4752 => x"84",
          4753 => x"38",
          4754 => x"06",
          4755 => x"33",
          4756 => x"89",
          4757 => x"08",
          4758 => x"54",
          4759 => x"fc",
          4760 => x"93",
          4761 => x"fe",
          4762 => x"ff",
          4763 => x"11",
          4764 => x"2b",
          4765 => x"81",
          4766 => x"2a",
          4767 => x"51",
          4768 => x"e2",
          4769 => x"ff",
          4770 => x"da",
          4771 => x"2a",
          4772 => x"05",
          4773 => x"fc",
          4774 => x"93",
          4775 => x"c6",
          4776 => x"83",
          4777 => x"05",
          4778 => x"f9",
          4779 => x"93",
          4780 => x"ff",
          4781 => x"ae",
          4782 => x"2a",
          4783 => x"05",
          4784 => x"fc",
          4785 => x"93",
          4786 => x"38",
          4787 => x"83",
          4788 => x"05",
          4789 => x"f8",
          4790 => x"93",
          4791 => x"0a",
          4792 => x"39",
          4793 => x"82",
          4794 => x"89",
          4795 => x"f8",
          4796 => x"7c",
          4797 => x"56",
          4798 => x"77",
          4799 => x"38",
          4800 => x"08",
          4801 => x"38",
          4802 => x"72",
          4803 => x"9d",
          4804 => x"24",
          4805 => x"81",
          4806 => x"82",
          4807 => x"83",
          4808 => x"38",
          4809 => x"76",
          4810 => x"70",
          4811 => x"18",
          4812 => x"76",
          4813 => x"9e",
          4814 => x"84",
          4815 => x"93",
          4816 => x"d9",
          4817 => x"ff",
          4818 => x"05",
          4819 => x"81",
          4820 => x"54",
          4821 => x"80",
          4822 => x"77",
          4823 => x"f0",
          4824 => x"8f",
          4825 => x"51",
          4826 => x"34",
          4827 => x"17",
          4828 => x"2a",
          4829 => x"05",
          4830 => x"fa",
          4831 => x"93",
          4832 => x"82",
          4833 => x"81",
          4834 => x"83",
          4835 => x"b4",
          4836 => x"2a",
          4837 => x"8f",
          4838 => x"2a",
          4839 => x"f0",
          4840 => x"06",
          4841 => x"72",
          4842 => x"ec",
          4843 => x"2a",
          4844 => x"05",
          4845 => x"fa",
          4846 => x"93",
          4847 => x"82",
          4848 => x"80",
          4849 => x"83",
          4850 => x"52",
          4851 => x"fe",
          4852 => x"b4",
          4853 => x"a4",
          4854 => x"76",
          4855 => x"17",
          4856 => x"75",
          4857 => x"3f",
          4858 => x"08",
          4859 => x"84",
          4860 => x"77",
          4861 => x"77",
          4862 => x"fc",
          4863 => x"b4",
          4864 => x"51",
          4865 => x"c9",
          4866 => x"84",
          4867 => x"06",
          4868 => x"72",
          4869 => x"3f",
          4870 => x"17",
          4871 => x"93",
          4872 => x"3d",
          4873 => x"3d",
          4874 => x"7e",
          4875 => x"56",
          4876 => x"75",
          4877 => x"74",
          4878 => x"27",
          4879 => x"80",
          4880 => x"ff",
          4881 => x"75",
          4882 => x"3f",
          4883 => x"08",
          4884 => x"84",
          4885 => x"38",
          4886 => x"54",
          4887 => x"81",
          4888 => x"39",
          4889 => x"08",
          4890 => x"39",
          4891 => x"51",
          4892 => x"82",
          4893 => x"58",
          4894 => x"08",
          4895 => x"c7",
          4896 => x"84",
          4897 => x"d2",
          4898 => x"84",
          4899 => x"cf",
          4900 => x"74",
          4901 => x"fc",
          4902 => x"93",
          4903 => x"38",
          4904 => x"fe",
          4905 => x"08",
          4906 => x"74",
          4907 => x"38",
          4908 => x"17",
          4909 => x"33",
          4910 => x"73",
          4911 => x"77",
          4912 => x"26",
          4913 => x"80",
          4914 => x"93",
          4915 => x"3d",
          4916 => x"3d",
          4917 => x"71",
          4918 => x"5b",
          4919 => x"8c",
          4920 => x"77",
          4921 => x"38",
          4922 => x"78",
          4923 => x"81",
          4924 => x"79",
          4925 => x"f9",
          4926 => x"55",
          4927 => x"84",
          4928 => x"e0",
          4929 => x"84",
          4930 => x"93",
          4931 => x"2e",
          4932 => x"98",
          4933 => x"93",
          4934 => x"82",
          4935 => x"58",
          4936 => x"70",
          4937 => x"80",
          4938 => x"38",
          4939 => x"09",
          4940 => x"e2",
          4941 => x"56",
          4942 => x"76",
          4943 => x"82",
          4944 => x"7a",
          4945 => x"3f",
          4946 => x"93",
          4947 => x"2e",
          4948 => x"86",
          4949 => x"84",
          4950 => x"93",
          4951 => x"70",
          4952 => x"07",
          4953 => x"7c",
          4954 => x"84",
          4955 => x"51",
          4956 => x"81",
          4957 => x"93",
          4958 => x"2e",
          4959 => x"17",
          4960 => x"74",
          4961 => x"73",
          4962 => x"27",
          4963 => x"58",
          4964 => x"80",
          4965 => x"56",
          4966 => x"98",
          4967 => x"26",
          4968 => x"56",
          4969 => x"81",
          4970 => x"52",
          4971 => x"c6",
          4972 => x"84",
          4973 => x"b8",
          4974 => x"82",
          4975 => x"81",
          4976 => x"06",
          4977 => x"93",
          4978 => x"82",
          4979 => x"09",
          4980 => x"72",
          4981 => x"70",
          4982 => x"51",
          4983 => x"80",
          4984 => x"78",
          4985 => x"06",
          4986 => x"73",
          4987 => x"39",
          4988 => x"52",
          4989 => x"f7",
          4990 => x"84",
          4991 => x"84",
          4992 => x"82",
          4993 => x"07",
          4994 => x"55",
          4995 => x"2e",
          4996 => x"80",
          4997 => x"75",
          4998 => x"76",
          4999 => x"3f",
          5000 => x"08",
          5001 => x"38",
          5002 => x"0c",
          5003 => x"fe",
          5004 => x"08",
          5005 => x"74",
          5006 => x"ff",
          5007 => x"0c",
          5008 => x"81",
          5009 => x"84",
          5010 => x"39",
          5011 => x"81",
          5012 => x"8c",
          5013 => x"8c",
          5014 => x"84",
          5015 => x"39",
          5016 => x"55",
          5017 => x"84",
          5018 => x"0d",
          5019 => x"0d",
          5020 => x"55",
          5021 => x"82",
          5022 => x"58",
          5023 => x"93",
          5024 => x"d8",
          5025 => x"74",
          5026 => x"3f",
          5027 => x"08",
          5028 => x"08",
          5029 => x"59",
          5030 => x"77",
          5031 => x"70",
          5032 => x"c8",
          5033 => x"84",
          5034 => x"56",
          5035 => x"58",
          5036 => x"97",
          5037 => x"75",
          5038 => x"52",
          5039 => x"51",
          5040 => x"82",
          5041 => x"80",
          5042 => x"8a",
          5043 => x"32",
          5044 => x"72",
          5045 => x"2a",
          5046 => x"56",
          5047 => x"84",
          5048 => x"0d",
          5049 => x"0d",
          5050 => x"08",
          5051 => x"74",
          5052 => x"26",
          5053 => x"74",
          5054 => x"72",
          5055 => x"74",
          5056 => x"88",
          5057 => x"73",
          5058 => x"33",
          5059 => x"27",
          5060 => x"16",
          5061 => x"9b",
          5062 => x"2a",
          5063 => x"88",
          5064 => x"58",
          5065 => x"80",
          5066 => x"16",
          5067 => x"0c",
          5068 => x"8a",
          5069 => x"89",
          5070 => x"72",
          5071 => x"38",
          5072 => x"51",
          5073 => x"82",
          5074 => x"54",
          5075 => x"08",
          5076 => x"38",
          5077 => x"93",
          5078 => x"8b",
          5079 => x"08",
          5080 => x"08",
          5081 => x"82",
          5082 => x"74",
          5083 => x"cb",
          5084 => x"75",
          5085 => x"3f",
          5086 => x"08",
          5087 => x"73",
          5088 => x"98",
          5089 => x"82",
          5090 => x"2e",
          5091 => x"39",
          5092 => x"39",
          5093 => x"13",
          5094 => x"74",
          5095 => x"16",
          5096 => x"18",
          5097 => x"77",
          5098 => x"0c",
          5099 => x"04",
          5100 => x"7a",
          5101 => x"12",
          5102 => x"59",
          5103 => x"80",
          5104 => x"86",
          5105 => x"98",
          5106 => x"14",
          5107 => x"55",
          5108 => x"81",
          5109 => x"83",
          5110 => x"77",
          5111 => x"81",
          5112 => x"0c",
          5113 => x"55",
          5114 => x"76",
          5115 => x"17",
          5116 => x"74",
          5117 => x"9b",
          5118 => x"39",
          5119 => x"ff",
          5120 => x"2a",
          5121 => x"81",
          5122 => x"52",
          5123 => x"e6",
          5124 => x"84",
          5125 => x"55",
          5126 => x"93",
          5127 => x"80",
          5128 => x"55",
          5129 => x"08",
          5130 => x"f4",
          5131 => x"08",
          5132 => x"08",
          5133 => x"38",
          5134 => x"77",
          5135 => x"84",
          5136 => x"39",
          5137 => x"52",
          5138 => x"86",
          5139 => x"84",
          5140 => x"55",
          5141 => x"08",
          5142 => x"c4",
          5143 => x"82",
          5144 => x"81",
          5145 => x"81",
          5146 => x"84",
          5147 => x"b0",
          5148 => x"84",
          5149 => x"51",
          5150 => x"82",
          5151 => x"a0",
          5152 => x"15",
          5153 => x"75",
          5154 => x"3f",
          5155 => x"08",
          5156 => x"76",
          5157 => x"77",
          5158 => x"9c",
          5159 => x"55",
          5160 => x"84",
          5161 => x"0d",
          5162 => x"0d",
          5163 => x"08",
          5164 => x"80",
          5165 => x"fc",
          5166 => x"93",
          5167 => x"82",
          5168 => x"80",
          5169 => x"93",
          5170 => x"98",
          5171 => x"78",
          5172 => x"3f",
          5173 => x"08",
          5174 => x"84",
          5175 => x"38",
          5176 => x"08",
          5177 => x"70",
          5178 => x"58",
          5179 => x"2e",
          5180 => x"83",
          5181 => x"82",
          5182 => x"55",
          5183 => x"81",
          5184 => x"07",
          5185 => x"2e",
          5186 => x"16",
          5187 => x"2e",
          5188 => x"88",
          5189 => x"82",
          5190 => x"56",
          5191 => x"51",
          5192 => x"82",
          5193 => x"54",
          5194 => x"08",
          5195 => x"9b",
          5196 => x"2e",
          5197 => x"83",
          5198 => x"73",
          5199 => x"0c",
          5200 => x"04",
          5201 => x"76",
          5202 => x"54",
          5203 => x"82",
          5204 => x"83",
          5205 => x"76",
          5206 => x"53",
          5207 => x"2e",
          5208 => x"90",
          5209 => x"51",
          5210 => x"82",
          5211 => x"90",
          5212 => x"53",
          5213 => x"84",
          5214 => x"0d",
          5215 => x"0d",
          5216 => x"83",
          5217 => x"54",
          5218 => x"55",
          5219 => x"3f",
          5220 => x"51",
          5221 => x"2e",
          5222 => x"8b",
          5223 => x"2a",
          5224 => x"51",
          5225 => x"86",
          5226 => x"f7",
          5227 => x"7d",
          5228 => x"75",
          5229 => x"98",
          5230 => x"2e",
          5231 => x"98",
          5232 => x"78",
          5233 => x"3f",
          5234 => x"08",
          5235 => x"84",
          5236 => x"38",
          5237 => x"70",
          5238 => x"73",
          5239 => x"58",
          5240 => x"8b",
          5241 => x"bf",
          5242 => x"ff",
          5243 => x"53",
          5244 => x"34",
          5245 => x"08",
          5246 => x"e5",
          5247 => x"81",
          5248 => x"2e",
          5249 => x"70",
          5250 => x"57",
          5251 => x"9e",
          5252 => x"2e",
          5253 => x"93",
          5254 => x"df",
          5255 => x"72",
          5256 => x"81",
          5257 => x"76",
          5258 => x"2e",
          5259 => x"52",
          5260 => x"fc",
          5261 => x"84",
          5262 => x"93",
          5263 => x"38",
          5264 => x"fe",
          5265 => x"39",
          5266 => x"16",
          5267 => x"93",
          5268 => x"3d",
          5269 => x"3d",
          5270 => x"08",
          5271 => x"52",
          5272 => x"c5",
          5273 => x"84",
          5274 => x"93",
          5275 => x"38",
          5276 => x"52",
          5277 => x"de",
          5278 => x"84",
          5279 => x"93",
          5280 => x"38",
          5281 => x"93",
          5282 => x"9c",
          5283 => x"ea",
          5284 => x"53",
          5285 => x"9c",
          5286 => x"ea",
          5287 => x"0b",
          5288 => x"74",
          5289 => x"0c",
          5290 => x"04",
          5291 => x"75",
          5292 => x"12",
          5293 => x"53",
          5294 => x"9a",
          5295 => x"84",
          5296 => x"9c",
          5297 => x"e5",
          5298 => x"0b",
          5299 => x"85",
          5300 => x"fa",
          5301 => x"7a",
          5302 => x"0b",
          5303 => x"98",
          5304 => x"2e",
          5305 => x"80",
          5306 => x"55",
          5307 => x"17",
          5308 => x"33",
          5309 => x"51",
          5310 => x"2e",
          5311 => x"85",
          5312 => x"06",
          5313 => x"e5",
          5314 => x"2e",
          5315 => x"8b",
          5316 => x"70",
          5317 => x"34",
          5318 => x"71",
          5319 => x"05",
          5320 => x"15",
          5321 => x"27",
          5322 => x"15",
          5323 => x"80",
          5324 => x"34",
          5325 => x"52",
          5326 => x"88",
          5327 => x"17",
          5328 => x"52",
          5329 => x"3f",
          5330 => x"08",
          5331 => x"12",
          5332 => x"3f",
          5333 => x"08",
          5334 => x"98",
          5335 => x"da",
          5336 => x"84",
          5337 => x"23",
          5338 => x"04",
          5339 => x"7f",
          5340 => x"5b",
          5341 => x"33",
          5342 => x"73",
          5343 => x"38",
          5344 => x"80",
          5345 => x"38",
          5346 => x"8c",
          5347 => x"08",
          5348 => x"aa",
          5349 => x"41",
          5350 => x"33",
          5351 => x"73",
          5352 => x"81",
          5353 => x"81",
          5354 => x"dc",
          5355 => x"70",
          5356 => x"07",
          5357 => x"73",
          5358 => x"88",
          5359 => x"70",
          5360 => x"73",
          5361 => x"38",
          5362 => x"ab",
          5363 => x"52",
          5364 => x"91",
          5365 => x"84",
          5366 => x"98",
          5367 => x"61",
          5368 => x"5a",
          5369 => x"a0",
          5370 => x"e7",
          5371 => x"70",
          5372 => x"79",
          5373 => x"73",
          5374 => x"81",
          5375 => x"38",
          5376 => x"33",
          5377 => x"ae",
          5378 => x"70",
          5379 => x"82",
          5380 => x"51",
          5381 => x"54",
          5382 => x"79",
          5383 => x"74",
          5384 => x"57",
          5385 => x"af",
          5386 => x"70",
          5387 => x"51",
          5388 => x"dc",
          5389 => x"73",
          5390 => x"38",
          5391 => x"82",
          5392 => x"19",
          5393 => x"54",
          5394 => x"82",
          5395 => x"54",
          5396 => x"78",
          5397 => x"81",
          5398 => x"54",
          5399 => x"81",
          5400 => x"af",
          5401 => x"77",
          5402 => x"70",
          5403 => x"25",
          5404 => x"07",
          5405 => x"51",
          5406 => x"2e",
          5407 => x"39",
          5408 => x"80",
          5409 => x"33",
          5410 => x"73",
          5411 => x"81",
          5412 => x"81",
          5413 => x"dc",
          5414 => x"70",
          5415 => x"07",
          5416 => x"73",
          5417 => x"b5",
          5418 => x"2e",
          5419 => x"83",
          5420 => x"76",
          5421 => x"07",
          5422 => x"2e",
          5423 => x"8b",
          5424 => x"77",
          5425 => x"30",
          5426 => x"71",
          5427 => x"53",
          5428 => x"55",
          5429 => x"38",
          5430 => x"5c",
          5431 => x"75",
          5432 => x"73",
          5433 => x"38",
          5434 => x"06",
          5435 => x"11",
          5436 => x"75",
          5437 => x"3f",
          5438 => x"08",
          5439 => x"38",
          5440 => x"33",
          5441 => x"54",
          5442 => x"e6",
          5443 => x"93",
          5444 => x"2e",
          5445 => x"ff",
          5446 => x"74",
          5447 => x"38",
          5448 => x"75",
          5449 => x"17",
          5450 => x"57",
          5451 => x"a7",
          5452 => x"81",
          5453 => x"e5",
          5454 => x"93",
          5455 => x"38",
          5456 => x"54",
          5457 => x"89",
          5458 => x"70",
          5459 => x"57",
          5460 => x"54",
          5461 => x"81",
          5462 => x"f7",
          5463 => x"7e",
          5464 => x"2e",
          5465 => x"33",
          5466 => x"e5",
          5467 => x"06",
          5468 => x"7a",
          5469 => x"a0",
          5470 => x"38",
          5471 => x"55",
          5472 => x"84",
          5473 => x"39",
          5474 => x"8b",
          5475 => x"7b",
          5476 => x"7a",
          5477 => x"3f",
          5478 => x"08",
          5479 => x"84",
          5480 => x"38",
          5481 => x"52",
          5482 => x"aa",
          5483 => x"84",
          5484 => x"93",
          5485 => x"c2",
          5486 => x"08",
          5487 => x"55",
          5488 => x"ff",
          5489 => x"15",
          5490 => x"54",
          5491 => x"34",
          5492 => x"70",
          5493 => x"81",
          5494 => x"58",
          5495 => x"8b",
          5496 => x"74",
          5497 => x"3f",
          5498 => x"08",
          5499 => x"38",
          5500 => x"51",
          5501 => x"ff",
          5502 => x"ab",
          5503 => x"55",
          5504 => x"bb",
          5505 => x"2e",
          5506 => x"80",
          5507 => x"85",
          5508 => x"06",
          5509 => x"58",
          5510 => x"80",
          5511 => x"75",
          5512 => x"73",
          5513 => x"b5",
          5514 => x"0b",
          5515 => x"80",
          5516 => x"39",
          5517 => x"54",
          5518 => x"85",
          5519 => x"75",
          5520 => x"81",
          5521 => x"73",
          5522 => x"1b",
          5523 => x"2a",
          5524 => x"51",
          5525 => x"80",
          5526 => x"90",
          5527 => x"ff",
          5528 => x"05",
          5529 => x"f5",
          5530 => x"93",
          5531 => x"1c",
          5532 => x"39",
          5533 => x"84",
          5534 => x"0d",
          5535 => x"0d",
          5536 => x"7b",
          5537 => x"73",
          5538 => x"55",
          5539 => x"2e",
          5540 => x"75",
          5541 => x"57",
          5542 => x"26",
          5543 => x"ba",
          5544 => x"70",
          5545 => x"ba",
          5546 => x"06",
          5547 => x"73",
          5548 => x"70",
          5549 => x"51",
          5550 => x"89",
          5551 => x"82",
          5552 => x"ff",
          5553 => x"56",
          5554 => x"2e",
          5555 => x"80",
          5556 => x"e0",
          5557 => x"08",
          5558 => x"76",
          5559 => x"58",
          5560 => x"81",
          5561 => x"ff",
          5562 => x"53",
          5563 => x"26",
          5564 => x"13",
          5565 => x"06",
          5566 => x"9f",
          5567 => x"99",
          5568 => x"e0",
          5569 => x"ff",
          5570 => x"72",
          5571 => x"2a",
          5572 => x"72",
          5573 => x"06",
          5574 => x"ff",
          5575 => x"30",
          5576 => x"70",
          5577 => x"07",
          5578 => x"9f",
          5579 => x"54",
          5580 => x"80",
          5581 => x"81",
          5582 => x"59",
          5583 => x"25",
          5584 => x"8b",
          5585 => x"24",
          5586 => x"76",
          5587 => x"78",
          5588 => x"82",
          5589 => x"51",
          5590 => x"84",
          5591 => x"0d",
          5592 => x"0d",
          5593 => x"0b",
          5594 => x"ff",
          5595 => x"0c",
          5596 => x"51",
          5597 => x"84",
          5598 => x"84",
          5599 => x"38",
          5600 => x"51",
          5601 => x"82",
          5602 => x"83",
          5603 => x"54",
          5604 => x"82",
          5605 => x"09",
          5606 => x"e3",
          5607 => x"b4",
          5608 => x"57",
          5609 => x"2e",
          5610 => x"83",
          5611 => x"74",
          5612 => x"70",
          5613 => x"25",
          5614 => x"51",
          5615 => x"38",
          5616 => x"2e",
          5617 => x"b5",
          5618 => x"81",
          5619 => x"80",
          5620 => x"e0",
          5621 => x"93",
          5622 => x"82",
          5623 => x"80",
          5624 => x"85",
          5625 => x"a4",
          5626 => x"16",
          5627 => x"3f",
          5628 => x"08",
          5629 => x"84",
          5630 => x"83",
          5631 => x"74",
          5632 => x"0c",
          5633 => x"04",
          5634 => x"61",
          5635 => x"80",
          5636 => x"58",
          5637 => x"0c",
          5638 => x"e1",
          5639 => x"84",
          5640 => x"56",
          5641 => x"93",
          5642 => x"86",
          5643 => x"93",
          5644 => x"29",
          5645 => x"05",
          5646 => x"53",
          5647 => x"80",
          5648 => x"38",
          5649 => x"76",
          5650 => x"74",
          5651 => x"72",
          5652 => x"38",
          5653 => x"51",
          5654 => x"82",
          5655 => x"81",
          5656 => x"81",
          5657 => x"72",
          5658 => x"80",
          5659 => x"38",
          5660 => x"70",
          5661 => x"53",
          5662 => x"86",
          5663 => x"a7",
          5664 => x"34",
          5665 => x"34",
          5666 => x"14",
          5667 => x"b2",
          5668 => x"84",
          5669 => x"06",
          5670 => x"54",
          5671 => x"72",
          5672 => x"76",
          5673 => x"38",
          5674 => x"70",
          5675 => x"53",
          5676 => x"85",
          5677 => x"70",
          5678 => x"5b",
          5679 => x"82",
          5680 => x"81",
          5681 => x"76",
          5682 => x"81",
          5683 => x"38",
          5684 => x"56",
          5685 => x"83",
          5686 => x"70",
          5687 => x"80",
          5688 => x"83",
          5689 => x"dc",
          5690 => x"93",
          5691 => x"76",
          5692 => x"05",
          5693 => x"16",
          5694 => x"56",
          5695 => x"d7",
          5696 => x"8d",
          5697 => x"72",
          5698 => x"54",
          5699 => x"57",
          5700 => x"95",
          5701 => x"73",
          5702 => x"3f",
          5703 => x"08",
          5704 => x"57",
          5705 => x"89",
          5706 => x"56",
          5707 => x"d7",
          5708 => x"76",
          5709 => x"f1",
          5710 => x"76",
          5711 => x"e9",
          5712 => x"51",
          5713 => x"82",
          5714 => x"83",
          5715 => x"53",
          5716 => x"2e",
          5717 => x"84",
          5718 => x"ca",
          5719 => x"da",
          5720 => x"84",
          5721 => x"ff",
          5722 => x"8d",
          5723 => x"14",
          5724 => x"3f",
          5725 => x"08",
          5726 => x"15",
          5727 => x"14",
          5728 => x"34",
          5729 => x"33",
          5730 => x"81",
          5731 => x"54",
          5732 => x"72",
          5733 => x"91",
          5734 => x"ff",
          5735 => x"29",
          5736 => x"33",
          5737 => x"72",
          5738 => x"72",
          5739 => x"38",
          5740 => x"06",
          5741 => x"2e",
          5742 => x"56",
          5743 => x"80",
          5744 => x"da",
          5745 => x"93",
          5746 => x"82",
          5747 => x"88",
          5748 => x"8f",
          5749 => x"56",
          5750 => x"38",
          5751 => x"51",
          5752 => x"82",
          5753 => x"83",
          5754 => x"55",
          5755 => x"80",
          5756 => x"da",
          5757 => x"93",
          5758 => x"80",
          5759 => x"da",
          5760 => x"93",
          5761 => x"ff",
          5762 => x"8d",
          5763 => x"2e",
          5764 => x"88",
          5765 => x"14",
          5766 => x"05",
          5767 => x"75",
          5768 => x"38",
          5769 => x"52",
          5770 => x"51",
          5771 => x"3f",
          5772 => x"08",
          5773 => x"84",
          5774 => x"82",
          5775 => x"93",
          5776 => x"ff",
          5777 => x"26",
          5778 => x"57",
          5779 => x"f5",
          5780 => x"82",
          5781 => x"f5",
          5782 => x"81",
          5783 => x"8d",
          5784 => x"2e",
          5785 => x"82",
          5786 => x"16",
          5787 => x"16",
          5788 => x"70",
          5789 => x"7a",
          5790 => x"0c",
          5791 => x"83",
          5792 => x"06",
          5793 => x"de",
          5794 => x"ae",
          5795 => x"84",
          5796 => x"ff",
          5797 => x"56",
          5798 => x"38",
          5799 => x"38",
          5800 => x"51",
          5801 => x"82",
          5802 => x"a8",
          5803 => x"82",
          5804 => x"39",
          5805 => x"80",
          5806 => x"38",
          5807 => x"15",
          5808 => x"53",
          5809 => x"8d",
          5810 => x"15",
          5811 => x"76",
          5812 => x"51",
          5813 => x"13",
          5814 => x"8d",
          5815 => x"15",
          5816 => x"c5",
          5817 => x"90",
          5818 => x"0b",
          5819 => x"ff",
          5820 => x"15",
          5821 => x"2e",
          5822 => x"81",
          5823 => x"e4",
          5824 => x"b6",
          5825 => x"84",
          5826 => x"ff",
          5827 => x"81",
          5828 => x"06",
          5829 => x"81",
          5830 => x"51",
          5831 => x"82",
          5832 => x"80",
          5833 => x"93",
          5834 => x"15",
          5835 => x"14",
          5836 => x"3f",
          5837 => x"08",
          5838 => x"06",
          5839 => x"d4",
          5840 => x"81",
          5841 => x"38",
          5842 => x"d8",
          5843 => x"93",
          5844 => x"8b",
          5845 => x"2e",
          5846 => x"b3",
          5847 => x"14",
          5848 => x"3f",
          5849 => x"08",
          5850 => x"e4",
          5851 => x"81",
          5852 => x"84",
          5853 => x"d7",
          5854 => x"93",
          5855 => x"15",
          5856 => x"14",
          5857 => x"3f",
          5858 => x"08",
          5859 => x"76",
          5860 => x"93",
          5861 => x"05",
          5862 => x"93",
          5863 => x"86",
          5864 => x"0b",
          5865 => x"80",
          5866 => x"93",
          5867 => x"3d",
          5868 => x"3d",
          5869 => x"89",
          5870 => x"2e",
          5871 => x"08",
          5872 => x"2e",
          5873 => x"33",
          5874 => x"2e",
          5875 => x"13",
          5876 => x"22",
          5877 => x"76",
          5878 => x"06",
          5879 => x"13",
          5880 => x"c0",
          5881 => x"84",
          5882 => x"52",
          5883 => x"71",
          5884 => x"55",
          5885 => x"53",
          5886 => x"0c",
          5887 => x"93",
          5888 => x"3d",
          5889 => x"3d",
          5890 => x"05",
          5891 => x"89",
          5892 => x"52",
          5893 => x"3f",
          5894 => x"0b",
          5895 => x"08",
          5896 => x"82",
          5897 => x"84",
          5898 => x"b4",
          5899 => x"55",
          5900 => x"2e",
          5901 => x"74",
          5902 => x"73",
          5903 => x"38",
          5904 => x"78",
          5905 => x"54",
          5906 => x"92",
          5907 => x"89",
          5908 => x"84",
          5909 => x"b0",
          5910 => x"84",
          5911 => x"82",
          5912 => x"88",
          5913 => x"eb",
          5914 => x"02",
          5915 => x"e7",
          5916 => x"59",
          5917 => x"80",
          5918 => x"38",
          5919 => x"70",
          5920 => x"d0",
          5921 => x"3d",
          5922 => x"58",
          5923 => x"82",
          5924 => x"55",
          5925 => x"08",
          5926 => x"7a",
          5927 => x"8c",
          5928 => x"56",
          5929 => x"82",
          5930 => x"55",
          5931 => x"08",
          5932 => x"80",
          5933 => x"70",
          5934 => x"57",
          5935 => x"83",
          5936 => x"77",
          5937 => x"73",
          5938 => x"ab",
          5939 => x"2e",
          5940 => x"84",
          5941 => x"06",
          5942 => x"51",
          5943 => x"82",
          5944 => x"55",
          5945 => x"b2",
          5946 => x"06",
          5947 => x"b8",
          5948 => x"2a",
          5949 => x"51",
          5950 => x"2e",
          5951 => x"55",
          5952 => x"77",
          5953 => x"74",
          5954 => x"77",
          5955 => x"81",
          5956 => x"73",
          5957 => x"af",
          5958 => x"7a",
          5959 => x"3f",
          5960 => x"08",
          5961 => x"b2",
          5962 => x"8e",
          5963 => x"ea",
          5964 => x"a0",
          5965 => x"34",
          5966 => x"52",
          5967 => x"bd",
          5968 => x"62",
          5969 => x"d4",
          5970 => x"54",
          5971 => x"15",
          5972 => x"2e",
          5973 => x"7a",
          5974 => x"51",
          5975 => x"75",
          5976 => x"d4",
          5977 => x"be",
          5978 => x"84",
          5979 => x"93",
          5980 => x"ca",
          5981 => x"74",
          5982 => x"02",
          5983 => x"70",
          5984 => x"81",
          5985 => x"56",
          5986 => x"86",
          5987 => x"82",
          5988 => x"81",
          5989 => x"06",
          5990 => x"80",
          5991 => x"75",
          5992 => x"73",
          5993 => x"38",
          5994 => x"92",
          5995 => x"7a",
          5996 => x"3f",
          5997 => x"08",
          5998 => x"8c",
          5999 => x"55",
          6000 => x"08",
          6001 => x"77",
          6002 => x"81",
          6003 => x"73",
          6004 => x"38",
          6005 => x"07",
          6006 => x"11",
          6007 => x"0c",
          6008 => x"0c",
          6009 => x"52",
          6010 => x"3f",
          6011 => x"08",
          6012 => x"08",
          6013 => x"63",
          6014 => x"5a",
          6015 => x"82",
          6016 => x"82",
          6017 => x"8c",
          6018 => x"7a",
          6019 => x"17",
          6020 => x"23",
          6021 => x"34",
          6022 => x"1a",
          6023 => x"9c",
          6024 => x"0b",
          6025 => x"77",
          6026 => x"81",
          6027 => x"73",
          6028 => x"8d",
          6029 => x"84",
          6030 => x"81",
          6031 => x"93",
          6032 => x"1a",
          6033 => x"22",
          6034 => x"7b",
          6035 => x"a8",
          6036 => x"78",
          6037 => x"3f",
          6038 => x"08",
          6039 => x"84",
          6040 => x"83",
          6041 => x"82",
          6042 => x"ff",
          6043 => x"06",
          6044 => x"55",
          6045 => x"56",
          6046 => x"76",
          6047 => x"51",
          6048 => x"27",
          6049 => x"70",
          6050 => x"5a",
          6051 => x"76",
          6052 => x"74",
          6053 => x"83",
          6054 => x"73",
          6055 => x"38",
          6056 => x"51",
          6057 => x"82",
          6058 => x"85",
          6059 => x"8e",
          6060 => x"2a",
          6061 => x"08",
          6062 => x"0c",
          6063 => x"79",
          6064 => x"73",
          6065 => x"0c",
          6066 => x"04",
          6067 => x"60",
          6068 => x"40",
          6069 => x"80",
          6070 => x"3d",
          6071 => x"78",
          6072 => x"3f",
          6073 => x"08",
          6074 => x"84",
          6075 => x"91",
          6076 => x"74",
          6077 => x"38",
          6078 => x"c4",
          6079 => x"33",
          6080 => x"87",
          6081 => x"2e",
          6082 => x"95",
          6083 => x"91",
          6084 => x"56",
          6085 => x"81",
          6086 => x"34",
          6087 => x"a0",
          6088 => x"08",
          6089 => x"31",
          6090 => x"27",
          6091 => x"5c",
          6092 => x"82",
          6093 => x"19",
          6094 => x"ff",
          6095 => x"74",
          6096 => x"7e",
          6097 => x"ff",
          6098 => x"2a",
          6099 => x"79",
          6100 => x"87",
          6101 => x"08",
          6102 => x"98",
          6103 => x"78",
          6104 => x"3f",
          6105 => x"08",
          6106 => x"27",
          6107 => x"74",
          6108 => x"a3",
          6109 => x"1a",
          6110 => x"08",
          6111 => x"d4",
          6112 => x"93",
          6113 => x"2e",
          6114 => x"82",
          6115 => x"1a",
          6116 => x"59",
          6117 => x"2e",
          6118 => x"77",
          6119 => x"11",
          6120 => x"55",
          6121 => x"85",
          6122 => x"31",
          6123 => x"76",
          6124 => x"81",
          6125 => x"ca",
          6126 => x"93",
          6127 => x"d7",
          6128 => x"11",
          6129 => x"74",
          6130 => x"38",
          6131 => x"77",
          6132 => x"78",
          6133 => x"84",
          6134 => x"16",
          6135 => x"08",
          6136 => x"2b",
          6137 => x"cf",
          6138 => x"89",
          6139 => x"39",
          6140 => x"0c",
          6141 => x"83",
          6142 => x"80",
          6143 => x"55",
          6144 => x"83",
          6145 => x"9c",
          6146 => x"7e",
          6147 => x"3f",
          6148 => x"08",
          6149 => x"75",
          6150 => x"08",
          6151 => x"1f",
          6152 => x"7c",
          6153 => x"3f",
          6154 => x"7e",
          6155 => x"0c",
          6156 => x"1b",
          6157 => x"1c",
          6158 => x"fd",
          6159 => x"56",
          6160 => x"84",
          6161 => x"0d",
          6162 => x"0d",
          6163 => x"64",
          6164 => x"58",
          6165 => x"90",
          6166 => x"52",
          6167 => x"d2",
          6168 => x"84",
          6169 => x"93",
          6170 => x"38",
          6171 => x"55",
          6172 => x"86",
          6173 => x"83",
          6174 => x"18",
          6175 => x"2a",
          6176 => x"51",
          6177 => x"56",
          6178 => x"83",
          6179 => x"39",
          6180 => x"19",
          6181 => x"83",
          6182 => x"0b",
          6183 => x"81",
          6184 => x"39",
          6185 => x"7c",
          6186 => x"74",
          6187 => x"38",
          6188 => x"7b",
          6189 => x"ec",
          6190 => x"08",
          6191 => x"06",
          6192 => x"81",
          6193 => x"8a",
          6194 => x"05",
          6195 => x"06",
          6196 => x"bf",
          6197 => x"38",
          6198 => x"55",
          6199 => x"7a",
          6200 => x"98",
          6201 => x"77",
          6202 => x"3f",
          6203 => x"08",
          6204 => x"84",
          6205 => x"82",
          6206 => x"81",
          6207 => x"38",
          6208 => x"ff",
          6209 => x"98",
          6210 => x"18",
          6211 => x"74",
          6212 => x"7e",
          6213 => x"08",
          6214 => x"2e",
          6215 => x"8d",
          6216 => x"ce",
          6217 => x"93",
          6218 => x"ee",
          6219 => x"08",
          6220 => x"d1",
          6221 => x"93",
          6222 => x"2e",
          6223 => x"82",
          6224 => x"1b",
          6225 => x"5a",
          6226 => x"2e",
          6227 => x"78",
          6228 => x"11",
          6229 => x"55",
          6230 => x"85",
          6231 => x"31",
          6232 => x"76",
          6233 => x"81",
          6234 => x"c8",
          6235 => x"93",
          6236 => x"a6",
          6237 => x"11",
          6238 => x"56",
          6239 => x"27",
          6240 => x"80",
          6241 => x"08",
          6242 => x"2b",
          6243 => x"b4",
          6244 => x"b5",
          6245 => x"80",
          6246 => x"34",
          6247 => x"56",
          6248 => x"8c",
          6249 => x"19",
          6250 => x"38",
          6251 => x"b6",
          6252 => x"84",
          6253 => x"38",
          6254 => x"12",
          6255 => x"9c",
          6256 => x"18",
          6257 => x"06",
          6258 => x"31",
          6259 => x"76",
          6260 => x"7b",
          6261 => x"08",
          6262 => x"cd",
          6263 => x"93",
          6264 => x"b6",
          6265 => x"7c",
          6266 => x"08",
          6267 => x"1f",
          6268 => x"cb",
          6269 => x"55",
          6270 => x"16",
          6271 => x"31",
          6272 => x"7f",
          6273 => x"94",
          6274 => x"70",
          6275 => x"8c",
          6276 => x"58",
          6277 => x"76",
          6278 => x"75",
          6279 => x"19",
          6280 => x"39",
          6281 => x"80",
          6282 => x"74",
          6283 => x"80",
          6284 => x"93",
          6285 => x"3d",
          6286 => x"3d",
          6287 => x"3d",
          6288 => x"70",
          6289 => x"ea",
          6290 => x"84",
          6291 => x"93",
          6292 => x"fb",
          6293 => x"33",
          6294 => x"70",
          6295 => x"55",
          6296 => x"2e",
          6297 => x"a0",
          6298 => x"78",
          6299 => x"3f",
          6300 => x"08",
          6301 => x"84",
          6302 => x"38",
          6303 => x"8b",
          6304 => x"07",
          6305 => x"8b",
          6306 => x"16",
          6307 => x"52",
          6308 => x"dd",
          6309 => x"16",
          6310 => x"15",
          6311 => x"3f",
          6312 => x"0a",
          6313 => x"51",
          6314 => x"76",
          6315 => x"51",
          6316 => x"78",
          6317 => x"83",
          6318 => x"51",
          6319 => x"82",
          6320 => x"90",
          6321 => x"bf",
          6322 => x"73",
          6323 => x"76",
          6324 => x"0c",
          6325 => x"04",
          6326 => x"76",
          6327 => x"fe",
          6328 => x"93",
          6329 => x"82",
          6330 => x"9c",
          6331 => x"fc",
          6332 => x"51",
          6333 => x"82",
          6334 => x"53",
          6335 => x"08",
          6336 => x"93",
          6337 => x"0c",
          6338 => x"84",
          6339 => x"0d",
          6340 => x"0d",
          6341 => x"e6",
          6342 => x"52",
          6343 => x"93",
          6344 => x"8b",
          6345 => x"84",
          6346 => x"c8",
          6347 => x"71",
          6348 => x"0c",
          6349 => x"04",
          6350 => x"80",
          6351 => x"d0",
          6352 => x"3d",
          6353 => x"3f",
          6354 => x"08",
          6355 => x"84",
          6356 => x"38",
          6357 => x"52",
          6358 => x"05",
          6359 => x"3f",
          6360 => x"08",
          6361 => x"84",
          6362 => x"02",
          6363 => x"33",
          6364 => x"55",
          6365 => x"25",
          6366 => x"7a",
          6367 => x"54",
          6368 => x"a2",
          6369 => x"84",
          6370 => x"06",
          6371 => x"73",
          6372 => x"38",
          6373 => x"70",
          6374 => x"a8",
          6375 => x"84",
          6376 => x"0c",
          6377 => x"93",
          6378 => x"2e",
          6379 => x"83",
          6380 => x"74",
          6381 => x"0c",
          6382 => x"04",
          6383 => x"6f",
          6384 => x"80",
          6385 => x"53",
          6386 => x"b8",
          6387 => x"3d",
          6388 => x"3f",
          6389 => x"08",
          6390 => x"84",
          6391 => x"38",
          6392 => x"7c",
          6393 => x"47",
          6394 => x"54",
          6395 => x"81",
          6396 => x"52",
          6397 => x"52",
          6398 => x"3f",
          6399 => x"08",
          6400 => x"84",
          6401 => x"38",
          6402 => x"51",
          6403 => x"82",
          6404 => x"57",
          6405 => x"08",
          6406 => x"69",
          6407 => x"da",
          6408 => x"93",
          6409 => x"76",
          6410 => x"d5",
          6411 => x"93",
          6412 => x"82",
          6413 => x"82",
          6414 => x"52",
          6415 => x"eb",
          6416 => x"84",
          6417 => x"93",
          6418 => x"38",
          6419 => x"51",
          6420 => x"73",
          6421 => x"08",
          6422 => x"76",
          6423 => x"d6",
          6424 => x"93",
          6425 => x"82",
          6426 => x"80",
          6427 => x"76",
          6428 => x"81",
          6429 => x"82",
          6430 => x"39",
          6431 => x"38",
          6432 => x"bc",
          6433 => x"51",
          6434 => x"76",
          6435 => x"11",
          6436 => x"51",
          6437 => x"73",
          6438 => x"38",
          6439 => x"55",
          6440 => x"16",
          6441 => x"56",
          6442 => x"38",
          6443 => x"73",
          6444 => x"90",
          6445 => x"2e",
          6446 => x"16",
          6447 => x"ff",
          6448 => x"ff",
          6449 => x"58",
          6450 => x"74",
          6451 => x"75",
          6452 => x"18",
          6453 => x"58",
          6454 => x"fe",
          6455 => x"7b",
          6456 => x"06",
          6457 => x"18",
          6458 => x"58",
          6459 => x"80",
          6460 => x"c8",
          6461 => x"29",
          6462 => x"05",
          6463 => x"33",
          6464 => x"56",
          6465 => x"2e",
          6466 => x"16",
          6467 => x"33",
          6468 => x"73",
          6469 => x"16",
          6470 => x"26",
          6471 => x"55",
          6472 => x"91",
          6473 => x"54",
          6474 => x"70",
          6475 => x"34",
          6476 => x"ec",
          6477 => x"70",
          6478 => x"34",
          6479 => x"09",
          6480 => x"38",
          6481 => x"39",
          6482 => x"19",
          6483 => x"33",
          6484 => x"05",
          6485 => x"78",
          6486 => x"80",
          6487 => x"82",
          6488 => x"9e",
          6489 => x"f7",
          6490 => x"7d",
          6491 => x"05",
          6492 => x"57",
          6493 => x"3f",
          6494 => x"08",
          6495 => x"84",
          6496 => x"38",
          6497 => x"53",
          6498 => x"38",
          6499 => x"54",
          6500 => x"92",
          6501 => x"33",
          6502 => x"70",
          6503 => x"54",
          6504 => x"38",
          6505 => x"15",
          6506 => x"70",
          6507 => x"58",
          6508 => x"82",
          6509 => x"8a",
          6510 => x"89",
          6511 => x"53",
          6512 => x"b7",
          6513 => x"ff",
          6514 => x"ff",
          6515 => x"93",
          6516 => x"15",
          6517 => x"53",
          6518 => x"fe",
          6519 => x"93",
          6520 => x"26",
          6521 => x"30",
          6522 => x"70",
          6523 => x"77",
          6524 => x"18",
          6525 => x"51",
          6526 => x"88",
          6527 => x"73",
          6528 => x"52",
          6529 => x"ca",
          6530 => x"84",
          6531 => x"93",
          6532 => x"2e",
          6533 => x"82",
          6534 => x"ff",
          6535 => x"38",
          6536 => x"08",
          6537 => x"73",
          6538 => x"73",
          6539 => x"9c",
          6540 => x"27",
          6541 => x"75",
          6542 => x"16",
          6543 => x"17",
          6544 => x"33",
          6545 => x"70",
          6546 => x"55",
          6547 => x"80",
          6548 => x"73",
          6549 => x"cc",
          6550 => x"93",
          6551 => x"82",
          6552 => x"94",
          6553 => x"84",
          6554 => x"39",
          6555 => x"51",
          6556 => x"82",
          6557 => x"54",
          6558 => x"be",
          6559 => x"27",
          6560 => x"53",
          6561 => x"08",
          6562 => x"73",
          6563 => x"ff",
          6564 => x"15",
          6565 => x"16",
          6566 => x"ff",
          6567 => x"80",
          6568 => x"73",
          6569 => x"c6",
          6570 => x"93",
          6571 => x"38",
          6572 => x"16",
          6573 => x"80",
          6574 => x"0b",
          6575 => x"81",
          6576 => x"75",
          6577 => x"93",
          6578 => x"58",
          6579 => x"54",
          6580 => x"74",
          6581 => x"73",
          6582 => x"90",
          6583 => x"c0",
          6584 => x"90",
          6585 => x"83",
          6586 => x"72",
          6587 => x"38",
          6588 => x"08",
          6589 => x"77",
          6590 => x"80",
          6591 => x"93",
          6592 => x"3d",
          6593 => x"3d",
          6594 => x"89",
          6595 => x"2e",
          6596 => x"80",
          6597 => x"fc",
          6598 => x"3d",
          6599 => x"e1",
          6600 => x"93",
          6601 => x"82",
          6602 => x"80",
          6603 => x"76",
          6604 => x"75",
          6605 => x"3f",
          6606 => x"08",
          6607 => x"84",
          6608 => x"38",
          6609 => x"70",
          6610 => x"57",
          6611 => x"a2",
          6612 => x"33",
          6613 => x"70",
          6614 => x"55",
          6615 => x"2e",
          6616 => x"16",
          6617 => x"51",
          6618 => x"82",
          6619 => x"88",
          6620 => x"54",
          6621 => x"84",
          6622 => x"52",
          6623 => x"e5",
          6624 => x"84",
          6625 => x"84",
          6626 => x"06",
          6627 => x"55",
          6628 => x"80",
          6629 => x"80",
          6630 => x"54",
          6631 => x"84",
          6632 => x"0d",
          6633 => x"0d",
          6634 => x"fc",
          6635 => x"52",
          6636 => x"3f",
          6637 => x"08",
          6638 => x"93",
          6639 => x"0c",
          6640 => x"04",
          6641 => x"77",
          6642 => x"fc",
          6643 => x"53",
          6644 => x"de",
          6645 => x"84",
          6646 => x"93",
          6647 => x"df",
          6648 => x"38",
          6649 => x"08",
          6650 => x"cd",
          6651 => x"93",
          6652 => x"80",
          6653 => x"93",
          6654 => x"73",
          6655 => x"3f",
          6656 => x"08",
          6657 => x"84",
          6658 => x"09",
          6659 => x"38",
          6660 => x"39",
          6661 => x"08",
          6662 => x"52",
          6663 => x"b3",
          6664 => x"73",
          6665 => x"3f",
          6666 => x"08",
          6667 => x"30",
          6668 => x"9f",
          6669 => x"93",
          6670 => x"51",
          6671 => x"72",
          6672 => x"0c",
          6673 => x"04",
          6674 => x"65",
          6675 => x"89",
          6676 => x"96",
          6677 => x"df",
          6678 => x"93",
          6679 => x"82",
          6680 => x"b2",
          6681 => x"75",
          6682 => x"3f",
          6683 => x"08",
          6684 => x"84",
          6685 => x"02",
          6686 => x"33",
          6687 => x"55",
          6688 => x"25",
          6689 => x"55",
          6690 => x"80",
          6691 => x"76",
          6692 => x"d4",
          6693 => x"82",
          6694 => x"94",
          6695 => x"f0",
          6696 => x"65",
          6697 => x"53",
          6698 => x"05",
          6699 => x"51",
          6700 => x"82",
          6701 => x"5b",
          6702 => x"08",
          6703 => x"7c",
          6704 => x"08",
          6705 => x"fe",
          6706 => x"08",
          6707 => x"55",
          6708 => x"91",
          6709 => x"0c",
          6710 => x"81",
          6711 => x"39",
          6712 => x"c7",
          6713 => x"84",
          6714 => x"55",
          6715 => x"2e",
          6716 => x"bf",
          6717 => x"5f",
          6718 => x"92",
          6719 => x"51",
          6720 => x"82",
          6721 => x"ff",
          6722 => x"82",
          6723 => x"81",
          6724 => x"82",
          6725 => x"30",
          6726 => x"84",
          6727 => x"25",
          6728 => x"19",
          6729 => x"5a",
          6730 => x"08",
          6731 => x"38",
          6732 => x"a4",
          6733 => x"93",
          6734 => x"58",
          6735 => x"77",
          6736 => x"7d",
          6737 => x"bf",
          6738 => x"93",
          6739 => x"82",
          6740 => x"80",
          6741 => x"70",
          6742 => x"ff",
          6743 => x"56",
          6744 => x"2e",
          6745 => x"9e",
          6746 => x"51",
          6747 => x"3f",
          6748 => x"08",
          6749 => x"06",
          6750 => x"80",
          6751 => x"19",
          6752 => x"54",
          6753 => x"14",
          6754 => x"c5",
          6755 => x"84",
          6756 => x"06",
          6757 => x"80",
          6758 => x"19",
          6759 => x"54",
          6760 => x"06",
          6761 => x"79",
          6762 => x"78",
          6763 => x"79",
          6764 => x"84",
          6765 => x"07",
          6766 => x"84",
          6767 => x"82",
          6768 => x"92",
          6769 => x"f9",
          6770 => x"8a",
          6771 => x"53",
          6772 => x"e3",
          6773 => x"93",
          6774 => x"82",
          6775 => x"81",
          6776 => x"17",
          6777 => x"81",
          6778 => x"17",
          6779 => x"2a",
          6780 => x"51",
          6781 => x"55",
          6782 => x"81",
          6783 => x"17",
          6784 => x"8c",
          6785 => x"81",
          6786 => x"9b",
          6787 => x"84",
          6788 => x"17",
          6789 => x"51",
          6790 => x"82",
          6791 => x"74",
          6792 => x"56",
          6793 => x"98",
          6794 => x"76",
          6795 => x"c6",
          6796 => x"84",
          6797 => x"09",
          6798 => x"38",
          6799 => x"93",
          6800 => x"2e",
          6801 => x"85",
          6802 => x"a3",
          6803 => x"38",
          6804 => x"93",
          6805 => x"15",
          6806 => x"38",
          6807 => x"53",
          6808 => x"08",
          6809 => x"c3",
          6810 => x"93",
          6811 => x"94",
          6812 => x"18",
          6813 => x"33",
          6814 => x"54",
          6815 => x"34",
          6816 => x"85",
          6817 => x"18",
          6818 => x"74",
          6819 => x"0c",
          6820 => x"04",
          6821 => x"82",
          6822 => x"ff",
          6823 => x"a1",
          6824 => x"e4",
          6825 => x"84",
          6826 => x"93",
          6827 => x"f5",
          6828 => x"a1",
          6829 => x"95",
          6830 => x"58",
          6831 => x"82",
          6832 => x"55",
          6833 => x"08",
          6834 => x"02",
          6835 => x"33",
          6836 => x"70",
          6837 => x"55",
          6838 => x"73",
          6839 => x"75",
          6840 => x"80",
          6841 => x"bd",
          6842 => x"d6",
          6843 => x"81",
          6844 => x"87",
          6845 => x"ad",
          6846 => x"78",
          6847 => x"3f",
          6848 => x"08",
          6849 => x"70",
          6850 => x"55",
          6851 => x"2e",
          6852 => x"78",
          6853 => x"84",
          6854 => x"08",
          6855 => x"38",
          6856 => x"93",
          6857 => x"76",
          6858 => x"70",
          6859 => x"b5",
          6860 => x"84",
          6861 => x"93",
          6862 => x"e9",
          6863 => x"84",
          6864 => x"51",
          6865 => x"82",
          6866 => x"55",
          6867 => x"08",
          6868 => x"55",
          6869 => x"82",
          6870 => x"84",
          6871 => x"82",
          6872 => x"80",
          6873 => x"51",
          6874 => x"82",
          6875 => x"82",
          6876 => x"30",
          6877 => x"84",
          6878 => x"25",
          6879 => x"75",
          6880 => x"38",
          6881 => x"8f",
          6882 => x"75",
          6883 => x"c1",
          6884 => x"93",
          6885 => x"74",
          6886 => x"51",
          6887 => x"3f",
          6888 => x"08",
          6889 => x"93",
          6890 => x"3d",
          6891 => x"3d",
          6892 => x"99",
          6893 => x"52",
          6894 => x"d8",
          6895 => x"93",
          6896 => x"82",
          6897 => x"82",
          6898 => x"5e",
          6899 => x"3d",
          6900 => x"cf",
          6901 => x"93",
          6902 => x"82",
          6903 => x"86",
          6904 => x"82",
          6905 => x"93",
          6906 => x"2e",
          6907 => x"82",
          6908 => x"80",
          6909 => x"70",
          6910 => x"06",
          6911 => x"54",
          6912 => x"38",
          6913 => x"52",
          6914 => x"52",
          6915 => x"3f",
          6916 => x"08",
          6917 => x"82",
          6918 => x"83",
          6919 => x"82",
          6920 => x"81",
          6921 => x"06",
          6922 => x"54",
          6923 => x"08",
          6924 => x"81",
          6925 => x"81",
          6926 => x"39",
          6927 => x"38",
          6928 => x"08",
          6929 => x"c4",
          6930 => x"93",
          6931 => x"82",
          6932 => x"81",
          6933 => x"53",
          6934 => x"19",
          6935 => x"8c",
          6936 => x"ae",
          6937 => x"34",
          6938 => x"0b",
          6939 => x"82",
          6940 => x"52",
          6941 => x"51",
          6942 => x"3f",
          6943 => x"b4",
          6944 => x"c9",
          6945 => x"53",
          6946 => x"53",
          6947 => x"51",
          6948 => x"3f",
          6949 => x"0b",
          6950 => x"34",
          6951 => x"80",
          6952 => x"51",
          6953 => x"78",
          6954 => x"83",
          6955 => x"51",
          6956 => x"82",
          6957 => x"54",
          6958 => x"08",
          6959 => x"88",
          6960 => x"64",
          6961 => x"ff",
          6962 => x"75",
          6963 => x"78",
          6964 => x"3f",
          6965 => x"0b",
          6966 => x"78",
          6967 => x"83",
          6968 => x"51",
          6969 => x"3f",
          6970 => x"08",
          6971 => x"80",
          6972 => x"76",
          6973 => x"ae",
          6974 => x"93",
          6975 => x"3d",
          6976 => x"3d",
          6977 => x"84",
          6978 => x"f1",
          6979 => x"a8",
          6980 => x"05",
          6981 => x"51",
          6982 => x"82",
          6983 => x"55",
          6984 => x"08",
          6985 => x"78",
          6986 => x"08",
          6987 => x"70",
          6988 => x"b8",
          6989 => x"84",
          6990 => x"93",
          6991 => x"b9",
          6992 => x"9b",
          6993 => x"a0",
          6994 => x"55",
          6995 => x"38",
          6996 => x"3d",
          6997 => x"3d",
          6998 => x"51",
          6999 => x"3f",
          7000 => x"52",
          7001 => x"52",
          7002 => x"dd",
          7003 => x"08",
          7004 => x"cb",
          7005 => x"93",
          7006 => x"82",
          7007 => x"95",
          7008 => x"2e",
          7009 => x"88",
          7010 => x"3d",
          7011 => x"38",
          7012 => x"e5",
          7013 => x"84",
          7014 => x"09",
          7015 => x"b8",
          7016 => x"c9",
          7017 => x"93",
          7018 => x"82",
          7019 => x"81",
          7020 => x"56",
          7021 => x"3d",
          7022 => x"52",
          7023 => x"ff",
          7024 => x"02",
          7025 => x"8b",
          7026 => x"16",
          7027 => x"2a",
          7028 => x"51",
          7029 => x"89",
          7030 => x"07",
          7031 => x"17",
          7032 => x"81",
          7033 => x"34",
          7034 => x"70",
          7035 => x"81",
          7036 => x"55",
          7037 => x"80",
          7038 => x"64",
          7039 => x"38",
          7040 => x"51",
          7041 => x"82",
          7042 => x"52",
          7043 => x"b7",
          7044 => x"55",
          7045 => x"08",
          7046 => x"dd",
          7047 => x"84",
          7048 => x"51",
          7049 => x"3f",
          7050 => x"08",
          7051 => x"11",
          7052 => x"82",
          7053 => x"80",
          7054 => x"16",
          7055 => x"ae",
          7056 => x"06",
          7057 => x"53",
          7058 => x"51",
          7059 => x"78",
          7060 => x"83",
          7061 => x"39",
          7062 => x"08",
          7063 => x"51",
          7064 => x"82",
          7065 => x"55",
          7066 => x"08",
          7067 => x"51",
          7068 => x"3f",
          7069 => x"08",
          7070 => x"93",
          7071 => x"3d",
          7072 => x"3d",
          7073 => x"db",
          7074 => x"84",
          7075 => x"05",
          7076 => x"82",
          7077 => x"d0",
          7078 => x"3d",
          7079 => x"3f",
          7080 => x"08",
          7081 => x"84",
          7082 => x"38",
          7083 => x"52",
          7084 => x"05",
          7085 => x"3f",
          7086 => x"08",
          7087 => x"84",
          7088 => x"02",
          7089 => x"33",
          7090 => x"54",
          7091 => x"aa",
          7092 => x"06",
          7093 => x"8b",
          7094 => x"06",
          7095 => x"07",
          7096 => x"56",
          7097 => x"34",
          7098 => x"0b",
          7099 => x"78",
          7100 => x"a9",
          7101 => x"84",
          7102 => x"82",
          7103 => x"95",
          7104 => x"ef",
          7105 => x"56",
          7106 => x"3d",
          7107 => x"94",
          7108 => x"f4",
          7109 => x"84",
          7110 => x"93",
          7111 => x"cb",
          7112 => x"63",
          7113 => x"d4",
          7114 => x"c0",
          7115 => x"84",
          7116 => x"93",
          7117 => x"38",
          7118 => x"05",
          7119 => x"06",
          7120 => x"73",
          7121 => x"16",
          7122 => x"22",
          7123 => x"07",
          7124 => x"1f",
          7125 => x"c2",
          7126 => x"81",
          7127 => x"34",
          7128 => x"b3",
          7129 => x"93",
          7130 => x"74",
          7131 => x"0c",
          7132 => x"04",
          7133 => x"69",
          7134 => x"80",
          7135 => x"d0",
          7136 => x"3d",
          7137 => x"3f",
          7138 => x"08",
          7139 => x"08",
          7140 => x"93",
          7141 => x"80",
          7142 => x"57",
          7143 => x"81",
          7144 => x"70",
          7145 => x"55",
          7146 => x"80",
          7147 => x"5d",
          7148 => x"52",
          7149 => x"52",
          7150 => x"a9",
          7151 => x"84",
          7152 => x"93",
          7153 => x"d1",
          7154 => x"73",
          7155 => x"3f",
          7156 => x"08",
          7157 => x"84",
          7158 => x"82",
          7159 => x"82",
          7160 => x"65",
          7161 => x"78",
          7162 => x"7b",
          7163 => x"55",
          7164 => x"34",
          7165 => x"8a",
          7166 => x"38",
          7167 => x"1a",
          7168 => x"34",
          7169 => x"9e",
          7170 => x"70",
          7171 => x"51",
          7172 => x"a0",
          7173 => x"8e",
          7174 => x"2e",
          7175 => x"86",
          7176 => x"34",
          7177 => x"30",
          7178 => x"80",
          7179 => x"7a",
          7180 => x"c1",
          7181 => x"2e",
          7182 => x"a0",
          7183 => x"51",
          7184 => x"3f",
          7185 => x"08",
          7186 => x"84",
          7187 => x"7b",
          7188 => x"55",
          7189 => x"73",
          7190 => x"38",
          7191 => x"73",
          7192 => x"38",
          7193 => x"15",
          7194 => x"ff",
          7195 => x"82",
          7196 => x"7b",
          7197 => x"93",
          7198 => x"3d",
          7199 => x"3d",
          7200 => x"9c",
          7201 => x"05",
          7202 => x"51",
          7203 => x"82",
          7204 => x"82",
          7205 => x"56",
          7206 => x"84",
          7207 => x"38",
          7208 => x"52",
          7209 => x"52",
          7210 => x"c0",
          7211 => x"70",
          7212 => x"ff",
          7213 => x"55",
          7214 => x"27",
          7215 => x"78",
          7216 => x"ff",
          7217 => x"05",
          7218 => x"55",
          7219 => x"3f",
          7220 => x"08",
          7221 => x"38",
          7222 => x"70",
          7223 => x"ff",
          7224 => x"82",
          7225 => x"80",
          7226 => x"74",
          7227 => x"07",
          7228 => x"4e",
          7229 => x"82",
          7230 => x"55",
          7231 => x"70",
          7232 => x"06",
          7233 => x"99",
          7234 => x"e0",
          7235 => x"ff",
          7236 => x"54",
          7237 => x"27",
          7238 => x"fe",
          7239 => x"55",
          7240 => x"a3",
          7241 => x"82",
          7242 => x"ff",
          7243 => x"82",
          7244 => x"93",
          7245 => x"75",
          7246 => x"76",
          7247 => x"38",
          7248 => x"77",
          7249 => x"86",
          7250 => x"39",
          7251 => x"27",
          7252 => x"88",
          7253 => x"78",
          7254 => x"5a",
          7255 => x"57",
          7256 => x"81",
          7257 => x"81",
          7258 => x"33",
          7259 => x"06",
          7260 => x"57",
          7261 => x"fe",
          7262 => x"3d",
          7263 => x"55",
          7264 => x"2e",
          7265 => x"76",
          7266 => x"38",
          7267 => x"55",
          7268 => x"33",
          7269 => x"a0",
          7270 => x"06",
          7271 => x"17",
          7272 => x"38",
          7273 => x"43",
          7274 => x"3d",
          7275 => x"ff",
          7276 => x"82",
          7277 => x"54",
          7278 => x"08",
          7279 => x"81",
          7280 => x"ff",
          7281 => x"82",
          7282 => x"54",
          7283 => x"08",
          7284 => x"80",
          7285 => x"54",
          7286 => x"80",
          7287 => x"93",
          7288 => x"2e",
          7289 => x"80",
          7290 => x"54",
          7291 => x"80",
          7292 => x"52",
          7293 => x"bd",
          7294 => x"93",
          7295 => x"82",
          7296 => x"b1",
          7297 => x"82",
          7298 => x"52",
          7299 => x"ab",
          7300 => x"54",
          7301 => x"15",
          7302 => x"78",
          7303 => x"ff",
          7304 => x"79",
          7305 => x"83",
          7306 => x"51",
          7307 => x"3f",
          7308 => x"08",
          7309 => x"74",
          7310 => x"0c",
          7311 => x"04",
          7312 => x"60",
          7313 => x"05",
          7314 => x"33",
          7315 => x"05",
          7316 => x"40",
          7317 => x"da",
          7318 => x"84",
          7319 => x"93",
          7320 => x"bd",
          7321 => x"33",
          7322 => x"b5",
          7323 => x"2e",
          7324 => x"1a",
          7325 => x"90",
          7326 => x"33",
          7327 => x"70",
          7328 => x"55",
          7329 => x"38",
          7330 => x"97",
          7331 => x"82",
          7332 => x"58",
          7333 => x"7e",
          7334 => x"70",
          7335 => x"55",
          7336 => x"56",
          7337 => x"b4",
          7338 => x"7d",
          7339 => x"70",
          7340 => x"2a",
          7341 => x"08",
          7342 => x"08",
          7343 => x"5d",
          7344 => x"77",
          7345 => x"98",
          7346 => x"26",
          7347 => x"57",
          7348 => x"59",
          7349 => x"52",
          7350 => x"ae",
          7351 => x"15",
          7352 => x"98",
          7353 => x"26",
          7354 => x"55",
          7355 => x"08",
          7356 => x"99",
          7357 => x"84",
          7358 => x"ff",
          7359 => x"93",
          7360 => x"38",
          7361 => x"75",
          7362 => x"81",
          7363 => x"93",
          7364 => x"80",
          7365 => x"2e",
          7366 => x"ff",
          7367 => x"58",
          7368 => x"7d",
          7369 => x"38",
          7370 => x"55",
          7371 => x"b4",
          7372 => x"56",
          7373 => x"09",
          7374 => x"38",
          7375 => x"53",
          7376 => x"51",
          7377 => x"3f",
          7378 => x"08",
          7379 => x"84",
          7380 => x"38",
          7381 => x"ff",
          7382 => x"5c",
          7383 => x"84",
          7384 => x"5c",
          7385 => x"12",
          7386 => x"80",
          7387 => x"78",
          7388 => x"7c",
          7389 => x"90",
          7390 => x"c0",
          7391 => x"90",
          7392 => x"15",
          7393 => x"90",
          7394 => x"54",
          7395 => x"91",
          7396 => x"31",
          7397 => x"84",
          7398 => x"07",
          7399 => x"16",
          7400 => x"73",
          7401 => x"0c",
          7402 => x"04",
          7403 => x"6b",
          7404 => x"05",
          7405 => x"33",
          7406 => x"5a",
          7407 => x"bd",
          7408 => x"80",
          7409 => x"84",
          7410 => x"f8",
          7411 => x"84",
          7412 => x"82",
          7413 => x"70",
          7414 => x"74",
          7415 => x"38",
          7416 => x"82",
          7417 => x"81",
          7418 => x"81",
          7419 => x"ff",
          7420 => x"82",
          7421 => x"81",
          7422 => x"81",
          7423 => x"83",
          7424 => x"c0",
          7425 => x"2a",
          7426 => x"51",
          7427 => x"74",
          7428 => x"99",
          7429 => x"53",
          7430 => x"51",
          7431 => x"3f",
          7432 => x"08",
          7433 => x"55",
          7434 => x"92",
          7435 => x"80",
          7436 => x"38",
          7437 => x"06",
          7438 => x"2e",
          7439 => x"48",
          7440 => x"87",
          7441 => x"79",
          7442 => x"78",
          7443 => x"26",
          7444 => x"19",
          7445 => x"74",
          7446 => x"38",
          7447 => x"e4",
          7448 => x"2a",
          7449 => x"70",
          7450 => x"59",
          7451 => x"7a",
          7452 => x"56",
          7453 => x"80",
          7454 => x"51",
          7455 => x"74",
          7456 => x"99",
          7457 => x"53",
          7458 => x"51",
          7459 => x"3f",
          7460 => x"93",
          7461 => x"ac",
          7462 => x"2a",
          7463 => x"82",
          7464 => x"43",
          7465 => x"83",
          7466 => x"66",
          7467 => x"60",
          7468 => x"90",
          7469 => x"31",
          7470 => x"80",
          7471 => x"8a",
          7472 => x"56",
          7473 => x"26",
          7474 => x"77",
          7475 => x"81",
          7476 => x"74",
          7477 => x"38",
          7478 => x"55",
          7479 => x"83",
          7480 => x"81",
          7481 => x"80",
          7482 => x"38",
          7483 => x"55",
          7484 => x"5e",
          7485 => x"89",
          7486 => x"5a",
          7487 => x"09",
          7488 => x"e1",
          7489 => x"38",
          7490 => x"57",
          7491 => x"81",
          7492 => x"5a",
          7493 => x"9d",
          7494 => x"26",
          7495 => x"81",
          7496 => x"10",
          7497 => x"22",
          7498 => x"74",
          7499 => x"38",
          7500 => x"ee",
          7501 => x"66",
          7502 => x"a0",
          7503 => x"84",
          7504 => x"84",
          7505 => x"89",
          7506 => x"a0",
          7507 => x"82",
          7508 => x"fc",
          7509 => x"56",
          7510 => x"f0",
          7511 => x"80",
          7512 => x"d3",
          7513 => x"38",
          7514 => x"57",
          7515 => x"81",
          7516 => x"5a",
          7517 => x"9d",
          7518 => x"26",
          7519 => x"81",
          7520 => x"10",
          7521 => x"22",
          7522 => x"74",
          7523 => x"38",
          7524 => x"ee",
          7525 => x"66",
          7526 => x"c0",
          7527 => x"84",
          7528 => x"05",
          7529 => x"84",
          7530 => x"26",
          7531 => x"0b",
          7532 => x"08",
          7533 => x"84",
          7534 => x"11",
          7535 => x"05",
          7536 => x"83",
          7537 => x"2a",
          7538 => x"a0",
          7539 => x"7d",
          7540 => x"69",
          7541 => x"05",
          7542 => x"72",
          7543 => x"5c",
          7544 => x"59",
          7545 => x"2e",
          7546 => x"89",
          7547 => x"60",
          7548 => x"84",
          7549 => x"5d",
          7550 => x"18",
          7551 => x"68",
          7552 => x"74",
          7553 => x"af",
          7554 => x"31",
          7555 => x"53",
          7556 => x"52",
          7557 => x"c4",
          7558 => x"84",
          7559 => x"83",
          7560 => x"06",
          7561 => x"93",
          7562 => x"ff",
          7563 => x"dd",
          7564 => x"83",
          7565 => x"2a",
          7566 => x"be",
          7567 => x"39",
          7568 => x"09",
          7569 => x"c5",
          7570 => x"f5",
          7571 => x"84",
          7572 => x"38",
          7573 => x"79",
          7574 => x"80",
          7575 => x"38",
          7576 => x"96",
          7577 => x"06",
          7578 => x"2e",
          7579 => x"5e",
          7580 => x"82",
          7581 => x"9f",
          7582 => x"38",
          7583 => x"38",
          7584 => x"81",
          7585 => x"fc",
          7586 => x"ab",
          7587 => x"7d",
          7588 => x"81",
          7589 => x"7d",
          7590 => x"78",
          7591 => x"74",
          7592 => x"8e",
          7593 => x"9c",
          7594 => x"53",
          7595 => x"51",
          7596 => x"3f",
          7597 => x"ff",
          7598 => x"51",
          7599 => x"3f",
          7600 => x"8b",
          7601 => x"a1",
          7602 => x"8d",
          7603 => x"83",
          7604 => x"52",
          7605 => x"ff",
          7606 => x"81",
          7607 => x"34",
          7608 => x"70",
          7609 => x"2a",
          7610 => x"54",
          7611 => x"1b",
          7612 => x"88",
          7613 => x"74",
          7614 => x"26",
          7615 => x"83",
          7616 => x"52",
          7617 => x"ff",
          7618 => x"8a",
          7619 => x"a0",
          7620 => x"a1",
          7621 => x"0b",
          7622 => x"bf",
          7623 => x"51",
          7624 => x"3f",
          7625 => x"9a",
          7626 => x"a0",
          7627 => x"52",
          7628 => x"ff",
          7629 => x"7d",
          7630 => x"81",
          7631 => x"38",
          7632 => x"0a",
          7633 => x"1b",
          7634 => x"ce",
          7635 => x"a4",
          7636 => x"a0",
          7637 => x"52",
          7638 => x"ff",
          7639 => x"81",
          7640 => x"51",
          7641 => x"3f",
          7642 => x"1b",
          7643 => x"8c",
          7644 => x"0b",
          7645 => x"34",
          7646 => x"c2",
          7647 => x"53",
          7648 => x"52",
          7649 => x"51",
          7650 => x"88",
          7651 => x"a7",
          7652 => x"a0",
          7653 => x"83",
          7654 => x"52",
          7655 => x"ff",
          7656 => x"ff",
          7657 => x"1c",
          7658 => x"a6",
          7659 => x"53",
          7660 => x"52",
          7661 => x"ff",
          7662 => x"82",
          7663 => x"83",
          7664 => x"52",
          7665 => x"b4",
          7666 => x"60",
          7667 => x"7e",
          7668 => x"d7",
          7669 => x"82",
          7670 => x"83",
          7671 => x"83",
          7672 => x"06",
          7673 => x"75",
          7674 => x"05",
          7675 => x"7e",
          7676 => x"b7",
          7677 => x"53",
          7678 => x"51",
          7679 => x"3f",
          7680 => x"a4",
          7681 => x"51",
          7682 => x"3f",
          7683 => x"e4",
          7684 => x"e4",
          7685 => x"9f",
          7686 => x"18",
          7687 => x"1b",
          7688 => x"f6",
          7689 => x"83",
          7690 => x"ff",
          7691 => x"82",
          7692 => x"78",
          7693 => x"c4",
          7694 => x"60",
          7695 => x"7a",
          7696 => x"ff",
          7697 => x"75",
          7698 => x"53",
          7699 => x"51",
          7700 => x"3f",
          7701 => x"52",
          7702 => x"9f",
          7703 => x"56",
          7704 => x"83",
          7705 => x"06",
          7706 => x"52",
          7707 => x"9e",
          7708 => x"52",
          7709 => x"ff",
          7710 => x"f0",
          7711 => x"1b",
          7712 => x"87",
          7713 => x"55",
          7714 => x"83",
          7715 => x"74",
          7716 => x"ff",
          7717 => x"7c",
          7718 => x"74",
          7719 => x"38",
          7720 => x"54",
          7721 => x"52",
          7722 => x"99",
          7723 => x"93",
          7724 => x"87",
          7725 => x"53",
          7726 => x"08",
          7727 => x"ff",
          7728 => x"76",
          7729 => x"31",
          7730 => x"cd",
          7731 => x"58",
          7732 => x"ff",
          7733 => x"55",
          7734 => x"83",
          7735 => x"61",
          7736 => x"26",
          7737 => x"57",
          7738 => x"53",
          7739 => x"51",
          7740 => x"3f",
          7741 => x"08",
          7742 => x"76",
          7743 => x"31",
          7744 => x"db",
          7745 => x"7d",
          7746 => x"38",
          7747 => x"83",
          7748 => x"8a",
          7749 => x"7d",
          7750 => x"38",
          7751 => x"81",
          7752 => x"80",
          7753 => x"80",
          7754 => x"7a",
          7755 => x"bc",
          7756 => x"d5",
          7757 => x"ff",
          7758 => x"83",
          7759 => x"77",
          7760 => x"0b",
          7761 => x"81",
          7762 => x"34",
          7763 => x"34",
          7764 => x"34",
          7765 => x"56",
          7766 => x"52",
          7767 => x"d7",
          7768 => x"0b",
          7769 => x"82",
          7770 => x"82",
          7771 => x"56",
          7772 => x"34",
          7773 => x"08",
          7774 => x"60",
          7775 => x"1b",
          7776 => x"96",
          7777 => x"83",
          7778 => x"ff",
          7779 => x"81",
          7780 => x"7a",
          7781 => x"ff",
          7782 => x"81",
          7783 => x"84",
          7784 => x"80",
          7785 => x"7e",
          7786 => x"e3",
          7787 => x"82",
          7788 => x"90",
          7789 => x"8e",
          7790 => x"81",
          7791 => x"82",
          7792 => x"56",
          7793 => x"84",
          7794 => x"0d",
          7795 => x"0d",
          7796 => x"59",
          7797 => x"ff",
          7798 => x"57",
          7799 => x"b4",
          7800 => x"f8",
          7801 => x"81",
          7802 => x"52",
          7803 => x"dc",
          7804 => x"2e",
          7805 => x"9c",
          7806 => x"33",
          7807 => x"2e",
          7808 => x"76",
          7809 => x"58",
          7810 => x"57",
          7811 => x"09",
          7812 => x"38",
          7813 => x"78",
          7814 => x"38",
          7815 => x"82",
          7816 => x"8d",
          7817 => x"f7",
          7818 => x"02",
          7819 => x"05",
          7820 => x"77",
          7821 => x"81",
          7822 => x"8d",
          7823 => x"e7",
          7824 => x"08",
          7825 => x"24",
          7826 => x"17",
          7827 => x"8c",
          7828 => x"77",
          7829 => x"16",
          7830 => x"25",
          7831 => x"3d",
          7832 => x"75",
          7833 => x"52",
          7834 => x"cb",
          7835 => x"76",
          7836 => x"70",
          7837 => x"2a",
          7838 => x"51",
          7839 => x"84",
          7840 => x"19",
          7841 => x"8b",
          7842 => x"f9",
          7843 => x"84",
          7844 => x"56",
          7845 => x"a7",
          7846 => x"fc",
          7847 => x"53",
          7848 => x"75",
          7849 => x"a1",
          7850 => x"84",
          7851 => x"84",
          7852 => x"2e",
          7853 => x"87",
          7854 => x"08",
          7855 => x"ff",
          7856 => x"93",
          7857 => x"3d",
          7858 => x"3d",
          7859 => x"80",
          7860 => x"52",
          7861 => x"9a",
          7862 => x"74",
          7863 => x"0d",
          7864 => x"0d",
          7865 => x"05",
          7866 => x"86",
          7867 => x"54",
          7868 => x"73",
          7869 => x"fe",
          7870 => x"51",
          7871 => x"98",
          7872 => x"f8",
          7873 => x"70",
          7874 => x"56",
          7875 => x"2e",
          7876 => x"8c",
          7877 => x"79",
          7878 => x"33",
          7879 => x"39",
          7880 => x"73",
          7881 => x"81",
          7882 => x"81",
          7883 => x"39",
          7884 => x"90",
          7885 => x"f4",
          7886 => x"52",
          7887 => x"af",
          7888 => x"84",
          7889 => x"84",
          7890 => x"53",
          7891 => x"58",
          7892 => x"3f",
          7893 => x"08",
          7894 => x"16",
          7895 => x"81",
          7896 => x"38",
          7897 => x"81",
          7898 => x"54",
          7899 => x"c2",
          7900 => x"73",
          7901 => x"0c",
          7902 => x"04",
          7903 => x"73",
          7904 => x"26",
          7905 => x"71",
          7906 => x"f6",
          7907 => x"71",
          7908 => x"82",
          7909 => x"80",
          7910 => x"d8",
          7911 => x"39",
          7912 => x"51",
          7913 => x"82",
          7914 => x"80",
          7915 => x"83",
          7916 => x"e4",
          7917 => x"a0",
          7918 => x"39",
          7919 => x"51",
          7920 => x"82",
          7921 => x"80",
          7922 => x"83",
          7923 => x"c8",
          7924 => x"f4",
          7925 => x"39",
          7926 => x"51",
          7927 => x"84",
          7928 => x"39",
          7929 => x"51",
          7930 => x"84",
          7931 => x"39",
          7932 => x"51",
          7933 => x"85",
          7934 => x"39",
          7935 => x"51",
          7936 => x"85",
          7937 => x"39",
          7938 => x"51",
          7939 => x"85",
          7940 => x"39",
          7941 => x"51",
          7942 => x"3f",
          7943 => x"04",
          7944 => x"77",
          7945 => x"74",
          7946 => x"8a",
          7947 => x"75",
          7948 => x"51",
          7949 => x"e8",
          7950 => x"fe",
          7951 => x"82",
          7952 => x"52",
          7953 => x"d2",
          7954 => x"93",
          7955 => x"79",
          7956 => x"82",
          7957 => x"fe",
          7958 => x"87",
          7959 => x"ec",
          7960 => x"02",
          7961 => x"e3",
          7962 => x"57",
          7963 => x"30",
          7964 => x"73",
          7965 => x"59",
          7966 => x"77",
          7967 => x"83",
          7968 => x"74",
          7969 => x"81",
          7970 => x"55",
          7971 => x"81",
          7972 => x"53",
          7973 => x"3d",
          7974 => x"ff",
          7975 => x"82",
          7976 => x"57",
          7977 => x"08",
          7978 => x"93",
          7979 => x"c0",
          7980 => x"82",
          7981 => x"59",
          7982 => x"05",
          7983 => x"53",
          7984 => x"51",
          7985 => x"82",
          7986 => x"57",
          7987 => x"08",
          7988 => x"55",
          7989 => x"89",
          7990 => x"75",
          7991 => x"d8",
          7992 => x"d8",
          7993 => x"f0",
          7994 => x"70",
          7995 => x"25",
          7996 => x"9f",
          7997 => x"51",
          7998 => x"74",
          7999 => x"38",
          8000 => x"53",
          8001 => x"88",
          8002 => x"51",
          8003 => x"76",
          8004 => x"93",
          8005 => x"3d",
          8006 => x"3d",
          8007 => x"84",
          8008 => x"33",
          8009 => x"57",
          8010 => x"52",
          8011 => x"af",
          8012 => x"84",
          8013 => x"75",
          8014 => x"38",
          8015 => x"98",
          8016 => x"60",
          8017 => x"82",
          8018 => x"7e",
          8019 => x"77",
          8020 => x"84",
          8021 => x"39",
          8022 => x"82",
          8023 => x"89",
          8024 => x"f3",
          8025 => x"61",
          8026 => x"05",
          8027 => x"33",
          8028 => x"68",
          8029 => x"5c",
          8030 => x"7a",
          8031 => x"c0",
          8032 => x"a9",
          8033 => x"c8",
          8034 => x"bd",
          8035 => x"74",
          8036 => x"fc",
          8037 => x"2e",
          8038 => x"a0",
          8039 => x"80",
          8040 => x"18",
          8041 => x"27",
          8042 => x"22",
          8043 => x"cc",
          8044 => x"f9",
          8045 => x"82",
          8046 => x"fe",
          8047 => x"82",
          8048 => x"c3",
          8049 => x"53",
          8050 => x"8e",
          8051 => x"52",
          8052 => x"51",
          8053 => x"3f",
          8054 => x"86",
          8055 => x"ee",
          8056 => x"15",
          8057 => x"74",
          8058 => x"7a",
          8059 => x"72",
          8060 => x"86",
          8061 => x"f4",
          8062 => x"39",
          8063 => x"51",
          8064 => x"3f",
          8065 => x"a0",
          8066 => x"e0",
          8067 => x"39",
          8068 => x"51",
          8069 => x"3f",
          8070 => x"79",
          8071 => x"74",
          8072 => x"55",
          8073 => x"72",
          8074 => x"38",
          8075 => x"53",
          8076 => x"83",
          8077 => x"75",
          8078 => x"81",
          8079 => x"53",
          8080 => x"8b",
          8081 => x"fe",
          8082 => x"73",
          8083 => x"a0",
          8084 => x"98",
          8085 => x"55",
          8086 => x"86",
          8087 => x"ed",
          8088 => x"18",
          8089 => x"58",
          8090 => x"3f",
          8091 => x"08",
          8092 => x"98",
          8093 => x"76",
          8094 => x"81",
          8095 => x"fe",
          8096 => x"82",
          8097 => x"98",
          8098 => x"2c",
          8099 => x"70",
          8100 => x"32",
          8101 => x"72",
          8102 => x"07",
          8103 => x"58",
          8104 => x"57",
          8105 => x"d7",
          8106 => x"2e",
          8107 => x"85",
          8108 => x"8c",
          8109 => x"53",
          8110 => x"fd",
          8111 => x"53",
          8112 => x"84",
          8113 => x"0d",
          8114 => x"0d",
          8115 => x"33",
          8116 => x"53",
          8117 => x"52",
          8118 => x"d1",
          8119 => x"b4",
          8120 => x"e6",
          8121 => x"87",
          8122 => x"87",
          8123 => x"8e",
          8124 => x"82",
          8125 => x"fe",
          8126 => x"74",
          8127 => x"38",
          8128 => x"3f",
          8129 => x"04",
          8130 => x"87",
          8131 => x"08",
          8132 => x"b1",
          8133 => x"fe",
          8134 => x"82",
          8135 => x"fe",
          8136 => x"80",
          8137 => x"eb",
          8138 => x"2a",
          8139 => x"51",
          8140 => x"2e",
          8141 => x"51",
          8142 => x"3f",
          8143 => x"51",
          8144 => x"3f",
          8145 => x"d8",
          8146 => x"82",
          8147 => x"06",
          8148 => x"80",
          8149 => x"81",
          8150 => x"b7",
          8151 => x"e8",
          8152 => x"af",
          8153 => x"fe",
          8154 => x"72",
          8155 => x"81",
          8156 => x"71",
          8157 => x"38",
          8158 => x"d8",
          8159 => x"87",
          8160 => x"da",
          8161 => x"51",
          8162 => x"3f",
          8163 => x"70",
          8164 => x"52",
          8165 => x"95",
          8166 => x"fe",
          8167 => x"82",
          8168 => x"fe",
          8169 => x"80",
          8170 => x"e7",
          8171 => x"2a",
          8172 => x"51",
          8173 => x"2e",
          8174 => x"51",
          8175 => x"3f",
          8176 => x"51",
          8177 => x"3f",
          8178 => x"d7",
          8179 => x"86",
          8180 => x"06",
          8181 => x"80",
          8182 => x"81",
          8183 => x"b3",
          8184 => x"b4",
          8185 => x"ab",
          8186 => x"fe",
          8187 => x"72",
          8188 => x"81",
          8189 => x"71",
          8190 => x"38",
          8191 => x"d7",
          8192 => x"88",
          8193 => x"d9",
          8194 => x"51",
          8195 => x"3f",
          8196 => x"70",
          8197 => x"52",
          8198 => x"95",
          8199 => x"fe",
          8200 => x"82",
          8201 => x"fe",
          8202 => x"80",
          8203 => x"e3",
          8204 => x"99",
          8205 => x"0d",
          8206 => x"0d",
          8207 => x"05",
          8208 => x"70",
          8209 => x"80",
          8210 => x"fe",
          8211 => x"82",
          8212 => x"54",
          8213 => x"81",
          8214 => x"9c",
          8215 => x"9c",
          8216 => x"83",
          8217 => x"84",
          8218 => x"82",
          8219 => x"07",
          8220 => x"71",
          8221 => x"54",
          8222 => x"f0",
          8223 => x"f0",
          8224 => x"81",
          8225 => x"06",
          8226 => x"aa",
          8227 => x"52",
          8228 => x"b9",
          8229 => x"84",
          8230 => x"8c",
          8231 => x"84",
          8232 => x"e9",
          8233 => x"39",
          8234 => x"51",
          8235 => x"82",
          8236 => x"f0",
          8237 => x"f0",
          8238 => x"82",
          8239 => x"06",
          8240 => x"52",
          8241 => x"fa",
          8242 => x"0b",
          8243 => x"0c",
          8244 => x"04",
          8245 => x"80",
          8246 => x"aa",
          8247 => x"5d",
          8248 => x"51",
          8249 => x"3f",
          8250 => x"08",
          8251 => x"59",
          8252 => x"09",
          8253 => x"38",
          8254 => x"52",
          8255 => x"52",
          8256 => x"bf",
          8257 => x"78",
          8258 => x"c8",
          8259 => x"f6",
          8260 => x"84",
          8261 => x"88",
          8262 => x"b0",
          8263 => x"39",
          8264 => x"5d",
          8265 => x"51",
          8266 => x"3f",
          8267 => x"46",
          8268 => x"52",
          8269 => x"81",
          8270 => x"ff",
          8271 => x"f3",
          8272 => x"93",
          8273 => x"2b",
          8274 => x"51",
          8275 => x"c1",
          8276 => x"38",
          8277 => x"24",
          8278 => x"78",
          8279 => x"c0",
          8280 => x"24",
          8281 => x"82",
          8282 => x"38",
          8283 => x"8a",
          8284 => x"2e",
          8285 => x"8f",
          8286 => x"84",
          8287 => x"38",
          8288 => x"82",
          8289 => x"96",
          8290 => x"2e",
          8291 => x"78",
          8292 => x"38",
          8293 => x"83",
          8294 => x"bc",
          8295 => x"38",
          8296 => x"78",
          8297 => x"d7",
          8298 => x"c0",
          8299 => x"38",
          8300 => x"78",
          8301 => x"8d",
          8302 => x"80",
          8303 => x"38",
          8304 => x"2e",
          8305 => x"78",
          8306 => x"92",
          8307 => x"c2",
          8308 => x"38",
          8309 => x"2e",
          8310 => x"8e",
          8311 => x"80",
          8312 => x"e9",
          8313 => x"d4",
          8314 => x"38",
          8315 => x"78",
          8316 => x"8e",
          8317 => x"81",
          8318 => x"38",
          8319 => x"2e",
          8320 => x"78",
          8321 => x"8d",
          8322 => x"92",
          8323 => x"83",
          8324 => x"38",
          8325 => x"2e",
          8326 => x"8e",
          8327 => x"3d",
          8328 => x"53",
          8329 => x"51",
          8330 => x"3f",
          8331 => x"08",
          8332 => x"89",
          8333 => x"e5",
          8334 => x"fe",
          8335 => x"ff",
          8336 => x"fe",
          8337 => x"82",
          8338 => x"80",
          8339 => x"81",
          8340 => x"38",
          8341 => x"80",
          8342 => x"52",
          8343 => x"05",
          8344 => x"83",
          8345 => x"93",
          8346 => x"ff",
          8347 => x"8e",
          8348 => x"fc",
          8349 => x"d1",
          8350 => x"fd",
          8351 => x"8a",
          8352 => x"b9",
          8353 => x"ff",
          8354 => x"ff",
          8355 => x"fe",
          8356 => x"82",
          8357 => x"80",
          8358 => x"38",
          8359 => x"52",
          8360 => x"05",
          8361 => x"87",
          8362 => x"93",
          8363 => x"82",
          8364 => x"8c",
          8365 => x"3d",
          8366 => x"53",
          8367 => x"51",
          8368 => x"3f",
          8369 => x"08",
          8370 => x"38",
          8371 => x"fc",
          8372 => x"3d",
          8373 => x"53",
          8374 => x"51",
          8375 => x"3f",
          8376 => x"08",
          8377 => x"93",
          8378 => x"63",
          8379 => x"ac",
          8380 => x"fe",
          8381 => x"02",
          8382 => x"33",
          8383 => x"63",
          8384 => x"82",
          8385 => x"51",
          8386 => x"3f",
          8387 => x"08",
          8388 => x"82",
          8389 => x"fe",
          8390 => x"81",
          8391 => x"39",
          8392 => x"84",
          8393 => x"cd",
          8394 => x"93",
          8395 => x"3d",
          8396 => x"52",
          8397 => x"ee",
          8398 => x"82",
          8399 => x"52",
          8400 => x"9b",
          8401 => x"39",
          8402 => x"84",
          8403 => x"cc",
          8404 => x"93",
          8405 => x"3d",
          8406 => x"52",
          8407 => x"c6",
          8408 => x"84",
          8409 => x"ff",
          8410 => x"5a",
          8411 => x"3f",
          8412 => x"08",
          8413 => x"84",
          8414 => x"fe",
          8415 => x"82",
          8416 => x"82",
          8417 => x"80",
          8418 => x"82",
          8419 => x"81",
          8420 => x"78",
          8421 => x"7a",
          8422 => x"3f",
          8423 => x"08",
          8424 => x"80",
          8425 => x"84",
          8426 => x"d0",
          8427 => x"39",
          8428 => x"80",
          8429 => x"84",
          8430 => x"ea",
          8431 => x"93",
          8432 => x"2e",
          8433 => x"b4",
          8434 => x"11",
          8435 => x"05",
          8436 => x"ce",
          8437 => x"84",
          8438 => x"fa",
          8439 => x"3d",
          8440 => x"53",
          8441 => x"51",
          8442 => x"3f",
          8443 => x"08",
          8444 => x"93",
          8445 => x"82",
          8446 => x"fe",
          8447 => x"63",
          8448 => x"79",
          8449 => x"f2",
          8450 => x"78",
          8451 => x"05",
          8452 => x"7a",
          8453 => x"81",
          8454 => x"3d",
          8455 => x"53",
          8456 => x"51",
          8457 => x"3f",
          8458 => x"08",
          8459 => x"f4",
          8460 => x"fe",
          8461 => x"ff",
          8462 => x"fe",
          8463 => x"82",
          8464 => x"80",
          8465 => x"38",
          8466 => x"f8",
          8467 => x"84",
          8468 => x"e9",
          8469 => x"93",
          8470 => x"2e",
          8471 => x"82",
          8472 => x"fe",
          8473 => x"63",
          8474 => x"27",
          8475 => x"61",
          8476 => x"81",
          8477 => x"79",
          8478 => x"05",
          8479 => x"b4",
          8480 => x"11",
          8481 => x"05",
          8482 => x"96",
          8483 => x"84",
          8484 => x"f9",
          8485 => x"3d",
          8486 => x"53",
          8487 => x"51",
          8488 => x"3f",
          8489 => x"08",
          8490 => x"f8",
          8491 => x"fe",
          8492 => x"ff",
          8493 => x"fe",
          8494 => x"82",
          8495 => x"80",
          8496 => x"38",
          8497 => x"51",
          8498 => x"3f",
          8499 => x"63",
          8500 => x"61",
          8501 => x"33",
          8502 => x"78",
          8503 => x"38",
          8504 => x"54",
          8505 => x"79",
          8506 => x"dc",
          8507 => x"bd",
          8508 => x"62",
          8509 => x"5a",
          8510 => x"89",
          8511 => x"bd",
          8512 => x"ff",
          8513 => x"ff",
          8514 => x"fe",
          8515 => x"82",
          8516 => x"80",
          8517 => x"8e",
          8518 => x"78",
          8519 => x"38",
          8520 => x"08",
          8521 => x"39",
          8522 => x"33",
          8523 => x"2e",
          8524 => x"8e",
          8525 => x"bc",
          8526 => x"ca",
          8527 => x"80",
          8528 => x"82",
          8529 => x"44",
          8530 => x"8e",
          8531 => x"78",
          8532 => x"38",
          8533 => x"08",
          8534 => x"82",
          8535 => x"59",
          8536 => x"88",
          8537 => x"a0",
          8538 => x"39",
          8539 => x"08",
          8540 => x"44",
          8541 => x"fc",
          8542 => x"84",
          8543 => x"e7",
          8544 => x"93",
          8545 => x"de",
          8546 => x"c8",
          8547 => x"80",
          8548 => x"82",
          8549 => x"43",
          8550 => x"82",
          8551 => x"59",
          8552 => x"88",
          8553 => x"8c",
          8554 => x"39",
          8555 => x"33",
          8556 => x"2e",
          8557 => x"8e",
          8558 => x"aa",
          8559 => x"cb",
          8560 => x"80",
          8561 => x"82",
          8562 => x"43",
          8563 => x"8e",
          8564 => x"78",
          8565 => x"38",
          8566 => x"08",
          8567 => x"82",
          8568 => x"88",
          8569 => x"3d",
          8570 => x"53",
          8571 => x"51",
          8572 => x"3f",
          8573 => x"08",
          8574 => x"38",
          8575 => x"5c",
          8576 => x"83",
          8577 => x"7a",
          8578 => x"30",
          8579 => x"9f",
          8580 => x"06",
          8581 => x"5a",
          8582 => x"88",
          8583 => x"2e",
          8584 => x"42",
          8585 => x"51",
          8586 => x"3f",
          8587 => x"54",
          8588 => x"52",
          8589 => x"ab",
          8590 => x"88",
          8591 => x"89",
          8592 => x"39",
          8593 => x"80",
          8594 => x"84",
          8595 => x"e5",
          8596 => x"93",
          8597 => x"2e",
          8598 => x"b4",
          8599 => x"11",
          8600 => x"05",
          8601 => x"ba",
          8602 => x"84",
          8603 => x"a5",
          8604 => x"02",
          8605 => x"33",
          8606 => x"81",
          8607 => x"3d",
          8608 => x"53",
          8609 => x"51",
          8610 => x"3f",
          8611 => x"08",
          8612 => x"90",
          8613 => x"33",
          8614 => x"8b",
          8615 => x"e3",
          8616 => x"f8",
          8617 => x"fe",
          8618 => x"79",
          8619 => x"59",
          8620 => x"f4",
          8621 => x"79",
          8622 => x"b4",
          8623 => x"11",
          8624 => x"05",
          8625 => x"da",
          8626 => x"84",
          8627 => x"91",
          8628 => x"02",
          8629 => x"33",
          8630 => x"81",
          8631 => x"b5",
          8632 => x"a0",
          8633 => x"e1",
          8634 => x"39",
          8635 => x"f4",
          8636 => x"84",
          8637 => x"e6",
          8638 => x"93",
          8639 => x"2e",
          8640 => x"b4",
          8641 => x"11",
          8642 => x"05",
          8643 => x"84",
          8644 => x"84",
          8645 => x"a6",
          8646 => x"02",
          8647 => x"79",
          8648 => x"5b",
          8649 => x"b4",
          8650 => x"11",
          8651 => x"05",
          8652 => x"e0",
          8653 => x"84",
          8654 => x"f3",
          8655 => x"70",
          8656 => x"82",
          8657 => x"fe",
          8658 => x"80",
          8659 => x"51",
          8660 => x"3f",
          8661 => x"33",
          8662 => x"2e",
          8663 => x"78",
          8664 => x"38",
          8665 => x"41",
          8666 => x"3d",
          8667 => x"53",
          8668 => x"51",
          8669 => x"3f",
          8670 => x"08",
          8671 => x"38",
          8672 => x"be",
          8673 => x"70",
          8674 => x"23",
          8675 => x"ae",
          8676 => x"a0",
          8677 => x"b1",
          8678 => x"39",
          8679 => x"f4",
          8680 => x"84",
          8681 => x"e4",
          8682 => x"93",
          8683 => x"2e",
          8684 => x"b4",
          8685 => x"11",
          8686 => x"05",
          8687 => x"d4",
          8688 => x"84",
          8689 => x"a1",
          8690 => x"71",
          8691 => x"84",
          8692 => x"3d",
          8693 => x"53",
          8694 => x"51",
          8695 => x"3f",
          8696 => x"08",
          8697 => x"bc",
          8698 => x"08",
          8699 => x"8b",
          8700 => x"e0",
          8701 => x"f8",
          8702 => x"fe",
          8703 => x"79",
          8704 => x"59",
          8705 => x"f2",
          8706 => x"79",
          8707 => x"b4",
          8708 => x"11",
          8709 => x"05",
          8710 => x"f8",
          8711 => x"84",
          8712 => x"8d",
          8713 => x"71",
          8714 => x"84",
          8715 => x"b9",
          8716 => x"a0",
          8717 => x"91",
          8718 => x"39",
          8719 => x"51",
          8720 => x"3f",
          8721 => x"d4",
          8722 => x"d8",
          8723 => x"d8",
          8724 => x"f5",
          8725 => x"fe",
          8726 => x"f1",
          8727 => x"8b",
          8728 => x"d9",
          8729 => x"80",
          8730 => x"c0",
          8731 => x"84",
          8732 => x"87",
          8733 => x"0c",
          8734 => x"82",
          8735 => x"fe",
          8736 => x"8c",
          8737 => x"87",
          8738 => x"0c",
          8739 => x"0b",
          8740 => x"94",
          8741 => x"39",
          8742 => x"80",
          8743 => x"84",
          8744 => x"e0",
          8745 => x"93",
          8746 => x"2e",
          8747 => x"63",
          8748 => x"98",
          8749 => x"f5",
          8750 => x"78",
          8751 => x"ff",
          8752 => x"ff",
          8753 => x"fe",
          8754 => x"82",
          8755 => x"80",
          8756 => x"38",
          8757 => x"8c",
          8758 => x"de",
          8759 => x"59",
          8760 => x"93",
          8761 => x"2e",
          8762 => x"82",
          8763 => x"52",
          8764 => x"51",
          8765 => x"3f",
          8766 => x"82",
          8767 => x"fe",
          8768 => x"fe",
          8769 => x"f0",
          8770 => x"8d",
          8771 => x"d8",
          8772 => x"59",
          8773 => x"fe",
          8774 => x"f0",
          8775 => x"45",
          8776 => x"78",
          8777 => x"fc",
          8778 => x"06",
          8779 => x"2e",
          8780 => x"b4",
          8781 => x"05",
          8782 => x"88",
          8783 => x"84",
          8784 => x"5c",
          8785 => x"b2",
          8786 => x"24",
          8787 => x"81",
          8788 => x"80",
          8789 => x"83",
          8790 => x"80",
          8791 => x"8d",
          8792 => x"55",
          8793 => x"54",
          8794 => x"8d",
          8795 => x"3d",
          8796 => x"51",
          8797 => x"3f",
          8798 => x"8d",
          8799 => x"3d",
          8800 => x"51",
          8801 => x"3f",
          8802 => x"55",
          8803 => x"54",
          8804 => x"8d",
          8805 => x"3d",
          8806 => x"51",
          8807 => x"3f",
          8808 => x"54",
          8809 => x"8d",
          8810 => x"3d",
          8811 => x"51",
          8812 => x"3f",
          8813 => x"58",
          8814 => x"57",
          8815 => x"55",
          8816 => x"80",
          8817 => x"80",
          8818 => x"3d",
          8819 => x"51",
          8820 => x"82",
          8821 => x"82",
          8822 => x"09",
          8823 => x"72",
          8824 => x"51",
          8825 => x"80",
          8826 => x"26",
          8827 => x"5a",
          8828 => x"59",
          8829 => x"8d",
          8830 => x"70",
          8831 => x"5d",
          8832 => x"c0",
          8833 => x"32",
          8834 => x"07",
          8835 => x"38",
          8836 => x"09",
          8837 => x"8c",
          8838 => x"c8",
          8839 => x"8d",
          8840 => x"39",
          8841 => x"80",
          8842 => x"cc",
          8843 => x"94",
          8844 => x"54",
          8845 => x"80",
          8846 => x"fe",
          8847 => x"82",
          8848 => x"90",
          8849 => x"55",
          8850 => x"80",
          8851 => x"fe",
          8852 => x"72",
          8853 => x"08",
          8854 => x"87",
          8855 => x"70",
          8856 => x"87",
          8857 => x"72",
          8858 => x"f0",
          8859 => x"84",
          8860 => x"75",
          8861 => x"87",
          8862 => x"73",
          8863 => x"dc",
          8864 => x"93",
          8865 => x"75",
          8866 => x"83",
          8867 => x"94",
          8868 => x"80",
          8869 => x"c0",
          8870 => x"b7",
          8871 => x"93",
          8872 => x"ad",
          8873 => x"9c",
          8874 => x"ab",
          8875 => x"95",
          8876 => x"d8",
          8877 => x"91",
          8878 => x"e4",
          8879 => x"89",
          8880 => x"87",
          8881 => x"b7",
          8882 => x"e7",
          8883 => x"84",
          8884 => x"00",
          8885 => x"22",
          8886 => x"22",
          8887 => x"22",
          8888 => x"22",
          8889 => x"22",
          8890 => x"30",
          8891 => x"30",
          8892 => x"31",
          8893 => x"31",
          8894 => x"31",
          8895 => x"32",
          8896 => x"2e",
          8897 => x"2e",
          8898 => x"32",
          8899 => x"33",
          8900 => x"33",
          8901 => x"33",
          8902 => x"6c",
          8903 => x"6b",
          8904 => x"6b",
          8905 => x"6b",
          8906 => x"6b",
          8907 => x"6b",
          8908 => x"6b",
          8909 => x"6b",
          8910 => x"6b",
          8911 => x"6b",
          8912 => x"6b",
          8913 => x"6b",
          8914 => x"6b",
          8915 => x"6b",
          8916 => x"6b",
          8917 => x"6b",
          8918 => x"6b",
          8919 => x"6b",
          8920 => x"6c",
          8921 => x"6c",
          8922 => x"2f",
          8923 => x"25",
          8924 => x"64",
          8925 => x"3a",
          8926 => x"25",
          8927 => x"0a",
          8928 => x"43",
          8929 => x"6e",
          8930 => x"75",
          8931 => x"69",
          8932 => x"00",
          8933 => x"66",
          8934 => x"20",
          8935 => x"20",
          8936 => x"66",
          8937 => x"00",
          8938 => x"44",
          8939 => x"63",
          8940 => x"69",
          8941 => x"65",
          8942 => x"74",
          8943 => x"0a",
          8944 => x"20",
          8945 => x"20",
          8946 => x"41",
          8947 => x"28",
          8948 => x"58",
          8949 => x"38",
          8950 => x"0a",
          8951 => x"20",
          8952 => x"52",
          8953 => x"20",
          8954 => x"28",
          8955 => x"58",
          8956 => x"38",
          8957 => x"0a",
          8958 => x"20",
          8959 => x"53",
          8960 => x"52",
          8961 => x"28",
          8962 => x"58",
          8963 => x"38",
          8964 => x"0a",
          8965 => x"20",
          8966 => x"41",
          8967 => x"20",
          8968 => x"28",
          8969 => x"58",
          8970 => x"38",
          8971 => x"0a",
          8972 => x"20",
          8973 => x"4d",
          8974 => x"20",
          8975 => x"28",
          8976 => x"58",
          8977 => x"38",
          8978 => x"0a",
          8979 => x"20",
          8980 => x"20",
          8981 => x"44",
          8982 => x"28",
          8983 => x"69",
          8984 => x"20",
          8985 => x"32",
          8986 => x"0a",
          8987 => x"20",
          8988 => x"4d",
          8989 => x"20",
          8990 => x"28",
          8991 => x"65",
          8992 => x"20",
          8993 => x"32",
          8994 => x"0a",
          8995 => x"20",
          8996 => x"54",
          8997 => x"54",
          8998 => x"28",
          8999 => x"6e",
          9000 => x"73",
          9001 => x"32",
          9002 => x"0a",
          9003 => x"20",
          9004 => x"53",
          9005 => x"4e",
          9006 => x"55",
          9007 => x"00",
          9008 => x"20",
          9009 => x"20",
          9010 => x"0a",
          9011 => x"20",
          9012 => x"43",
          9013 => x"00",
          9014 => x"20",
          9015 => x"32",
          9016 => x"00",
          9017 => x"20",
          9018 => x"49",
          9019 => x"00",
          9020 => x"64",
          9021 => x"73",
          9022 => x"0a",
          9023 => x"20",
          9024 => x"55",
          9025 => x"73",
          9026 => x"56",
          9027 => x"6f",
          9028 => x"64",
          9029 => x"73",
          9030 => x"20",
          9031 => x"58",
          9032 => x"00",
          9033 => x"20",
          9034 => x"55",
          9035 => x"6d",
          9036 => x"20",
          9037 => x"72",
          9038 => x"64",
          9039 => x"73",
          9040 => x"20",
          9041 => x"58",
          9042 => x"00",
          9043 => x"20",
          9044 => x"61",
          9045 => x"53",
          9046 => x"74",
          9047 => x"64",
          9048 => x"73",
          9049 => x"20",
          9050 => x"20",
          9051 => x"58",
          9052 => x"00",
          9053 => x"73",
          9054 => x"00",
          9055 => x"20",
          9056 => x"55",
          9057 => x"20",
          9058 => x"20",
          9059 => x"20",
          9060 => x"20",
          9061 => x"20",
          9062 => x"20",
          9063 => x"58",
          9064 => x"00",
          9065 => x"20",
          9066 => x"73",
          9067 => x"20",
          9068 => x"63",
          9069 => x"72",
          9070 => x"20",
          9071 => x"20",
          9072 => x"20",
          9073 => x"25",
          9074 => x"4d",
          9075 => x"00",
          9076 => x"20",
          9077 => x"52",
          9078 => x"43",
          9079 => x"6b",
          9080 => x"65",
          9081 => x"20",
          9082 => x"20",
          9083 => x"20",
          9084 => x"25",
          9085 => x"4d",
          9086 => x"00",
          9087 => x"20",
          9088 => x"73",
          9089 => x"6e",
          9090 => x"44",
          9091 => x"20",
          9092 => x"63",
          9093 => x"72",
          9094 => x"20",
          9095 => x"25",
          9096 => x"4d",
          9097 => x"00",
          9098 => x"61",
          9099 => x"00",
          9100 => x"64",
          9101 => x"00",
          9102 => x"65",
          9103 => x"00",
          9104 => x"4f",
          9105 => x"4f",
          9106 => x"00",
          9107 => x"6b",
          9108 => x"6e",
          9109 => x"73",
          9110 => x"79",
          9111 => x"74",
          9112 => x"73",
          9113 => x"79",
          9114 => x"73",
          9115 => x"00",
          9116 => x"00",
          9117 => x"34",
          9118 => x"25",
          9119 => x"00",
          9120 => x"69",
          9121 => x"20",
          9122 => x"72",
          9123 => x"74",
          9124 => x"65",
          9125 => x"73",
          9126 => x"79",
          9127 => x"6c",
          9128 => x"6f",
          9129 => x"46",
          9130 => x"00",
          9131 => x"6e",
          9132 => x"20",
          9133 => x"6e",
          9134 => x"65",
          9135 => x"20",
          9136 => x"74",
          9137 => x"20",
          9138 => x"65",
          9139 => x"69",
          9140 => x"6c",
          9141 => x"2e",
          9142 => x"00",
          9143 => x"7f",
          9144 => x"00",
          9145 => x"00",
          9146 => x"7f",
          9147 => x"00",
          9148 => x"00",
          9149 => x"7f",
          9150 => x"00",
          9151 => x"00",
          9152 => x"7f",
          9153 => x"00",
          9154 => x"00",
          9155 => x"7f",
          9156 => x"00",
          9157 => x"00",
          9158 => x"7f",
          9159 => x"00",
          9160 => x"00",
          9161 => x"7f",
          9162 => x"00",
          9163 => x"00",
          9164 => x"7f",
          9165 => x"00",
          9166 => x"00",
          9167 => x"7f",
          9168 => x"00",
          9169 => x"00",
          9170 => x"7f",
          9171 => x"00",
          9172 => x"00",
          9173 => x"7f",
          9174 => x"00",
          9175 => x"00",
          9176 => x"44",
          9177 => x"43",
          9178 => x"42",
          9179 => x"41",
          9180 => x"36",
          9181 => x"35",
          9182 => x"34",
          9183 => x"33",
          9184 => x"31",
          9185 => x"00",
          9186 => x"00",
          9187 => x"00",
          9188 => x"2b",
          9189 => x"3c",
          9190 => x"5b",
          9191 => x"00",
          9192 => x"54",
          9193 => x"54",
          9194 => x"00",
          9195 => x"90",
          9196 => x"4f",
          9197 => x"30",
          9198 => x"20",
          9199 => x"45",
          9200 => x"20",
          9201 => x"33",
          9202 => x"20",
          9203 => x"20",
          9204 => x"45",
          9205 => x"20",
          9206 => x"20",
          9207 => x"20",
          9208 => x"7f",
          9209 => x"00",
          9210 => x"00",
          9211 => x"00",
          9212 => x"45",
          9213 => x"8f",
          9214 => x"45",
          9215 => x"8e",
          9216 => x"92",
          9217 => x"55",
          9218 => x"9a",
          9219 => x"9e",
          9220 => x"4f",
          9221 => x"a6",
          9222 => x"aa",
          9223 => x"ae",
          9224 => x"b2",
          9225 => x"b6",
          9226 => x"ba",
          9227 => x"be",
          9228 => x"c2",
          9229 => x"c6",
          9230 => x"ca",
          9231 => x"ce",
          9232 => x"d2",
          9233 => x"d6",
          9234 => x"da",
          9235 => x"de",
          9236 => x"e2",
          9237 => x"e6",
          9238 => x"ea",
          9239 => x"ee",
          9240 => x"f2",
          9241 => x"f6",
          9242 => x"fa",
          9243 => x"fe",
          9244 => x"2c",
          9245 => x"5d",
          9246 => x"2a",
          9247 => x"3f",
          9248 => x"00",
          9249 => x"00",
          9250 => x"00",
          9251 => x"02",
          9252 => x"00",
          9253 => x"00",
          9254 => x"00",
          9255 => x"00",
          9256 => x"00",
          9257 => x"6e",
          9258 => x"00",
          9259 => x"6f",
          9260 => x"00",
          9261 => x"6e",
          9262 => x"00",
          9263 => x"6f",
          9264 => x"00",
          9265 => x"78",
          9266 => x"00",
          9267 => x"6c",
          9268 => x"00",
          9269 => x"6f",
          9270 => x"00",
          9271 => x"69",
          9272 => x"00",
          9273 => x"75",
          9274 => x"00",
          9275 => x"62",
          9276 => x"68",
          9277 => x"77",
          9278 => x"64",
          9279 => x"65",
          9280 => x"64",
          9281 => x"65",
          9282 => x"6c",
          9283 => x"00",
          9284 => x"70",
          9285 => x"73",
          9286 => x"74",
          9287 => x"73",
          9288 => x"00",
          9289 => x"66",
          9290 => x"00",
          9291 => x"73",
          9292 => x"00",
          9293 => x"61",
          9294 => x"00",
          9295 => x"61",
          9296 => x"00",
          9297 => x"6c",
          9298 => x"00",
          9299 => x"73",
          9300 => x"72",
          9301 => x"0a",
          9302 => x"74",
          9303 => x"61",
          9304 => x"72",
          9305 => x"2e",
          9306 => x"00",
          9307 => x"73",
          9308 => x"6f",
          9309 => x"65",
          9310 => x"2e",
          9311 => x"00",
          9312 => x"20",
          9313 => x"65",
          9314 => x"75",
          9315 => x"0a",
          9316 => x"20",
          9317 => x"68",
          9318 => x"75",
          9319 => x"0a",
          9320 => x"76",
          9321 => x"64",
          9322 => x"6c",
          9323 => x"6d",
          9324 => x"00",
          9325 => x"63",
          9326 => x"20",
          9327 => x"69",
          9328 => x"0a",
          9329 => x"6c",
          9330 => x"6c",
          9331 => x"64",
          9332 => x"78",
          9333 => x"73",
          9334 => x"00",
          9335 => x"6c",
          9336 => x"61",
          9337 => x"65",
          9338 => x"76",
          9339 => x"64",
          9340 => x"00",
          9341 => x"20",
          9342 => x"77",
          9343 => x"65",
          9344 => x"6f",
          9345 => x"74",
          9346 => x"0a",
          9347 => x"69",
          9348 => x"6e",
          9349 => x"65",
          9350 => x"73",
          9351 => x"76",
          9352 => x"64",
          9353 => x"00",
          9354 => x"73",
          9355 => x"6f",
          9356 => x"6e",
          9357 => x"65",
          9358 => x"00",
          9359 => x"20",
          9360 => x"70",
          9361 => x"62",
          9362 => x"66",
          9363 => x"73",
          9364 => x"65",
          9365 => x"6f",
          9366 => x"20",
          9367 => x"64",
          9368 => x"2e",
          9369 => x"00",
          9370 => x"72",
          9371 => x"20",
          9372 => x"72",
          9373 => x"2e",
          9374 => x"00",
          9375 => x"6d",
          9376 => x"74",
          9377 => x"70",
          9378 => x"74",
          9379 => x"20",
          9380 => x"63",
          9381 => x"65",
          9382 => x"00",
          9383 => x"6c",
          9384 => x"73",
          9385 => x"63",
          9386 => x"2e",
          9387 => x"00",
          9388 => x"73",
          9389 => x"69",
          9390 => x"6e",
          9391 => x"65",
          9392 => x"79",
          9393 => x"00",
          9394 => x"6f",
          9395 => x"6e",
          9396 => x"70",
          9397 => x"66",
          9398 => x"73",
          9399 => x"00",
          9400 => x"72",
          9401 => x"74",
          9402 => x"20",
          9403 => x"6f",
          9404 => x"63",
          9405 => x"00",
          9406 => x"63",
          9407 => x"73",
          9408 => x"00",
          9409 => x"6b",
          9410 => x"6e",
          9411 => x"72",
          9412 => x"0a",
          9413 => x"6c",
          9414 => x"79",
          9415 => x"20",
          9416 => x"61",
          9417 => x"6c",
          9418 => x"79",
          9419 => x"2f",
          9420 => x"2e",
          9421 => x"00",
          9422 => x"61",
          9423 => x"00",
          9424 => x"38",
          9425 => x"00",
          9426 => x"20",
          9427 => x"34",
          9428 => x"00",
          9429 => x"20",
          9430 => x"20",
          9431 => x"00",
          9432 => x"32",
          9433 => x"00",
          9434 => x"00",
          9435 => x"00",
          9436 => x"0a",
          9437 => x"55",
          9438 => x"00",
          9439 => x"2a",
          9440 => x"20",
          9441 => x"00",
          9442 => x"2f",
          9443 => x"32",
          9444 => x"00",
          9445 => x"2e",
          9446 => x"00",
          9447 => x"50",
          9448 => x"72",
          9449 => x"25",
          9450 => x"29",
          9451 => x"20",
          9452 => x"2a",
          9453 => x"00",
          9454 => x"55",
          9455 => x"49",
          9456 => x"72",
          9457 => x"74",
          9458 => x"6e",
          9459 => x"72",
          9460 => x"00",
          9461 => x"6d",
          9462 => x"69",
          9463 => x"72",
          9464 => x"74",
          9465 => x"00",
          9466 => x"32",
          9467 => x"74",
          9468 => x"75",
          9469 => x"00",
          9470 => x"43",
          9471 => x"52",
          9472 => x"6e",
          9473 => x"72",
          9474 => x"0a",
          9475 => x"43",
          9476 => x"57",
          9477 => x"6e",
          9478 => x"72",
          9479 => x"0a",
          9480 => x"52",
          9481 => x"52",
          9482 => x"6e",
          9483 => x"72",
          9484 => x"0a",
          9485 => x"52",
          9486 => x"54",
          9487 => x"6e",
          9488 => x"72",
          9489 => x"0a",
          9490 => x"52",
          9491 => x"52",
          9492 => x"6e",
          9493 => x"72",
          9494 => x"0a",
          9495 => x"52",
          9496 => x"54",
          9497 => x"6e",
          9498 => x"72",
          9499 => x"0a",
          9500 => x"74",
          9501 => x"67",
          9502 => x"20",
          9503 => x"65",
          9504 => x"2e",
          9505 => x"00",
          9506 => x"61",
          9507 => x"6e",
          9508 => x"69",
          9509 => x"2e",
          9510 => x"00",
          9511 => x"74",
          9512 => x"65",
          9513 => x"61",
          9514 => x"00",
          9515 => x"00",
          9516 => x"69",
          9517 => x"20",
          9518 => x"69",
          9519 => x"69",
          9520 => x"73",
          9521 => x"64",
          9522 => x"72",
          9523 => x"2c",
          9524 => x"65",
          9525 => x"20",
          9526 => x"74",
          9527 => x"6e",
          9528 => x"6c",
          9529 => x"00",
          9530 => x"00",
          9531 => x"64",
          9532 => x"73",
          9533 => x"64",
          9534 => x"00",
          9535 => x"69",
          9536 => x"6c",
          9537 => x"64",
          9538 => x"00",
          9539 => x"69",
          9540 => x"20",
          9541 => x"69",
          9542 => x"69",
          9543 => x"73",
          9544 => x"00",
          9545 => x"3d",
          9546 => x"00",
          9547 => x"3a",
          9548 => x"65",
          9549 => x"6e",
          9550 => x"2e",
          9551 => x"00",
          9552 => x"70",
          9553 => x"67",
          9554 => x"00",
          9555 => x"6d",
          9556 => x"69",
          9557 => x"2e",
          9558 => x"00",
          9559 => x"38",
          9560 => x"25",
          9561 => x"29",
          9562 => x"30",
          9563 => x"28",
          9564 => x"78",
          9565 => x"00",
          9566 => x"6d",
          9567 => x"65",
          9568 => x"79",
          9569 => x"00",
          9570 => x"6f",
          9571 => x"65",
          9572 => x"0a",
          9573 => x"38",
          9574 => x"30",
          9575 => x"00",
          9576 => x"3f",
          9577 => x"00",
          9578 => x"38",
          9579 => x"30",
          9580 => x"00",
          9581 => x"38",
          9582 => x"30",
          9583 => x"00",
          9584 => x"73",
          9585 => x"69",
          9586 => x"69",
          9587 => x"72",
          9588 => x"74",
          9589 => x"00",
          9590 => x"61",
          9591 => x"6e",
          9592 => x"6e",
          9593 => x"72",
          9594 => x"73",
          9595 => x"00",
          9596 => x"73",
          9597 => x"65",
          9598 => x"61",
          9599 => x"66",
          9600 => x"0a",
          9601 => x"61",
          9602 => x"6e",
          9603 => x"61",
          9604 => x"66",
          9605 => x"0a",
          9606 => x"65",
          9607 => x"69",
          9608 => x"63",
          9609 => x"20",
          9610 => x"30",
          9611 => x"2e",
          9612 => x"00",
          9613 => x"6c",
          9614 => x"67",
          9615 => x"64",
          9616 => x"20",
          9617 => x"78",
          9618 => x"2e",
          9619 => x"00",
          9620 => x"6c",
          9621 => x"65",
          9622 => x"6e",
          9623 => x"63",
          9624 => x"20",
          9625 => x"29",
          9626 => x"00",
          9627 => x"73",
          9628 => x"74",
          9629 => x"20",
          9630 => x"6c",
          9631 => x"74",
          9632 => x"2e",
          9633 => x"00",
          9634 => x"6c",
          9635 => x"65",
          9636 => x"74",
          9637 => x"2e",
          9638 => x"00",
          9639 => x"55",
          9640 => x"6e",
          9641 => x"3a",
          9642 => x"5c",
          9643 => x"25",
          9644 => x"00",
          9645 => x"3a",
          9646 => x"5c",
          9647 => x"00",
          9648 => x"3a",
          9649 => x"00",
          9650 => x"64",
          9651 => x"6d",
          9652 => x"64",
          9653 => x"00",
          9654 => x"6e",
          9655 => x"67",
          9656 => x"0a",
          9657 => x"61",
          9658 => x"6e",
          9659 => x"6e",
          9660 => x"72",
          9661 => x"73",
          9662 => x"0a",
          9663 => x"00",
          9664 => x"00",
          9665 => x"7f",
          9666 => x"00",
          9667 => x"7f",
          9668 => x"00",
          9669 => x"7f",
          9670 => x"00",
          9671 => x"00",
          9672 => x"00",
          9673 => x"ff",
          9674 => x"00",
          9675 => x"00",
          9676 => x"78",
          9677 => x"00",
          9678 => x"e1",
          9679 => x"e1",
          9680 => x"e1",
          9681 => x"00",
          9682 => x"01",
          9683 => x"01",
          9684 => x"10",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"87",
          9690 => x"87",
          9691 => x"87",
          9692 => x"87",
          9693 => x"7e",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"7e",
          9718 => x"00",
          9719 => x"7e",
          9720 => x"00",
          9721 => x"7e",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"80",
          9726 => x"01",
          9727 => x"00",
          9728 => x"00",
          9729 => x"80",
          9730 => x"01",
          9731 => x"00",
          9732 => x"00",
          9733 => x"80",
          9734 => x"03",
          9735 => x"00",
          9736 => x"00",
          9737 => x"80",
          9738 => x"03",
          9739 => x"00",
          9740 => x"00",
          9741 => x"80",
          9742 => x"03",
          9743 => x"00",
          9744 => x"00",
          9745 => x"80",
          9746 => x"04",
          9747 => x"00",
          9748 => x"00",
          9749 => x"80",
          9750 => x"04",
          9751 => x"00",
          9752 => x"00",
          9753 => x"80",
          9754 => x"04",
          9755 => x"00",
          9756 => x"00",
          9757 => x"80",
          9758 => x"04",
          9759 => x"00",
          9760 => x"00",
          9761 => x"80",
          9762 => x"04",
          9763 => x"00",
          9764 => x"00",
          9765 => x"80",
          9766 => x"04",
          9767 => x"00",
          9768 => x"00",
          9769 => x"80",
          9770 => x"04",
          9771 => x"00",
          9772 => x"00",
          9773 => x"80",
          9774 => x"05",
          9775 => x"00",
          9776 => x"00",
          9777 => x"80",
          9778 => x"05",
          9779 => x"00",
          9780 => x"00",
          9781 => x"81",
          9782 => x"05",
          9783 => x"00",
          9784 => x"00",
          9785 => x"81",
          9786 => x"05",
          9787 => x"00",
          9788 => x"00",
          9789 => x"81",
          9790 => x"07",
          9791 => x"00",
          9792 => x"00",
          9793 => x"81",
          9794 => x"07",
          9795 => x"00",
          9796 => x"00",
          9797 => x"81",
          9798 => x"08",
          9799 => x"00",
          9800 => x"00",
          9801 => x"81",
          9802 => x"08",
          9803 => x"00",
          9804 => x"00",
          9805 => x"81",
          9806 => x"08",
          9807 => x"00",
          9808 => x"00",
          9809 => x"81",
          9810 => x"08",
          9811 => x"00",
          9812 => x"00",
          9813 => x"81",
          9814 => x"09",
          9815 => x"00",
          9816 => x"00",
          9817 => x"81",
          9818 => x"09",
          9819 => x"00",
          9820 => x"00",
          9821 => x"81",
          9822 => x"09",
          9823 => x"00",
          9824 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"04",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"08",
             9 => x"08",
            10 => x"88",
            11 => x"90",
            12 => x"88",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"fd",
            17 => x"83",
            18 => x"05",
            19 => x"2b",
            20 => x"ff",
            21 => x"00",
            22 => x"00",
            23 => x"00",
            24 => x"fd",
            25 => x"ff",
            26 => x"06",
            27 => x"82",
            28 => x"2b",
            29 => x"83",
            30 => x"0b",
            31 => x"a5",
            32 => x"09",
            33 => x"05",
            34 => x"06",
            35 => x"09",
            36 => x"0a",
            37 => x"51",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"2e",
            42 => x"04",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"73",
            49 => x"06",
            50 => x"81",
            51 => x"10",
            52 => x"10",
            53 => x"0a",
            54 => x"51",
            55 => x"00",
            56 => x"72",
            57 => x"2e",
            58 => x"04",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"04",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"0a",
            81 => x"53",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"81",
            90 => x"0b",
            91 => x"04",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"9f",
            98 => x"74",
            99 => x"06",
           100 => x"07",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"06",
           106 => x"09",
           107 => x"05",
           108 => x"2b",
           109 => x"06",
           110 => x"04",
           111 => x"00",
           112 => x"09",
           113 => x"05",
           114 => x"05",
           115 => x"81",
           116 => x"04",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"09",
           121 => x"05",
           122 => x"05",
           123 => x"09",
           124 => x"51",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"09",
           129 => x"04",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"00",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"09",
           145 => x"73",
           146 => x"53",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"fc",
           153 => x"83",
           154 => x"05",
           155 => x"10",
           156 => x"ff",
           157 => x"00",
           158 => x"00",
           159 => x"00",
           160 => x"fc",
           161 => x"0b",
           162 => x"73",
           163 => x"10",
           164 => x"0b",
           165 => x"ac",
           166 => x"00",
           167 => x"00",
           168 => x"08",
           169 => x"08",
           170 => x"0b",
           171 => x"2d",
           172 => x"08",
           173 => x"8c",
           174 => x"51",
           175 => x"00",
           176 => x"08",
           177 => x"08",
           178 => x"0b",
           179 => x"2d",
           180 => x"08",
           181 => x"8c",
           182 => x"51",
           183 => x"00",
           184 => x"09",
           185 => x"09",
           186 => x"06",
           187 => x"54",
           188 => x"09",
           189 => x"ff",
           190 => x"51",
           191 => x"00",
           192 => x"09",
           193 => x"09",
           194 => x"81",
           195 => x"70",
           196 => x"73",
           197 => x"05",
           198 => x"07",
           199 => x"04",
           200 => x"ff",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"00",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"81",
           217 => x"00",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"00",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"84",
           233 => x"10",
           234 => x"00",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"71",
           250 => x"0d",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"00",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"04",
           267 => x"81",
           268 => x"83",
           269 => x"05",
           270 => x"10",
           271 => x"72",
           272 => x"51",
           273 => x"72",
           274 => x"06",
           275 => x"72",
           276 => x"10",
           277 => x"10",
           278 => x"ed",
           279 => x"53",
           280 => x"f4",
           281 => x"27",
           282 => x"71",
           283 => x"53",
           284 => x"0b",
           285 => x"88",
           286 => x"9d",
           287 => x"04",
           288 => x"04",
           289 => x"94",
           290 => x"0c",
           291 => x"80",
           292 => x"8c",
           293 => x"94",
           294 => x"08",
           295 => x"3f",
           296 => x"88",
           297 => x"3d",
           298 => x"04",
           299 => x"94",
           300 => x"0d",
           301 => x"08",
           302 => x"52",
           303 => x"05",
           304 => x"b9",
           305 => x"70",
           306 => x"85",
           307 => x"0c",
           308 => x"02",
           309 => x"3d",
           310 => x"94",
           311 => x"0c",
           312 => x"05",
           313 => x"ab",
           314 => x"88",
           315 => x"94",
           316 => x"0c",
           317 => x"08",
           318 => x"94",
           319 => x"08",
           320 => x"0b",
           321 => x"05",
           322 => x"f4",
           323 => x"08",
           324 => x"94",
           325 => x"08",
           326 => x"38",
           327 => x"05",
           328 => x"08",
           329 => x"80",
           330 => x"f0",
           331 => x"08",
           332 => x"88",
           333 => x"94",
           334 => x"0c",
           335 => x"05",
           336 => x"fc",
           337 => x"53",
           338 => x"05",
           339 => x"08",
           340 => x"51",
           341 => x"88",
           342 => x"08",
           343 => x"54",
           344 => x"05",
           345 => x"8c",
           346 => x"f8",
           347 => x"94",
           348 => x"0c",
           349 => x"05",
           350 => x"0c",
           351 => x"0d",
           352 => x"94",
           353 => x"0c",
           354 => x"80",
           355 => x"fc",
           356 => x"08",
           357 => x"80",
           358 => x"94",
           359 => x"08",
           360 => x"88",
           361 => x"0b",
           362 => x"05",
           363 => x"8c",
           364 => x"25",
           365 => x"08",
           366 => x"30",
           367 => x"05",
           368 => x"94",
           369 => x"08",
           370 => x"88",
           371 => x"ad",
           372 => x"70",
           373 => x"05",
           374 => x"08",
           375 => x"80",
           376 => x"94",
           377 => x"08",
           378 => x"f8",
           379 => x"08",
           380 => x"70",
           381 => x"87",
           382 => x"0c",
           383 => x"02",
           384 => x"3d",
           385 => x"94",
           386 => x"0c",
           387 => x"08",
           388 => x"94",
           389 => x"08",
           390 => x"05",
           391 => x"38",
           392 => x"05",
           393 => x"a3",
           394 => x"94",
           395 => x"08",
           396 => x"94",
           397 => x"08",
           398 => x"8c",
           399 => x"08",
           400 => x"10",
           401 => x"05",
           402 => x"94",
           403 => x"08",
           404 => x"c9",
           405 => x"8c",
           406 => x"08",
           407 => x"26",
           408 => x"08",
           409 => x"94",
           410 => x"08",
           411 => x"88",
           412 => x"08",
           413 => x"94",
           414 => x"08",
           415 => x"f8",
           416 => x"08",
           417 => x"81",
           418 => x"fc",
           419 => x"08",
           420 => x"81",
           421 => x"8c",
           422 => x"af",
           423 => x"90",
           424 => x"2e",
           425 => x"08",
           426 => x"70",
           427 => x"05",
           428 => x"39",
           429 => x"05",
           430 => x"08",
           431 => x"51",
           432 => x"05",
           433 => x"85",
           434 => x"0c",
           435 => x"0d",
           436 => x"87",
           437 => x"0c",
           438 => x"c0",
           439 => x"85",
           440 => x"98",
           441 => x"c0",
           442 => x"70",
           443 => x"51",
           444 => x"8a",
           445 => x"98",
           446 => x"70",
           447 => x"c0",
           448 => x"fc",
           449 => x"52",
           450 => x"87",
           451 => x"08",
           452 => x"2e",
           453 => x"0b",
           454 => x"f0",
           455 => x"0b",
           456 => x"88",
           457 => x"0d",
           458 => x"0d",
           459 => x"56",
           460 => x"0b",
           461 => x"9f",
           462 => x"06",
           463 => x"52",
           464 => x"09",
           465 => x"9e",
           466 => x"87",
           467 => x"0c",
           468 => x"92",
           469 => x"0b",
           470 => x"8c",
           471 => x"92",
           472 => x"85",
           473 => x"06",
           474 => x"70",
           475 => x"38",
           476 => x"84",
           477 => x"ff",
           478 => x"27",
           479 => x"73",
           480 => x"38",
           481 => x"8b",
           482 => x"70",
           483 => x"34",
           484 => x"81",
           485 => x"a2",
           486 => x"80",
           487 => x"87",
           488 => x"08",
           489 => x"b5",
           490 => x"98",
           491 => x"70",
           492 => x"0b",
           493 => x"8c",
           494 => x"92",
           495 => x"82",
           496 => x"70",
           497 => x"73",
           498 => x"06",
           499 => x"72",
           500 => x"06",
           501 => x"c0",
           502 => x"51",
           503 => x"09",
           504 => x"38",
           505 => x"88",
           506 => x"0d",
           507 => x"0d",
           508 => x"33",
           509 => x"88",
           510 => x"0c",
           511 => x"3d",
           512 => x"3d",
           513 => x"11",
           514 => x"33",
           515 => x"71",
           516 => x"81",
           517 => x"72",
           518 => x"75",
           519 => x"88",
           520 => x"54",
           521 => x"85",
           522 => x"f9",
           523 => x"0b",
           524 => x"f4",
           525 => x"81",
           526 => x"ed",
           527 => x"17",
           528 => x"e5",
           529 => x"55",
           530 => x"89",
           531 => x"2e",
           532 => x"d5",
           533 => x"76",
           534 => x"06",
           535 => x"2a",
           536 => x"05",
           537 => x"70",
           538 => x"bd",
           539 => x"b9",
           540 => x"fe",
           541 => x"08",
           542 => x"06",
           543 => x"84",
           544 => x"2b",
           545 => x"53",
           546 => x"8c",
           547 => x"52",
           548 => x"52",
           549 => x"3f",
           550 => x"38",
           551 => x"e2",
           552 => x"f0",
           553 => x"83",
           554 => x"74",
           555 => x"3d",
           556 => x"3d",
           557 => x"0b",
           558 => x"fe",
           559 => x"08",
           560 => x"56",
           561 => x"74",
           562 => x"38",
           563 => x"75",
           564 => x"16",
           565 => x"53",
           566 => x"87",
           567 => x"fd",
           568 => x"54",
           569 => x"0b",
           570 => x"08",
           571 => x"53",
           572 => x"2e",
           573 => x"8c",
           574 => x"51",
           575 => x"88",
           576 => x"53",
           577 => x"fd",
           578 => x"08",
           579 => x"06",
           580 => x"0c",
           581 => x"04",
           582 => x"76",
           583 => x"9f",
           584 => x"55",
           585 => x"88",
           586 => x"72",
           587 => x"38",
           588 => x"73",
           589 => x"81",
           590 => x"72",
           591 => x"33",
           592 => x"2e",
           593 => x"85",
           594 => x"08",
           595 => x"16",
           596 => x"2e",
           597 => x"51",
           598 => x"88",
           599 => x"39",
           600 => x"52",
           601 => x"0c",
           602 => x"88",
           603 => x"0d",
           604 => x"0d",
           605 => x"0b",
           606 => x"71",
           607 => x"70",
           608 => x"06",
           609 => x"55",
           610 => x"88",
           611 => x"08",
           612 => x"38",
           613 => x"dc",
           614 => x"06",
           615 => x"cf",
           616 => x"90",
           617 => x"15",
           618 => x"8f",
           619 => x"84",
           620 => x"52",
           621 => x"bc",
           622 => x"82",
           623 => x"05",
           624 => x"06",
           625 => x"38",
           626 => x"df",
           627 => x"71",
           628 => x"a0",
           629 => x"88",
           630 => x"08",
           631 => x"88",
           632 => x"0c",
           633 => x"fd",
           634 => x"08",
           635 => x"73",
           636 => x"52",
           637 => x"88",
           638 => x"f2",
           639 => x"62",
           640 => x"5c",
           641 => x"74",
           642 => x"81",
           643 => x"81",
           644 => x"56",
           645 => x"70",
           646 => x"74",
           647 => x"81",
           648 => x"81",
           649 => x"0b",
           650 => x"62",
           651 => x"55",
           652 => x"8f",
           653 => x"fd",
           654 => x"08",
           655 => x"34",
           656 => x"93",
           657 => x"08",
           658 => x"5f",
           659 => x"76",
           660 => x"58",
           661 => x"55",
           662 => x"09",
           663 => x"38",
           664 => x"5b",
           665 => x"5f",
           666 => x"1c",
           667 => x"06",
           668 => x"33",
           669 => x"70",
           670 => x"27",
           671 => x"07",
           672 => x"5b",
           673 => x"55",
           674 => x"38",
           675 => x"09",
           676 => x"38",
           677 => x"7a",
           678 => x"55",
           679 => x"9f",
           680 => x"32",
           681 => x"ae",
           682 => x"70",
           683 => x"2a",
           684 => x"51",
           685 => x"38",
           686 => x"5a",
           687 => x"77",
           688 => x"81",
           689 => x"1c",
           690 => x"55",
           691 => x"ff",
           692 => x"1e",
           693 => x"55",
           694 => x"83",
           695 => x"74",
           696 => x"7b",
           697 => x"3f",
           698 => x"ef",
           699 => x"7b",
           700 => x"2b",
           701 => x"54",
           702 => x"08",
           703 => x"f8",
           704 => x"08",
           705 => x"80",
           706 => x"33",
           707 => x"2e",
           708 => x"8b",
           709 => x"83",
           710 => x"06",
           711 => x"74",
           712 => x"7d",
           713 => x"88",
           714 => x"5b",
           715 => x"58",
           716 => x"9a",
           717 => x"81",
           718 => x"79",
           719 => x"5b",
           720 => x"31",
           721 => x"75",
           722 => x"38",
           723 => x"80",
           724 => x"7b",
           725 => x"3f",
           726 => x"88",
           727 => x"08",
           728 => x"39",
           729 => x"1c",
           730 => x"33",
           731 => x"a5",
           732 => x"33",
           733 => x"70",
           734 => x"56",
           735 => x"38",
           736 => x"39",
           737 => x"39",
           738 => x"d3",
           739 => x"88",
           740 => x"af",
           741 => x"0c",
           742 => x"04",
           743 => x"79",
           744 => x"82",
           745 => x"53",
           746 => x"51",
           747 => x"83",
           748 => x"80",
           749 => x"51",
           750 => x"88",
           751 => x"ff",
           752 => x"56",
           753 => x"d5",
           754 => x"06",
           755 => x"75",
           756 => x"77",
           757 => x"f6",
           758 => x"08",
           759 => x"94",
           760 => x"f8",
           761 => x"08",
           762 => x"06",
           763 => x"82",
           764 => x"38",
           765 => x"d2",
           766 => x"76",
           767 => x"3f",
           768 => x"88",
           769 => x"76",
           770 => x"3f",
           771 => x"ff",
           772 => x"74",
           773 => x"2e",
           774 => x"56",
           775 => x"89",
           776 => x"ed",
           777 => x"59",
           778 => x"0b",
           779 => x"0c",
           780 => x"88",
           781 => x"55",
           782 => x"82",
           783 => x"75",
           784 => x"70",
           785 => x"fe",
           786 => x"08",
           787 => x"57",
           788 => x"09",
           789 => x"38",
           790 => x"be",
           791 => x"75",
           792 => x"3f",
           793 => x"38",
           794 => x"55",
           795 => x"ac",
           796 => x"e4",
           797 => x"8a",
           798 => x"88",
           799 => x"52",
           800 => x"3f",
           801 => x"ff",
           802 => x"83",
           803 => x"06",
           804 => x"56",
           805 => x"76",
           806 => x"38",
           807 => x"8f",
           808 => x"8d",
           809 => x"75",
           810 => x"3f",
           811 => x"08",
           812 => x"95",
           813 => x"51",
           814 => x"88",
           815 => x"ff",
           816 => x"8c",
           817 => x"f3",
           818 => x"b6",
           819 => x"58",
           820 => x"33",
           821 => x"02",
           822 => x"05",
           823 => x"59",
           824 => x"3f",
           825 => x"ff",
           826 => x"05",
           827 => x"8c",
           828 => x"1a",
           829 => x"e0",
           830 => x"f1",
           831 => x"84",
           832 => x"3d",
           833 => x"f5",
           834 => x"08",
           835 => x"06",
           836 => x"38",
           837 => x"05",
           838 => x"3f",
           839 => x"7a",
           840 => x"3f",
           841 => x"ff",
           842 => x"71",
           843 => x"84",
           844 => x"84",
           845 => x"33",
           846 => x"31",
           847 => x"51",
           848 => x"3f",
           849 => x"05",
           850 => x"0c",
           851 => x"8a",
           852 => x"74",
           853 => x"26",
           854 => x"57",
           855 => x"76",
           856 => x"83",
           857 => x"86",
           858 => x"2e",
           859 => x"76",
           860 => x"83",
           861 => x"06",
           862 => x"3d",
           863 => x"f5",
           864 => x"08",
           865 => x"88",
           866 => x"08",
           867 => x"0c",
           868 => x"ff",
           869 => x"08",
           870 => x"2a",
           871 => x"0c",
           872 => x"81",
           873 => x"0b",
           874 => x"f4",
           875 => x"75",
           876 => x"3d",
           877 => x"3d",
           878 => x"0b",
           879 => x"55",
           880 => x"80",
           881 => x"38",
           882 => x"16",
           883 => x"e0",
           884 => x"54",
           885 => x"54",
           886 => x"51",
           887 => x"88",
           888 => x"08",
           889 => x"88",
           890 => x"73",
           891 => x"38",
           892 => x"33",
           893 => x"70",
           894 => x"55",
           895 => x"2e",
           896 => x"54",
           897 => x"51",
           898 => x"88",
           899 => x"0c",
           900 => x"05",
           901 => x"3f",
           902 => x"16",
           903 => x"16",
           904 => x"81",
           905 => x"88",
           906 => x"0d",
           907 => x"0d",
           908 => x"0b",
           909 => x"f4",
           910 => x"5c",
           911 => x"0c",
           912 => x"80",
           913 => x"38",
           914 => x"81",
           915 => x"57",
           916 => x"81",
           917 => x"39",
           918 => x"34",
           919 => x"0b",
           920 => x"81",
           921 => x"39",
           922 => x"98",
           923 => x"55",
           924 => x"83",
           925 => x"77",
           926 => x"9a",
           927 => x"08",
           928 => x"06",
           929 => x"80",
           930 => x"16",
           931 => x"77",
           932 => x"70",
           933 => x"5b",
           934 => x"38",
           935 => x"a0",
           936 => x"8b",
           937 => x"08",
           938 => x"3f",
           939 => x"81",
           940 => x"aa",
           941 => x"17",
           942 => x"08",
           943 => x"3f",
           944 => x"88",
           945 => x"ff",
           946 => x"08",
           947 => x"0c",
           948 => x"83",
           949 => x"80",
           950 => x"55",
           951 => x"83",
           952 => x"74",
           953 => x"08",
           954 => x"53",
           955 => x"52",
           956 => x"b5",
           957 => x"fe",
           958 => x"16",
           959 => x"17",
           960 => x"31",
           961 => x"7c",
           962 => x"80",
           963 => x"38",
           964 => x"fe",
           965 => x"57",
           966 => x"8c",
           967 => x"fb",
           968 => x"c0",
           969 => x"54",
           970 => x"52",
           971 => x"d7",
           972 => x"90",
           973 => x"94",
           974 => x"54",
           975 => x"52",
           976 => x"c3",
           977 => x"08",
           978 => x"94",
           979 => x"c0",
           980 => x"54",
           981 => x"52",
           982 => x"ab",
           983 => x"90",
           984 => x"94",
           985 => x"54",
           986 => x"52",
           987 => x"97",
           988 => x"08",
           989 => x"94",
           990 => x"80",
           991 => x"c0",
           992 => x"8c",
           993 => x"87",
           994 => x"0c",
           995 => x"f9",
           996 => x"08",
           997 => x"e0",
           998 => x"3f",
           999 => x"38",
          1000 => x"88",
          1001 => x"98",
          1002 => x"87",
          1003 => x"53",
          1004 => x"74",
          1005 => x"3f",
          1006 => x"38",
          1007 => x"80",
          1008 => x"73",
          1009 => x"39",
          1010 => x"73",
          1011 => x"fb",
          1012 => x"ff",
          1013 => x"00",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"4f",
          1017 => x"49",
          1018 => x"52",
          1019 => x"00",
          1020 => x"00",
          2048 => x"0b",
          2049 => x"0b",
          2050 => x"aa",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"04",
          2058 => x"a4",
          2059 => x"0b",
          2060 => x"04",
          2061 => x"a4",
          2062 => x"0b",
          2063 => x"04",
          2064 => x"a4",
          2065 => x"0b",
          2066 => x"04",
          2067 => x"a4",
          2068 => x"0b",
          2069 => x"04",
          2070 => x"a5",
          2071 => x"0b",
          2072 => x"04",
          2073 => x"a5",
          2074 => x"0b",
          2075 => x"04",
          2076 => x"a5",
          2077 => x"0b",
          2078 => x"04",
          2079 => x"a5",
          2080 => x"0b",
          2081 => x"04",
          2082 => x"a6",
          2083 => x"0b",
          2084 => x"04",
          2085 => x"a6",
          2086 => x"0b",
          2087 => x"04",
          2088 => x"a6",
          2089 => x"0b",
          2090 => x"04",
          2091 => x"a6",
          2092 => x"0b",
          2093 => x"04",
          2094 => x"a6",
          2095 => x"0b",
          2096 => x"04",
          2097 => x"a7",
          2098 => x"0b",
          2099 => x"04",
          2100 => x"a7",
          2101 => x"0b",
          2102 => x"04",
          2103 => x"a7",
          2104 => x"0b",
          2105 => x"04",
          2106 => x"a7",
          2107 => x"0b",
          2108 => x"04",
          2109 => x"a8",
          2110 => x"0b",
          2111 => x"04",
          2112 => x"a8",
          2113 => x"0b",
          2114 => x"04",
          2115 => x"a8",
          2116 => x"0b",
          2117 => x"04",
          2118 => x"a8",
          2119 => x"0b",
          2120 => x"04",
          2121 => x"a9",
          2122 => x"0b",
          2123 => x"04",
          2124 => x"a9",
          2125 => x"0b",
          2126 => x"04",
          2127 => x"a9",
          2128 => x"0b",
          2129 => x"04",
          2130 => x"a9",
          2131 => x"0b",
          2132 => x"04",
          2133 => x"aa",
          2134 => x"0b",
          2135 => x"04",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"a4",
          2177 => x"93",
          2178 => x"a0",
          2179 => x"90",
          2180 => x"90",
          2181 => x"90",
          2182 => x"eb",
          2183 => x"90",
          2184 => x"90",
          2185 => x"90",
          2186 => x"aa",
          2187 => x"90",
          2188 => x"90",
          2189 => x"90",
          2190 => x"c8",
          2191 => x"90",
          2192 => x"90",
          2193 => x"90",
          2194 => x"86",
          2195 => x"90",
          2196 => x"90",
          2197 => x"90",
          2198 => x"84",
          2199 => x"90",
          2200 => x"90",
          2201 => x"90",
          2202 => x"eb",
          2203 => x"90",
          2204 => x"90",
          2205 => x"90",
          2206 => x"a1",
          2207 => x"90",
          2208 => x"90",
          2209 => x"90",
          2210 => x"93",
          2211 => x"90",
          2212 => x"90",
          2213 => x"90",
          2214 => x"ac",
          2215 => x"90",
          2216 => x"90",
          2217 => x"90",
          2218 => x"9d",
          2219 => x"90",
          2220 => x"90",
          2221 => x"90",
          2222 => x"c2",
          2223 => x"90",
          2224 => x"90",
          2225 => x"90",
          2226 => x"e6",
          2227 => x"90",
          2228 => x"90",
          2229 => x"90",
          2230 => x"2d",
          2231 => x"08",
          2232 => x"04",
          2233 => x"0c",
          2234 => x"82",
          2235 => x"83",
          2236 => x"82",
          2237 => x"b3",
          2238 => x"93",
          2239 => x"80",
          2240 => x"93",
          2241 => x"cf",
          2242 => x"90",
          2243 => x"90",
          2244 => x"90",
          2245 => x"2d",
          2246 => x"08",
          2247 => x"04",
          2248 => x"0c",
          2249 => x"2d",
          2250 => x"08",
          2251 => x"04",
          2252 => x"0c",
          2253 => x"2d",
          2254 => x"08",
          2255 => x"04",
          2256 => x"0c",
          2257 => x"2d",
          2258 => x"08",
          2259 => x"04",
          2260 => x"0c",
          2261 => x"2d",
          2262 => x"08",
          2263 => x"04",
          2264 => x"0c",
          2265 => x"2d",
          2266 => x"08",
          2267 => x"04",
          2268 => x"0c",
          2269 => x"2d",
          2270 => x"08",
          2271 => x"04",
          2272 => x"0c",
          2273 => x"2d",
          2274 => x"08",
          2275 => x"04",
          2276 => x"0c",
          2277 => x"2d",
          2278 => x"08",
          2279 => x"04",
          2280 => x"0c",
          2281 => x"2d",
          2282 => x"08",
          2283 => x"04",
          2284 => x"0c",
          2285 => x"2d",
          2286 => x"08",
          2287 => x"04",
          2288 => x"0c",
          2289 => x"2d",
          2290 => x"08",
          2291 => x"04",
          2292 => x"0c",
          2293 => x"2d",
          2294 => x"08",
          2295 => x"04",
          2296 => x"0c",
          2297 => x"2d",
          2298 => x"08",
          2299 => x"04",
          2300 => x"0c",
          2301 => x"2d",
          2302 => x"08",
          2303 => x"04",
          2304 => x"0c",
          2305 => x"2d",
          2306 => x"08",
          2307 => x"04",
          2308 => x"0c",
          2309 => x"2d",
          2310 => x"08",
          2311 => x"04",
          2312 => x"0c",
          2313 => x"2d",
          2314 => x"08",
          2315 => x"04",
          2316 => x"0c",
          2317 => x"2d",
          2318 => x"08",
          2319 => x"04",
          2320 => x"0c",
          2321 => x"2d",
          2322 => x"08",
          2323 => x"04",
          2324 => x"0c",
          2325 => x"2d",
          2326 => x"08",
          2327 => x"04",
          2328 => x"0c",
          2329 => x"2d",
          2330 => x"08",
          2331 => x"04",
          2332 => x"0c",
          2333 => x"2d",
          2334 => x"08",
          2335 => x"04",
          2336 => x"0c",
          2337 => x"2d",
          2338 => x"08",
          2339 => x"04",
          2340 => x"0c",
          2341 => x"2d",
          2342 => x"08",
          2343 => x"04",
          2344 => x"0c",
          2345 => x"2d",
          2346 => x"08",
          2347 => x"04",
          2348 => x"0c",
          2349 => x"2d",
          2350 => x"08",
          2351 => x"04",
          2352 => x"0c",
          2353 => x"2d",
          2354 => x"08",
          2355 => x"04",
          2356 => x"0c",
          2357 => x"2d",
          2358 => x"08",
          2359 => x"04",
          2360 => x"0c",
          2361 => x"2d",
          2362 => x"08",
          2363 => x"04",
          2364 => x"0c",
          2365 => x"2d",
          2366 => x"08",
          2367 => x"04",
          2368 => x"0c",
          2369 => x"82",
          2370 => x"83",
          2371 => x"82",
          2372 => x"b4",
          2373 => x"93",
          2374 => x"80",
          2375 => x"93",
          2376 => x"92",
          2377 => x"90",
          2378 => x"90",
          2379 => x"90",
          2380 => x"fb",
          2381 => x"90",
          2382 => x"90",
          2383 => x"84",
          2384 => x"c4",
          2385 => x"80",
          2386 => x"05",
          2387 => x"0b",
          2388 => x"04",
          2389 => x"81",
          2390 => x"3c",
          2391 => x"90",
          2392 => x"93",
          2393 => x"3d",
          2394 => x"82",
          2395 => x"8c",
          2396 => x"82",
          2397 => x"88",
          2398 => x"80",
          2399 => x"93",
          2400 => x"82",
          2401 => x"54",
          2402 => x"82",
          2403 => x"04",
          2404 => x"08",
          2405 => x"90",
          2406 => x"0d",
          2407 => x"93",
          2408 => x"05",
          2409 => x"93",
          2410 => x"05",
          2411 => x"3f",
          2412 => x"08",
          2413 => x"84",
          2414 => x"3d",
          2415 => x"90",
          2416 => x"93",
          2417 => x"82",
          2418 => x"fd",
          2419 => x"0b",
          2420 => x"08",
          2421 => x"80",
          2422 => x"90",
          2423 => x"0c",
          2424 => x"08",
          2425 => x"82",
          2426 => x"88",
          2427 => x"b9",
          2428 => x"90",
          2429 => x"08",
          2430 => x"38",
          2431 => x"93",
          2432 => x"05",
          2433 => x"38",
          2434 => x"08",
          2435 => x"10",
          2436 => x"08",
          2437 => x"82",
          2438 => x"fc",
          2439 => x"82",
          2440 => x"fc",
          2441 => x"b8",
          2442 => x"90",
          2443 => x"08",
          2444 => x"e1",
          2445 => x"90",
          2446 => x"08",
          2447 => x"08",
          2448 => x"26",
          2449 => x"93",
          2450 => x"05",
          2451 => x"90",
          2452 => x"08",
          2453 => x"90",
          2454 => x"0c",
          2455 => x"08",
          2456 => x"82",
          2457 => x"fc",
          2458 => x"82",
          2459 => x"f8",
          2460 => x"93",
          2461 => x"05",
          2462 => x"82",
          2463 => x"fc",
          2464 => x"93",
          2465 => x"05",
          2466 => x"82",
          2467 => x"8c",
          2468 => x"95",
          2469 => x"90",
          2470 => x"08",
          2471 => x"38",
          2472 => x"08",
          2473 => x"70",
          2474 => x"08",
          2475 => x"51",
          2476 => x"93",
          2477 => x"05",
          2478 => x"93",
          2479 => x"05",
          2480 => x"93",
          2481 => x"05",
          2482 => x"84",
          2483 => x"0d",
          2484 => x"0c",
          2485 => x"0d",
          2486 => x"7b",
          2487 => x"55",
          2488 => x"8c",
          2489 => x"07",
          2490 => x"70",
          2491 => x"38",
          2492 => x"71",
          2493 => x"38",
          2494 => x"05",
          2495 => x"70",
          2496 => x"34",
          2497 => x"71",
          2498 => x"81",
          2499 => x"74",
          2500 => x"0c",
          2501 => x"04",
          2502 => x"70",
          2503 => x"08",
          2504 => x"05",
          2505 => x"70",
          2506 => x"08",
          2507 => x"05",
          2508 => x"70",
          2509 => x"08",
          2510 => x"05",
          2511 => x"70",
          2512 => x"08",
          2513 => x"05",
          2514 => x"12",
          2515 => x"26",
          2516 => x"72",
          2517 => x"72",
          2518 => x"54",
          2519 => x"84",
          2520 => x"fc",
          2521 => x"83",
          2522 => x"70",
          2523 => x"39",
          2524 => x"76",
          2525 => x"8c",
          2526 => x"33",
          2527 => x"55",
          2528 => x"8a",
          2529 => x"06",
          2530 => x"2e",
          2531 => x"12",
          2532 => x"2e",
          2533 => x"73",
          2534 => x"55",
          2535 => x"52",
          2536 => x"09",
          2537 => x"38",
          2538 => x"84",
          2539 => x"0d",
          2540 => x"88",
          2541 => x"70",
          2542 => x"07",
          2543 => x"8f",
          2544 => x"38",
          2545 => x"84",
          2546 => x"72",
          2547 => x"05",
          2548 => x"71",
          2549 => x"53",
          2550 => x"70",
          2551 => x"0c",
          2552 => x"71",
          2553 => x"38",
          2554 => x"90",
          2555 => x"70",
          2556 => x"0c",
          2557 => x"71",
          2558 => x"38",
          2559 => x"8e",
          2560 => x"0d",
          2561 => x"70",
          2562 => x"06",
          2563 => x"55",
          2564 => x"38",
          2565 => x"70",
          2566 => x"fb",
          2567 => x"06",
          2568 => x"82",
          2569 => x"51",
          2570 => x"54",
          2571 => x"84",
          2572 => x"70",
          2573 => x"0c",
          2574 => x"09",
          2575 => x"fd",
          2576 => x"70",
          2577 => x"81",
          2578 => x"51",
          2579 => x"70",
          2580 => x"38",
          2581 => x"70",
          2582 => x"33",
          2583 => x"70",
          2584 => x"34",
          2585 => x"74",
          2586 => x"0c",
          2587 => x"04",
          2588 => x"75",
          2589 => x"06",
          2590 => x"70",
          2591 => x"70",
          2592 => x"f7",
          2593 => x"12",
          2594 => x"84",
          2595 => x"06",
          2596 => x"53",
          2597 => x"84",
          2598 => x"70",
          2599 => x"fd",
          2600 => x"70",
          2601 => x"81",
          2602 => x"51",
          2603 => x"80",
          2604 => x"72",
          2605 => x"51",
          2606 => x"8a",
          2607 => x"70",
          2608 => x"70",
          2609 => x"74",
          2610 => x"84",
          2611 => x"0d",
          2612 => x"0d",
          2613 => x"70",
          2614 => x"52",
          2615 => x"80",
          2616 => x"74",
          2617 => x"51",
          2618 => x"80",
          2619 => x"13",
          2620 => x"2e",
          2621 => x"33",
          2622 => x"51",
          2623 => x"09",
          2624 => x"38",
          2625 => x"81",
          2626 => x"81",
          2627 => x"70",
          2628 => x"fe",
          2629 => x"81",
          2630 => x"55",
          2631 => x"ff",
          2632 => x"06",
          2633 => x"33",
          2634 => x"51",
          2635 => x"06",
          2636 => x"06",
          2637 => x"51",
          2638 => x"82",
          2639 => x"88",
          2640 => x"71",
          2641 => x"83",
          2642 => x"38",
          2643 => x"08",
          2644 => x"74",
          2645 => x"ff",
          2646 => x"13",
          2647 => x"2e",
          2648 => x"08",
          2649 => x"fb",
          2650 => x"06",
          2651 => x"82",
          2652 => x"51",
          2653 => x"9a",
          2654 => x"84",
          2655 => x"83",
          2656 => x"38",
          2657 => x"08",
          2658 => x"74",
          2659 => x"fe",
          2660 => x"0b",
          2661 => x"0c",
          2662 => x"04",
          2663 => x"80",
          2664 => x"71",
          2665 => x"87",
          2666 => x"93",
          2667 => x"ff",
          2668 => x"ff",
          2669 => x"72",
          2670 => x"38",
          2671 => x"84",
          2672 => x"0d",
          2673 => x"0d",
          2674 => x"70",
          2675 => x"71",
          2676 => x"ca",
          2677 => x"51",
          2678 => x"09",
          2679 => x"38",
          2680 => x"f1",
          2681 => x"84",
          2682 => x"53",
          2683 => x"70",
          2684 => x"53",
          2685 => x"a0",
          2686 => x"81",
          2687 => x"2e",
          2688 => x"e5",
          2689 => x"ff",
          2690 => x"a0",
          2691 => x"06",
          2692 => x"73",
          2693 => x"55",
          2694 => x"0c",
          2695 => x"82",
          2696 => x"87",
          2697 => x"fc",
          2698 => x"53",
          2699 => x"2e",
          2700 => x"3d",
          2701 => x"72",
          2702 => x"3f",
          2703 => x"08",
          2704 => x"53",
          2705 => x"53",
          2706 => x"84",
          2707 => x"0d",
          2708 => x"0d",
          2709 => x"33",
          2710 => x"53",
          2711 => x"8b",
          2712 => x"38",
          2713 => x"ff",
          2714 => x"52",
          2715 => x"81",
          2716 => x"13",
          2717 => x"52",
          2718 => x"80",
          2719 => x"13",
          2720 => x"52",
          2721 => x"80",
          2722 => x"13",
          2723 => x"52",
          2724 => x"80",
          2725 => x"13",
          2726 => x"52",
          2727 => x"26",
          2728 => x"8a",
          2729 => x"87",
          2730 => x"e7",
          2731 => x"38",
          2732 => x"c0",
          2733 => x"72",
          2734 => x"98",
          2735 => x"13",
          2736 => x"98",
          2737 => x"13",
          2738 => x"98",
          2739 => x"13",
          2740 => x"98",
          2741 => x"13",
          2742 => x"98",
          2743 => x"13",
          2744 => x"98",
          2745 => x"87",
          2746 => x"0c",
          2747 => x"98",
          2748 => x"0b",
          2749 => x"9c",
          2750 => x"71",
          2751 => x"0c",
          2752 => x"04",
          2753 => x"7f",
          2754 => x"98",
          2755 => x"7d",
          2756 => x"98",
          2757 => x"7d",
          2758 => x"c0",
          2759 => x"5a",
          2760 => x"34",
          2761 => x"b4",
          2762 => x"83",
          2763 => x"c0",
          2764 => x"5a",
          2765 => x"34",
          2766 => x"ac",
          2767 => x"85",
          2768 => x"c0",
          2769 => x"5a",
          2770 => x"34",
          2771 => x"a4",
          2772 => x"88",
          2773 => x"c0",
          2774 => x"5a",
          2775 => x"23",
          2776 => x"79",
          2777 => x"06",
          2778 => x"ff",
          2779 => x"86",
          2780 => x"85",
          2781 => x"84",
          2782 => x"83",
          2783 => x"82",
          2784 => x"7d",
          2785 => x"06",
          2786 => x"e8",
          2787 => x"3f",
          2788 => x"04",
          2789 => x"02",
          2790 => x"70",
          2791 => x"2a",
          2792 => x"70",
          2793 => x"8d",
          2794 => x"3d",
          2795 => x"3d",
          2796 => x"0b",
          2797 => x"33",
          2798 => x"06",
          2799 => x"87",
          2800 => x"51",
          2801 => x"86",
          2802 => x"94",
          2803 => x"08",
          2804 => x"70",
          2805 => x"54",
          2806 => x"2e",
          2807 => x"91",
          2808 => x"06",
          2809 => x"d7",
          2810 => x"32",
          2811 => x"51",
          2812 => x"2e",
          2813 => x"93",
          2814 => x"06",
          2815 => x"ff",
          2816 => x"81",
          2817 => x"87",
          2818 => x"52",
          2819 => x"86",
          2820 => x"94",
          2821 => x"72",
          2822 => x"93",
          2823 => x"3d",
          2824 => x"3d",
          2825 => x"05",
          2826 => x"82",
          2827 => x"70",
          2828 => x"57",
          2829 => x"c0",
          2830 => x"74",
          2831 => x"38",
          2832 => x"94",
          2833 => x"70",
          2834 => x"81",
          2835 => x"52",
          2836 => x"8c",
          2837 => x"2a",
          2838 => x"51",
          2839 => x"38",
          2840 => x"70",
          2841 => x"51",
          2842 => x"8d",
          2843 => x"2a",
          2844 => x"51",
          2845 => x"be",
          2846 => x"ff",
          2847 => x"c0",
          2848 => x"70",
          2849 => x"38",
          2850 => x"90",
          2851 => x"0c",
          2852 => x"04",
          2853 => x"79",
          2854 => x"33",
          2855 => x"06",
          2856 => x"70",
          2857 => x"fe",
          2858 => x"ff",
          2859 => x"0b",
          2860 => x"fc",
          2861 => x"ff",
          2862 => x"55",
          2863 => x"94",
          2864 => x"80",
          2865 => x"87",
          2866 => x"51",
          2867 => x"96",
          2868 => x"06",
          2869 => x"70",
          2870 => x"38",
          2871 => x"70",
          2872 => x"51",
          2873 => x"72",
          2874 => x"81",
          2875 => x"70",
          2876 => x"38",
          2877 => x"70",
          2878 => x"51",
          2879 => x"38",
          2880 => x"06",
          2881 => x"94",
          2882 => x"80",
          2883 => x"87",
          2884 => x"52",
          2885 => x"81",
          2886 => x"70",
          2887 => x"53",
          2888 => x"ff",
          2889 => x"82",
          2890 => x"89",
          2891 => x"fe",
          2892 => x"0b",
          2893 => x"33",
          2894 => x"06",
          2895 => x"c0",
          2896 => x"72",
          2897 => x"38",
          2898 => x"94",
          2899 => x"70",
          2900 => x"81",
          2901 => x"51",
          2902 => x"e2",
          2903 => x"ff",
          2904 => x"c0",
          2905 => x"70",
          2906 => x"38",
          2907 => x"90",
          2908 => x"70",
          2909 => x"82",
          2910 => x"51",
          2911 => x"04",
          2912 => x"0b",
          2913 => x"fc",
          2914 => x"ff",
          2915 => x"87",
          2916 => x"52",
          2917 => x"86",
          2918 => x"94",
          2919 => x"08",
          2920 => x"70",
          2921 => x"51",
          2922 => x"70",
          2923 => x"38",
          2924 => x"06",
          2925 => x"94",
          2926 => x"80",
          2927 => x"87",
          2928 => x"52",
          2929 => x"98",
          2930 => x"2c",
          2931 => x"71",
          2932 => x"0c",
          2933 => x"04",
          2934 => x"87",
          2935 => x"08",
          2936 => x"8a",
          2937 => x"70",
          2938 => x"b4",
          2939 => x"9e",
          2940 => x"8e",
          2941 => x"c0",
          2942 => x"82",
          2943 => x"87",
          2944 => x"08",
          2945 => x"0c",
          2946 => x"98",
          2947 => x"8c",
          2948 => x"9e",
          2949 => x"8e",
          2950 => x"c0",
          2951 => x"82",
          2952 => x"87",
          2953 => x"08",
          2954 => x"0c",
          2955 => x"b0",
          2956 => x"9c",
          2957 => x"9e",
          2958 => x"8e",
          2959 => x"c0",
          2960 => x"82",
          2961 => x"87",
          2962 => x"08",
          2963 => x"0c",
          2964 => x"c0",
          2965 => x"ac",
          2966 => x"9e",
          2967 => x"8e",
          2968 => x"c0",
          2969 => x"51",
          2970 => x"b4",
          2971 => x"9e",
          2972 => x"8e",
          2973 => x"c0",
          2974 => x"82",
          2975 => x"87",
          2976 => x"08",
          2977 => x"0c",
          2978 => x"8e",
          2979 => x"0b",
          2980 => x"90",
          2981 => x"80",
          2982 => x"52",
          2983 => x"2e",
          2984 => x"52",
          2985 => x"c5",
          2986 => x"87",
          2987 => x"08",
          2988 => x"0a",
          2989 => x"52",
          2990 => x"83",
          2991 => x"71",
          2992 => x"34",
          2993 => x"c0",
          2994 => x"70",
          2995 => x"06",
          2996 => x"70",
          2997 => x"38",
          2998 => x"82",
          2999 => x"80",
          3000 => x"9e",
          3001 => x"88",
          3002 => x"51",
          3003 => x"80",
          3004 => x"81",
          3005 => x"8e",
          3006 => x"0b",
          3007 => x"90",
          3008 => x"80",
          3009 => x"52",
          3010 => x"2e",
          3011 => x"52",
          3012 => x"c9",
          3013 => x"87",
          3014 => x"08",
          3015 => x"80",
          3016 => x"52",
          3017 => x"83",
          3018 => x"71",
          3019 => x"34",
          3020 => x"c0",
          3021 => x"70",
          3022 => x"06",
          3023 => x"70",
          3024 => x"38",
          3025 => x"82",
          3026 => x"80",
          3027 => x"9e",
          3028 => x"82",
          3029 => x"51",
          3030 => x"80",
          3031 => x"81",
          3032 => x"8e",
          3033 => x"0b",
          3034 => x"90",
          3035 => x"80",
          3036 => x"52",
          3037 => x"2e",
          3038 => x"52",
          3039 => x"cd",
          3040 => x"87",
          3041 => x"08",
          3042 => x"80",
          3043 => x"52",
          3044 => x"83",
          3045 => x"71",
          3046 => x"34",
          3047 => x"c0",
          3048 => x"70",
          3049 => x"51",
          3050 => x"80",
          3051 => x"81",
          3052 => x"8e",
          3053 => x"c0",
          3054 => x"70",
          3055 => x"70",
          3056 => x"51",
          3057 => x"8e",
          3058 => x"0b",
          3059 => x"90",
          3060 => x"80",
          3061 => x"52",
          3062 => x"83",
          3063 => x"71",
          3064 => x"34",
          3065 => x"90",
          3066 => x"f0",
          3067 => x"2a",
          3068 => x"70",
          3069 => x"34",
          3070 => x"c0",
          3071 => x"70",
          3072 => x"52",
          3073 => x"2e",
          3074 => x"52",
          3075 => x"d3",
          3076 => x"9e",
          3077 => x"87",
          3078 => x"70",
          3079 => x"34",
          3080 => x"04",
          3081 => x"81",
          3082 => x"8a",
          3083 => x"8e",
          3084 => x"73",
          3085 => x"38",
          3086 => x"51",
          3087 => x"81",
          3088 => x"8a",
          3089 => x"8e",
          3090 => x"73",
          3091 => x"38",
          3092 => x"08",
          3093 => x"08",
          3094 => x"81",
          3095 => x"8f",
          3096 => x"8e",
          3097 => x"73",
          3098 => x"38",
          3099 => x"08",
          3100 => x"08",
          3101 => x"81",
          3102 => x"8f",
          3103 => x"8e",
          3104 => x"73",
          3105 => x"38",
          3106 => x"08",
          3107 => x"08",
          3108 => x"81",
          3109 => x"8f",
          3110 => x"8e",
          3111 => x"73",
          3112 => x"38",
          3113 => x"08",
          3114 => x"08",
          3115 => x"81",
          3116 => x"8e",
          3117 => x"8e",
          3118 => x"73",
          3119 => x"38",
          3120 => x"08",
          3121 => x"08",
          3122 => x"81",
          3123 => x"8e",
          3124 => x"8e",
          3125 => x"73",
          3126 => x"38",
          3127 => x"33",
          3128 => x"cc",
          3129 => x"3f",
          3130 => x"33",
          3131 => x"2e",
          3132 => x"8e",
          3133 => x"81",
          3134 => x"8e",
          3135 => x"8e",
          3136 => x"73",
          3137 => x"38",
          3138 => x"33",
          3139 => x"8c",
          3140 => x"3f",
          3141 => x"33",
          3142 => x"2e",
          3143 => x"f9",
          3144 => x"a6",
          3145 => x"c7",
          3146 => x"80",
          3147 => x"81",
          3148 => x"88",
          3149 => x"8e",
          3150 => x"73",
          3151 => x"38",
          3152 => x"51",
          3153 => x"82",
          3154 => x"54",
          3155 => x"88",
          3156 => x"d8",
          3157 => x"3f",
          3158 => x"33",
          3159 => x"2e",
          3160 => x"f9",
          3161 => x"e2",
          3162 => x"f0",
          3163 => x"3f",
          3164 => x"08",
          3165 => x"fc",
          3166 => x"3f",
          3167 => x"08",
          3168 => x"a4",
          3169 => x"3f",
          3170 => x"08",
          3171 => x"cc",
          3172 => x"3f",
          3173 => x"51",
          3174 => x"82",
          3175 => x"52",
          3176 => x"51",
          3177 => x"82",
          3178 => x"56",
          3179 => x"52",
          3180 => x"a9",
          3181 => x"84",
          3182 => x"c0",
          3183 => x"31",
          3184 => x"93",
          3185 => x"81",
          3186 => x"8c",
          3187 => x"8e",
          3188 => x"73",
          3189 => x"38",
          3190 => x"08",
          3191 => x"c0",
          3192 => x"e6",
          3193 => x"93",
          3194 => x"84",
          3195 => x"71",
          3196 => x"82",
          3197 => x"52",
          3198 => x"51",
          3199 => x"82",
          3200 => x"54",
          3201 => x"a8",
          3202 => x"c0",
          3203 => x"84",
          3204 => x"51",
          3205 => x"82",
          3206 => x"bd",
          3207 => x"76",
          3208 => x"54",
          3209 => x"08",
          3210 => x"fc",
          3211 => x"3f",
          3212 => x"51",
          3213 => x"87",
          3214 => x"fe",
          3215 => x"92",
          3216 => x"05",
          3217 => x"26",
          3218 => x"84",
          3219 => x"81",
          3220 => x"52",
          3221 => x"81",
          3222 => x"9d",
          3223 => x"b0",
          3224 => x"81",
          3225 => x"91",
          3226 => x"c0",
          3227 => x"81",
          3228 => x"85",
          3229 => x"cc",
          3230 => x"3f",
          3231 => x"04",
          3232 => x"0c",
          3233 => x"0d",
          3234 => x"84",
          3235 => x"52",
          3236 => x"70",
          3237 => x"82",
          3238 => x"72",
          3239 => x"0d",
          3240 => x"0d",
          3241 => x"84",
          3242 => x"8e",
          3243 => x"80",
          3244 => x"09",
          3245 => x"d8",
          3246 => x"82",
          3247 => x"73",
          3248 => x"3d",
          3249 => x"0b",
          3250 => x"84",
          3251 => x"8e",
          3252 => x"c0",
          3253 => x"04",
          3254 => x"82",
          3255 => x"89",
          3256 => x"c4",
          3257 => x"94",
          3258 => x"94",
          3259 => x"52",
          3260 => x"70",
          3261 => x"26",
          3262 => x"82",
          3263 => x"71",
          3264 => x"93",
          3265 => x"3d",
          3266 => x"3d",
          3267 => x"84",
          3268 => x"12",
          3269 => x"94",
          3270 => x"16",
          3271 => x"54",
          3272 => x"70",
          3273 => x"38",
          3274 => x"14",
          3275 => x"81",
          3276 => x"76",
          3277 => x"0c",
          3278 => x"75",
          3279 => x"72",
          3280 => x"71",
          3281 => x"70",
          3282 => x"70",
          3283 => x"73",
          3284 => x"74",
          3285 => x"70",
          3286 => x"70",
          3287 => x"8c",
          3288 => x"0c",
          3289 => x"0c",
          3290 => x"0c",
          3291 => x"84",
          3292 => x"0d",
          3293 => x"0d",
          3294 => x"08",
          3295 => x"56",
          3296 => x"08",
          3297 => x"81",
          3298 => x"84",
          3299 => x"13",
          3300 => x"73",
          3301 => x"06",
          3302 => x"13",
          3303 => x"13",
          3304 => x"13",
          3305 => x"15",
          3306 => x"9f",
          3307 => x"0c",
          3308 => x"08",
          3309 => x"82",
          3310 => x"94",
          3311 => x"82",
          3312 => x"90",
          3313 => x"94",
          3314 => x"73",
          3315 => x"09",
          3316 => x"38",
          3317 => x"70",
          3318 => x"70",
          3319 => x"81",
          3320 => x"84",
          3321 => x"84",
          3322 => x"14",
          3323 => x"08",
          3324 => x"0c",
          3325 => x"0c",
          3326 => x"88",
          3327 => x"88",
          3328 => x"8c",
          3329 => x"82",
          3330 => x"86",
          3331 => x"f9",
          3332 => x"70",
          3333 => x"80",
          3334 => x"38",
          3335 => x"06",
          3336 => x"08",
          3337 => x"08",
          3338 => x"38",
          3339 => x"77",
          3340 => x"38",
          3341 => x"56",
          3342 => x"ff",
          3343 => x"80",
          3344 => x"52",
          3345 => x"3f",
          3346 => x"08",
          3347 => x"08",
          3348 => x"93",
          3349 => x"80",
          3350 => x"84",
          3351 => x"30",
          3352 => x"80",
          3353 => x"53",
          3354 => x"54",
          3355 => x"72",
          3356 => x"81",
          3357 => x"38",
          3358 => x"52",
          3359 => x"c8",
          3360 => x"82",
          3361 => x"0c",
          3362 => x"84",
          3363 => x"0c",
          3364 => x"08",
          3365 => x"82",
          3366 => x"75",
          3367 => x"38",
          3368 => x"53",
          3369 => x"13",
          3370 => x"0c",
          3371 => x"0c",
          3372 => x"0c",
          3373 => x"76",
          3374 => x"53",
          3375 => x"b5",
          3376 => x"82",
          3377 => x"51",
          3378 => x"82",
          3379 => x"54",
          3380 => x"84",
          3381 => x"0d",
          3382 => x"0d",
          3383 => x"80",
          3384 => x"f0",
          3385 => x"8d",
          3386 => x"0d",
          3387 => x"0d",
          3388 => x"33",
          3389 => x"2e",
          3390 => x"85",
          3391 => x"ed",
          3392 => x"a0",
          3393 => x"80",
          3394 => x"72",
          3395 => x"93",
          3396 => x"05",
          3397 => x"0c",
          3398 => x"93",
          3399 => x"71",
          3400 => x"38",
          3401 => x"2d",
          3402 => x"04",
          3403 => x"02",
          3404 => x"82",
          3405 => x"76",
          3406 => x"0c",
          3407 => x"ad",
          3408 => x"93",
          3409 => x"3d",
          3410 => x"3d",
          3411 => x"73",
          3412 => x"ff",
          3413 => x"71",
          3414 => x"38",
          3415 => x"06",
          3416 => x"54",
          3417 => x"e7",
          3418 => x"0d",
          3419 => x"0d",
          3420 => x"98",
          3421 => x"93",
          3422 => x"54",
          3423 => x"81",
          3424 => x"53",
          3425 => x"8e",
          3426 => x"ff",
          3427 => x"14",
          3428 => x"3f",
          3429 => x"82",
          3430 => x"86",
          3431 => x"ec",
          3432 => x"68",
          3433 => x"70",
          3434 => x"33",
          3435 => x"2e",
          3436 => x"75",
          3437 => x"81",
          3438 => x"38",
          3439 => x"70",
          3440 => x"33",
          3441 => x"75",
          3442 => x"81",
          3443 => x"81",
          3444 => x"75",
          3445 => x"81",
          3446 => x"82",
          3447 => x"81",
          3448 => x"56",
          3449 => x"09",
          3450 => x"38",
          3451 => x"71",
          3452 => x"81",
          3453 => x"59",
          3454 => x"9d",
          3455 => x"53",
          3456 => x"95",
          3457 => x"29",
          3458 => x"76",
          3459 => x"79",
          3460 => x"5b",
          3461 => x"e5",
          3462 => x"ec",
          3463 => x"70",
          3464 => x"25",
          3465 => x"32",
          3466 => x"72",
          3467 => x"73",
          3468 => x"58",
          3469 => x"73",
          3470 => x"38",
          3471 => x"79",
          3472 => x"5b",
          3473 => x"75",
          3474 => x"de",
          3475 => x"80",
          3476 => x"89",
          3477 => x"70",
          3478 => x"55",
          3479 => x"cf",
          3480 => x"38",
          3481 => x"24",
          3482 => x"80",
          3483 => x"8e",
          3484 => x"c3",
          3485 => x"73",
          3486 => x"81",
          3487 => x"99",
          3488 => x"c4",
          3489 => x"38",
          3490 => x"73",
          3491 => x"81",
          3492 => x"80",
          3493 => x"38",
          3494 => x"2e",
          3495 => x"f9",
          3496 => x"d8",
          3497 => x"38",
          3498 => x"77",
          3499 => x"08",
          3500 => x"80",
          3501 => x"55",
          3502 => x"8d",
          3503 => x"70",
          3504 => x"51",
          3505 => x"f5",
          3506 => x"2a",
          3507 => x"74",
          3508 => x"53",
          3509 => x"8f",
          3510 => x"fc",
          3511 => x"81",
          3512 => x"80",
          3513 => x"73",
          3514 => x"3f",
          3515 => x"56",
          3516 => x"27",
          3517 => x"a0",
          3518 => x"3f",
          3519 => x"84",
          3520 => x"33",
          3521 => x"93",
          3522 => x"95",
          3523 => x"91",
          3524 => x"8d",
          3525 => x"89",
          3526 => x"fb",
          3527 => x"86",
          3528 => x"2a",
          3529 => x"51",
          3530 => x"2e",
          3531 => x"84",
          3532 => x"86",
          3533 => x"78",
          3534 => x"08",
          3535 => x"32",
          3536 => x"72",
          3537 => x"51",
          3538 => x"74",
          3539 => x"38",
          3540 => x"88",
          3541 => x"7a",
          3542 => x"55",
          3543 => x"3d",
          3544 => x"52",
          3545 => x"a8",
          3546 => x"84",
          3547 => x"06",
          3548 => x"52",
          3549 => x"3f",
          3550 => x"08",
          3551 => x"27",
          3552 => x"14",
          3553 => x"f8",
          3554 => x"87",
          3555 => x"81",
          3556 => x"b0",
          3557 => x"7d",
          3558 => x"5f",
          3559 => x"75",
          3560 => x"07",
          3561 => x"54",
          3562 => x"26",
          3563 => x"ff",
          3564 => x"84",
          3565 => x"06",
          3566 => x"80",
          3567 => x"96",
          3568 => x"e0",
          3569 => x"73",
          3570 => x"57",
          3571 => x"06",
          3572 => x"54",
          3573 => x"a0",
          3574 => x"2a",
          3575 => x"54",
          3576 => x"38",
          3577 => x"76",
          3578 => x"38",
          3579 => x"fd",
          3580 => x"06",
          3581 => x"38",
          3582 => x"56",
          3583 => x"26",
          3584 => x"3d",
          3585 => x"05",
          3586 => x"ff",
          3587 => x"53",
          3588 => x"d9",
          3589 => x"38",
          3590 => x"56",
          3591 => x"27",
          3592 => x"a0",
          3593 => x"3f",
          3594 => x"3d",
          3595 => x"3d",
          3596 => x"70",
          3597 => x"52",
          3598 => x"73",
          3599 => x"3f",
          3600 => x"04",
          3601 => x"74",
          3602 => x"0c",
          3603 => x"05",
          3604 => x"fa",
          3605 => x"93",
          3606 => x"80",
          3607 => x"0b",
          3608 => x"0c",
          3609 => x"04",
          3610 => x"82",
          3611 => x"76",
          3612 => x"0c",
          3613 => x"05",
          3614 => x"53",
          3615 => x"72",
          3616 => x"0c",
          3617 => x"04",
          3618 => x"77",
          3619 => x"9c",
          3620 => x"54",
          3621 => x"54",
          3622 => x"80",
          3623 => x"93",
          3624 => x"71",
          3625 => x"84",
          3626 => x"06",
          3627 => x"2e",
          3628 => x"72",
          3629 => x"38",
          3630 => x"70",
          3631 => x"25",
          3632 => x"73",
          3633 => x"38",
          3634 => x"86",
          3635 => x"54",
          3636 => x"73",
          3637 => x"ff",
          3638 => x"72",
          3639 => x"74",
          3640 => x"72",
          3641 => x"54",
          3642 => x"81",
          3643 => x"39",
          3644 => x"80",
          3645 => x"51",
          3646 => x"81",
          3647 => x"93",
          3648 => x"3d",
          3649 => x"3d",
          3650 => x"9c",
          3651 => x"93",
          3652 => x"53",
          3653 => x"fe",
          3654 => x"82",
          3655 => x"84",
          3656 => x"f8",
          3657 => x"7c",
          3658 => x"70",
          3659 => x"75",
          3660 => x"55",
          3661 => x"2e",
          3662 => x"87",
          3663 => x"76",
          3664 => x"73",
          3665 => x"81",
          3666 => x"81",
          3667 => x"77",
          3668 => x"70",
          3669 => x"58",
          3670 => x"09",
          3671 => x"c2",
          3672 => x"81",
          3673 => x"75",
          3674 => x"55",
          3675 => x"e2",
          3676 => x"90",
          3677 => x"f8",
          3678 => x"8f",
          3679 => x"81",
          3680 => x"75",
          3681 => x"55",
          3682 => x"81",
          3683 => x"27",
          3684 => x"d0",
          3685 => x"55",
          3686 => x"73",
          3687 => x"80",
          3688 => x"14",
          3689 => x"72",
          3690 => x"e0",
          3691 => x"80",
          3692 => x"39",
          3693 => x"55",
          3694 => x"80",
          3695 => x"e0",
          3696 => x"38",
          3697 => x"81",
          3698 => x"53",
          3699 => x"81",
          3700 => x"53",
          3701 => x"8e",
          3702 => x"70",
          3703 => x"55",
          3704 => x"27",
          3705 => x"77",
          3706 => x"74",
          3707 => x"76",
          3708 => x"77",
          3709 => x"70",
          3710 => x"55",
          3711 => x"77",
          3712 => x"38",
          3713 => x"74",
          3714 => x"55",
          3715 => x"84",
          3716 => x"0d",
          3717 => x"0d",
          3718 => x"56",
          3719 => x"0c",
          3720 => x"70",
          3721 => x"73",
          3722 => x"81",
          3723 => x"81",
          3724 => x"ed",
          3725 => x"2e",
          3726 => x"8e",
          3727 => x"08",
          3728 => x"76",
          3729 => x"56",
          3730 => x"b0",
          3731 => x"06",
          3732 => x"75",
          3733 => x"76",
          3734 => x"70",
          3735 => x"73",
          3736 => x"8b",
          3737 => x"73",
          3738 => x"85",
          3739 => x"82",
          3740 => x"76",
          3741 => x"70",
          3742 => x"ac",
          3743 => x"a0",
          3744 => x"fa",
          3745 => x"53",
          3746 => x"57",
          3747 => x"98",
          3748 => x"39",
          3749 => x"80",
          3750 => x"26",
          3751 => x"86",
          3752 => x"80",
          3753 => x"57",
          3754 => x"74",
          3755 => x"38",
          3756 => x"27",
          3757 => x"14",
          3758 => x"06",
          3759 => x"14",
          3760 => x"06",
          3761 => x"74",
          3762 => x"f9",
          3763 => x"ff",
          3764 => x"89",
          3765 => x"38",
          3766 => x"c5",
          3767 => x"29",
          3768 => x"81",
          3769 => x"76",
          3770 => x"56",
          3771 => x"ba",
          3772 => x"2e",
          3773 => x"30",
          3774 => x"0c",
          3775 => x"82",
          3776 => x"8a",
          3777 => x"fd",
          3778 => x"98",
          3779 => x"2c",
          3780 => x"70",
          3781 => x"10",
          3782 => x"2b",
          3783 => x"54",
          3784 => x"0b",
          3785 => x"12",
          3786 => x"71",
          3787 => x"38",
          3788 => x"11",
          3789 => x"84",
          3790 => x"33",
          3791 => x"52",
          3792 => x"2e",
          3793 => x"83",
          3794 => x"72",
          3795 => x"0c",
          3796 => x"04",
          3797 => x"78",
          3798 => x"9f",
          3799 => x"33",
          3800 => x"71",
          3801 => x"38",
          3802 => x"81",
          3803 => x"f2",
          3804 => x"51",
          3805 => x"72",
          3806 => x"52",
          3807 => x"71",
          3808 => x"52",
          3809 => x"51",
          3810 => x"73",
          3811 => x"3d",
          3812 => x"3d",
          3813 => x"84",
          3814 => x"33",
          3815 => x"bb",
          3816 => x"8f",
          3817 => x"84",
          3818 => x"f8",
          3819 => x"51",
          3820 => x"58",
          3821 => x"2e",
          3822 => x"51",
          3823 => x"82",
          3824 => x"70",
          3825 => x"8e",
          3826 => x"19",
          3827 => x"56",
          3828 => x"3f",
          3829 => x"08",
          3830 => x"8f",
          3831 => x"84",
          3832 => x"f8",
          3833 => x"51",
          3834 => x"80",
          3835 => x"75",
          3836 => x"74",
          3837 => x"3f",
          3838 => x"33",
          3839 => x"74",
          3840 => x"34",
          3841 => x"06",
          3842 => x"27",
          3843 => x"0b",
          3844 => x"34",
          3845 => x"b6",
          3846 => x"cc",
          3847 => x"80",
          3848 => x"82",
          3849 => x"55",
          3850 => x"8c",
          3851 => x"54",
          3852 => x"52",
          3853 => x"c8",
          3854 => x"8f",
          3855 => x"8a",
          3856 => x"9e",
          3857 => x"cc",
          3858 => x"cb",
          3859 => x"3d",
          3860 => x"3d",
          3861 => x"80",
          3862 => x"cc",
          3863 => x"d2",
          3864 => x"93",
          3865 => x"d1",
          3866 => x"cc",
          3867 => x"f8",
          3868 => x"70",
          3869 => x"fa",
          3870 => x"93",
          3871 => x"2e",
          3872 => x"51",
          3873 => x"82",
          3874 => x"55",
          3875 => x"93",
          3876 => x"9c",
          3877 => x"84",
          3878 => x"70",
          3879 => x"80",
          3880 => x"53",
          3881 => x"17",
          3882 => x"52",
          3883 => x"3f",
          3884 => x"09",
          3885 => x"b1",
          3886 => x"0d",
          3887 => x"0d",
          3888 => x"ad",
          3889 => x"5a",
          3890 => x"58",
          3891 => x"8f",
          3892 => x"80",
          3893 => x"82",
          3894 => x"81",
          3895 => x"0b",
          3896 => x"08",
          3897 => x"f8",
          3898 => x"70",
          3899 => x"f9",
          3900 => x"93",
          3901 => x"2e",
          3902 => x"51",
          3903 => x"82",
          3904 => x"81",
          3905 => x"80",
          3906 => x"84",
          3907 => x"38",
          3908 => x"08",
          3909 => x"17",
          3910 => x"74",
          3911 => x"70",
          3912 => x"07",
          3913 => x"55",
          3914 => x"2e",
          3915 => x"ff",
          3916 => x"8f",
          3917 => x"11",
          3918 => x"80",
          3919 => x"82",
          3920 => x"80",
          3921 => x"81",
          3922 => x"ef",
          3923 => x"77",
          3924 => x"06",
          3925 => x"52",
          3926 => x"a5",
          3927 => x"d6",
          3928 => x"3d",
          3929 => x"93",
          3930 => x"34",
          3931 => x"82",
          3932 => x"a9",
          3933 => x"f6",
          3934 => x"7e",
          3935 => x"72",
          3936 => x"5a",
          3937 => x"2e",
          3938 => x"a2",
          3939 => x"78",
          3940 => x"76",
          3941 => x"81",
          3942 => x"70",
          3943 => x"58",
          3944 => x"2e",
          3945 => x"86",
          3946 => x"26",
          3947 => x"54",
          3948 => x"82",
          3949 => x"70",
          3950 => x"d5",
          3951 => x"93",
          3952 => x"79",
          3953 => x"51",
          3954 => x"82",
          3955 => x"80",
          3956 => x"15",
          3957 => x"81",
          3958 => x"74",
          3959 => x"38",
          3960 => x"ee",
          3961 => x"81",
          3962 => x"3d",
          3963 => x"f8",
          3964 => x"af",
          3965 => x"84",
          3966 => x"99",
          3967 => x"78",
          3968 => x"fd",
          3969 => x"93",
          3970 => x"ff",
          3971 => x"85",
          3972 => x"91",
          3973 => x"70",
          3974 => x"51",
          3975 => x"27",
          3976 => x"80",
          3977 => x"93",
          3978 => x"3d",
          3979 => x"3d",
          3980 => x"08",
          3981 => x"81",
          3982 => x"5f",
          3983 => x"af",
          3984 => x"8f",
          3985 => x"82",
          3986 => x"81",
          3987 => x"8f",
          3988 => x"73",
          3989 => x"a8",
          3990 => x"3f",
          3991 => x"08",
          3992 => x"0c",
          3993 => x"08",
          3994 => x"fe",
          3995 => x"82",
          3996 => x"52",
          3997 => x"08",
          3998 => x"3f",
          3999 => x"08",
          4000 => x"38",
          4001 => x"51",
          4002 => x"80",
          4003 => x"8f",
          4004 => x"80",
          4005 => x"3d",
          4006 => x"80",
          4007 => x"82",
          4008 => x"56",
          4009 => x"08",
          4010 => x"81",
          4011 => x"38",
          4012 => x"08",
          4013 => x"3f",
          4014 => x"08",
          4015 => x"82",
          4016 => x"25",
          4017 => x"93",
          4018 => x"05",
          4019 => x"55",
          4020 => x"80",
          4021 => x"ff",
          4022 => x"51",
          4023 => x"74",
          4024 => x"81",
          4025 => x"38",
          4026 => x"0b",
          4027 => x"34",
          4028 => x"dd",
          4029 => x"93",
          4030 => x"2b",
          4031 => x"51",
          4032 => x"2e",
          4033 => x"81",
          4034 => x"93",
          4035 => x"98",
          4036 => x"2c",
          4037 => x"33",
          4038 => x"70",
          4039 => x"98",
          4040 => x"84",
          4041 => x"dc",
          4042 => x"15",
          4043 => x"51",
          4044 => x"59",
          4045 => x"58",
          4046 => x"78",
          4047 => x"38",
          4048 => x"b4",
          4049 => x"80",
          4050 => x"ff",
          4051 => x"98",
          4052 => x"80",
          4053 => x"ce",
          4054 => x"74",
          4055 => x"f7",
          4056 => x"93",
          4057 => x"ff",
          4058 => x"80",
          4059 => x"74",
          4060 => x"34",
          4061 => x"39",
          4062 => x"0a",
          4063 => x"0a",
          4064 => x"2c",
          4065 => x"06",
          4066 => x"73",
          4067 => x"38",
          4068 => x"52",
          4069 => x"ef",
          4070 => x"84",
          4071 => x"06",
          4072 => x"38",
          4073 => x"56",
          4074 => x"80",
          4075 => x"1c",
          4076 => x"93",
          4077 => x"98",
          4078 => x"2c",
          4079 => x"33",
          4080 => x"70",
          4081 => x"10",
          4082 => x"2b",
          4083 => x"11",
          4084 => x"51",
          4085 => x"51",
          4086 => x"2e",
          4087 => x"fe",
          4088 => x"fd",
          4089 => x"7d",
          4090 => x"82",
          4091 => x"80",
          4092 => x"a4",
          4093 => x"75",
          4094 => x"34",
          4095 => x"a4",
          4096 => x"3d",
          4097 => x"0c",
          4098 => x"8b",
          4099 => x"38",
          4100 => x"81",
          4101 => x"54",
          4102 => x"82",
          4103 => x"54",
          4104 => x"fd",
          4105 => x"93",
          4106 => x"73",
          4107 => x"38",
          4108 => x"70",
          4109 => x"55",
          4110 => x"9e",
          4111 => x"54",
          4112 => x"15",
          4113 => x"80",
          4114 => x"ff",
          4115 => x"98",
          4116 => x"b0",
          4117 => x"55",
          4118 => x"93",
          4119 => x"11",
          4120 => x"82",
          4121 => x"73",
          4122 => x"3d",
          4123 => x"82",
          4124 => x"54",
          4125 => x"89",
          4126 => x"54",
          4127 => x"ac",
          4128 => x"b0",
          4129 => x"80",
          4130 => x"ff",
          4131 => x"98",
          4132 => x"ac",
          4133 => x"56",
          4134 => x"25",
          4135 => x"1a",
          4136 => x"54",
          4137 => x"74",
          4138 => x"29",
          4139 => x"05",
          4140 => x"82",
          4141 => x"56",
          4142 => x"75",
          4143 => x"82",
          4144 => x"70",
          4145 => x"98",
          4146 => x"ac",
          4147 => x"56",
          4148 => x"25",
          4149 => x"88",
          4150 => x"3f",
          4151 => x"0a",
          4152 => x"0a",
          4153 => x"2c",
          4154 => x"33",
          4155 => x"73",
          4156 => x"38",
          4157 => x"82",
          4158 => x"70",
          4159 => x"55",
          4160 => x"2e",
          4161 => x"82",
          4162 => x"ff",
          4163 => x"82",
          4164 => x"ff",
          4165 => x"82",
          4166 => x"88",
          4167 => x"3f",
          4168 => x"33",
          4169 => x"70",
          4170 => x"93",
          4171 => x"51",
          4172 => x"74",
          4173 => x"74",
          4174 => x"14",
          4175 => x"73",
          4176 => x"a9",
          4177 => x"80",
          4178 => x"80",
          4179 => x"98",
          4180 => x"ac",
          4181 => x"55",
          4182 => x"db",
          4183 => x"e7",
          4184 => x"93",
          4185 => x"98",
          4186 => x"2c",
          4187 => x"33",
          4188 => x"57",
          4189 => x"fa",
          4190 => x"51",
          4191 => x"74",
          4192 => x"29",
          4193 => x"05",
          4194 => x"82",
          4195 => x"58",
          4196 => x"75",
          4197 => x"fa",
          4198 => x"93",
          4199 => x"05",
          4200 => x"34",
          4201 => x"c5",
          4202 => x"ac",
          4203 => x"f7",
          4204 => x"93",
          4205 => x"ff",
          4206 => x"98",
          4207 => x"ac",
          4208 => x"80",
          4209 => x"38",
          4210 => x"52",
          4211 => x"c2",
          4212 => x"39",
          4213 => x"84",
          4214 => x"93",
          4215 => x"73",
          4216 => x"8c",
          4217 => x"e6",
          4218 => x"93",
          4219 => x"05",
          4220 => x"93",
          4221 => x"81",
          4222 => x"e3",
          4223 => x"b0",
          4224 => x"ac",
          4225 => x"73",
          4226 => x"e4",
          4227 => x"54",
          4228 => x"ac",
          4229 => x"2b",
          4230 => x"75",
          4231 => x"56",
          4232 => x"74",
          4233 => x"74",
          4234 => x"14",
          4235 => x"73",
          4236 => x"b9",
          4237 => x"80",
          4238 => x"80",
          4239 => x"98",
          4240 => x"ac",
          4241 => x"55",
          4242 => x"db",
          4243 => x"e5",
          4244 => x"93",
          4245 => x"98",
          4246 => x"2c",
          4247 => x"33",
          4248 => x"57",
          4249 => x"f9",
          4250 => x"51",
          4251 => x"74",
          4252 => x"29",
          4253 => x"05",
          4254 => x"82",
          4255 => x"58",
          4256 => x"75",
          4257 => x"f8",
          4258 => x"93",
          4259 => x"81",
          4260 => x"93",
          4261 => x"56",
          4262 => x"27",
          4263 => x"81",
          4264 => x"82",
          4265 => x"74",
          4266 => x"52",
          4267 => x"3f",
          4268 => x"33",
          4269 => x"06",
          4270 => x"33",
          4271 => x"75",
          4272 => x"38",
          4273 => x"7a",
          4274 => x"8f",
          4275 => x"74",
          4276 => x"38",
          4277 => x"98",
          4278 => x"84",
          4279 => x"ac",
          4280 => x"84",
          4281 => x"06",
          4282 => x"74",
          4283 => x"c7",
          4284 => x"5b",
          4285 => x"7a",
          4286 => x"8e",
          4287 => x"11",
          4288 => x"74",
          4289 => x"38",
          4290 => x"e4",
          4291 => x"84",
          4292 => x"ac",
          4293 => x"84",
          4294 => x"06",
          4295 => x"74",
          4296 => x"c7",
          4297 => x"1b",
          4298 => x"39",
          4299 => x"74",
          4300 => x"bc",
          4301 => x"ca",
          4302 => x"e2",
          4303 => x"2e",
          4304 => x"93",
          4305 => x"f8",
          4306 => x"80",
          4307 => x"74",
          4308 => x"3f",
          4309 => x"7a",
          4310 => x"8e",
          4311 => x"11",
          4312 => x"74",
          4313 => x"38",
          4314 => x"84",
          4315 => x"84",
          4316 => x"ac",
          4317 => x"84",
          4318 => x"06",
          4319 => x"74",
          4320 => x"c6",
          4321 => x"1b",
          4322 => x"ff",
          4323 => x"39",
          4324 => x"74",
          4325 => x"d8",
          4326 => x"c9",
          4327 => x"93",
          4328 => x"93",
          4329 => x"93",
          4330 => x"ff",
          4331 => x"53",
          4332 => x"51",
          4333 => x"82",
          4334 => x"82",
          4335 => x"52",
          4336 => x"90",
          4337 => x"39",
          4338 => x"33",
          4339 => x"06",
          4340 => x"33",
          4341 => x"74",
          4342 => x"94",
          4343 => x"54",
          4344 => x"b0",
          4345 => x"70",
          4346 => x"e2",
          4347 => x"80",
          4348 => x"b0",
          4349 => x"80",
          4350 => x"38",
          4351 => x"ed",
          4352 => x"b0",
          4353 => x"54",
          4354 => x"b0",
          4355 => x"39",
          4356 => x"93",
          4357 => x"0b",
          4358 => x"34",
          4359 => x"84",
          4360 => x"0d",
          4361 => x"0d",
          4362 => x"33",
          4363 => x"70",
          4364 => x"38",
          4365 => x"11",
          4366 => x"82",
          4367 => x"83",
          4368 => x"fc",
          4369 => x"9b",
          4370 => x"84",
          4371 => x"33",
          4372 => x"51",
          4373 => x"80",
          4374 => x"84",
          4375 => x"92",
          4376 => x"51",
          4377 => x"80",
          4378 => x"81",
          4379 => x"72",
          4380 => x"92",
          4381 => x"81",
          4382 => x"0b",
          4383 => x"8c",
          4384 => x"71",
          4385 => x"06",
          4386 => x"80",
          4387 => x"87",
          4388 => x"08",
          4389 => x"38",
          4390 => x"80",
          4391 => x"71",
          4392 => x"c0",
          4393 => x"51",
          4394 => x"87",
          4395 => x"8f",
          4396 => x"82",
          4397 => x"33",
          4398 => x"93",
          4399 => x"3d",
          4400 => x"3d",
          4401 => x"64",
          4402 => x"bf",
          4403 => x"40",
          4404 => x"74",
          4405 => x"cd",
          4406 => x"84",
          4407 => x"7a",
          4408 => x"81",
          4409 => x"72",
          4410 => x"87",
          4411 => x"11",
          4412 => x"8c",
          4413 => x"92",
          4414 => x"5a",
          4415 => x"58",
          4416 => x"c0",
          4417 => x"76",
          4418 => x"76",
          4419 => x"70",
          4420 => x"81",
          4421 => x"54",
          4422 => x"8e",
          4423 => x"52",
          4424 => x"81",
          4425 => x"81",
          4426 => x"74",
          4427 => x"53",
          4428 => x"83",
          4429 => x"78",
          4430 => x"8f",
          4431 => x"2e",
          4432 => x"c0",
          4433 => x"52",
          4434 => x"87",
          4435 => x"08",
          4436 => x"2e",
          4437 => x"84",
          4438 => x"38",
          4439 => x"87",
          4440 => x"15",
          4441 => x"70",
          4442 => x"52",
          4443 => x"ff",
          4444 => x"39",
          4445 => x"81",
          4446 => x"ff",
          4447 => x"57",
          4448 => x"90",
          4449 => x"80",
          4450 => x"71",
          4451 => x"78",
          4452 => x"38",
          4453 => x"80",
          4454 => x"80",
          4455 => x"81",
          4456 => x"72",
          4457 => x"0c",
          4458 => x"04",
          4459 => x"60",
          4460 => x"8c",
          4461 => x"33",
          4462 => x"5b",
          4463 => x"74",
          4464 => x"e1",
          4465 => x"84",
          4466 => x"79",
          4467 => x"78",
          4468 => x"06",
          4469 => x"77",
          4470 => x"87",
          4471 => x"11",
          4472 => x"8c",
          4473 => x"92",
          4474 => x"59",
          4475 => x"85",
          4476 => x"98",
          4477 => x"7d",
          4478 => x"0c",
          4479 => x"08",
          4480 => x"70",
          4481 => x"53",
          4482 => x"2e",
          4483 => x"70",
          4484 => x"33",
          4485 => x"18",
          4486 => x"2a",
          4487 => x"51",
          4488 => x"2e",
          4489 => x"c0",
          4490 => x"52",
          4491 => x"87",
          4492 => x"08",
          4493 => x"2e",
          4494 => x"84",
          4495 => x"38",
          4496 => x"87",
          4497 => x"15",
          4498 => x"70",
          4499 => x"52",
          4500 => x"ff",
          4501 => x"39",
          4502 => x"81",
          4503 => x"80",
          4504 => x"52",
          4505 => x"90",
          4506 => x"80",
          4507 => x"71",
          4508 => x"7a",
          4509 => x"38",
          4510 => x"80",
          4511 => x"80",
          4512 => x"81",
          4513 => x"72",
          4514 => x"0c",
          4515 => x"04",
          4516 => x"7a",
          4517 => x"a3",
          4518 => x"88",
          4519 => x"33",
          4520 => x"56",
          4521 => x"3f",
          4522 => x"08",
          4523 => x"83",
          4524 => x"fe",
          4525 => x"87",
          4526 => x"0c",
          4527 => x"76",
          4528 => x"38",
          4529 => x"93",
          4530 => x"2b",
          4531 => x"8c",
          4532 => x"71",
          4533 => x"38",
          4534 => x"71",
          4535 => x"c6",
          4536 => x"39",
          4537 => x"81",
          4538 => x"06",
          4539 => x"71",
          4540 => x"38",
          4541 => x"8c",
          4542 => x"e8",
          4543 => x"98",
          4544 => x"71",
          4545 => x"73",
          4546 => x"92",
          4547 => x"72",
          4548 => x"06",
          4549 => x"f7",
          4550 => x"80",
          4551 => x"88",
          4552 => x"0c",
          4553 => x"80",
          4554 => x"56",
          4555 => x"56",
          4556 => x"82",
          4557 => x"88",
          4558 => x"fe",
          4559 => x"81",
          4560 => x"33",
          4561 => x"07",
          4562 => x"0c",
          4563 => x"3d",
          4564 => x"3d",
          4565 => x"11",
          4566 => x"33",
          4567 => x"71",
          4568 => x"81",
          4569 => x"72",
          4570 => x"75",
          4571 => x"82",
          4572 => x"52",
          4573 => x"54",
          4574 => x"0d",
          4575 => x"0d",
          4576 => x"05",
          4577 => x"52",
          4578 => x"70",
          4579 => x"34",
          4580 => x"51",
          4581 => x"83",
          4582 => x"ff",
          4583 => x"75",
          4584 => x"72",
          4585 => x"54",
          4586 => x"2a",
          4587 => x"70",
          4588 => x"34",
          4589 => x"51",
          4590 => x"81",
          4591 => x"70",
          4592 => x"70",
          4593 => x"3d",
          4594 => x"3d",
          4595 => x"77",
          4596 => x"70",
          4597 => x"38",
          4598 => x"05",
          4599 => x"70",
          4600 => x"34",
          4601 => x"eb",
          4602 => x"0d",
          4603 => x"0d",
          4604 => x"54",
          4605 => x"72",
          4606 => x"54",
          4607 => x"51",
          4608 => x"84",
          4609 => x"fc",
          4610 => x"77",
          4611 => x"53",
          4612 => x"05",
          4613 => x"70",
          4614 => x"33",
          4615 => x"ff",
          4616 => x"52",
          4617 => x"2e",
          4618 => x"80",
          4619 => x"71",
          4620 => x"0c",
          4621 => x"04",
          4622 => x"74",
          4623 => x"89",
          4624 => x"2e",
          4625 => x"11",
          4626 => x"52",
          4627 => x"70",
          4628 => x"84",
          4629 => x"0d",
          4630 => x"82",
          4631 => x"04",
          4632 => x"93",
          4633 => x"f7",
          4634 => x"56",
          4635 => x"17",
          4636 => x"74",
          4637 => x"d6",
          4638 => x"b0",
          4639 => x"b4",
          4640 => x"81",
          4641 => x"59",
          4642 => x"82",
          4643 => x"7a",
          4644 => x"06",
          4645 => x"93",
          4646 => x"17",
          4647 => x"08",
          4648 => x"08",
          4649 => x"08",
          4650 => x"74",
          4651 => x"38",
          4652 => x"55",
          4653 => x"09",
          4654 => x"38",
          4655 => x"18",
          4656 => x"81",
          4657 => x"f9",
          4658 => x"39",
          4659 => x"82",
          4660 => x"8b",
          4661 => x"fa",
          4662 => x"7a",
          4663 => x"57",
          4664 => x"08",
          4665 => x"75",
          4666 => x"3f",
          4667 => x"08",
          4668 => x"84",
          4669 => x"81",
          4670 => x"b4",
          4671 => x"16",
          4672 => x"be",
          4673 => x"84",
          4674 => x"85",
          4675 => x"81",
          4676 => x"17",
          4677 => x"93",
          4678 => x"3d",
          4679 => x"3d",
          4680 => x"52",
          4681 => x"3f",
          4682 => x"08",
          4683 => x"84",
          4684 => x"38",
          4685 => x"74",
          4686 => x"81",
          4687 => x"38",
          4688 => x"59",
          4689 => x"09",
          4690 => x"e3",
          4691 => x"53",
          4692 => x"08",
          4693 => x"70",
          4694 => x"91",
          4695 => x"d5",
          4696 => x"17",
          4697 => x"3f",
          4698 => x"a4",
          4699 => x"51",
          4700 => x"86",
          4701 => x"f2",
          4702 => x"17",
          4703 => x"3f",
          4704 => x"52",
          4705 => x"51",
          4706 => x"8c",
          4707 => x"84",
          4708 => x"fc",
          4709 => x"17",
          4710 => x"70",
          4711 => x"79",
          4712 => x"52",
          4713 => x"51",
          4714 => x"77",
          4715 => x"80",
          4716 => x"81",
          4717 => x"f9",
          4718 => x"93",
          4719 => x"2e",
          4720 => x"58",
          4721 => x"84",
          4722 => x"0d",
          4723 => x"0d",
          4724 => x"98",
          4725 => x"05",
          4726 => x"80",
          4727 => x"27",
          4728 => x"14",
          4729 => x"29",
          4730 => x"05",
          4731 => x"82",
          4732 => x"87",
          4733 => x"f9",
          4734 => x"7a",
          4735 => x"54",
          4736 => x"27",
          4737 => x"76",
          4738 => x"27",
          4739 => x"ff",
          4740 => x"58",
          4741 => x"80",
          4742 => x"82",
          4743 => x"72",
          4744 => x"38",
          4745 => x"72",
          4746 => x"8e",
          4747 => x"39",
          4748 => x"17",
          4749 => x"a4",
          4750 => x"53",
          4751 => x"fd",
          4752 => x"93",
          4753 => x"9f",
          4754 => x"ff",
          4755 => x"11",
          4756 => x"70",
          4757 => x"18",
          4758 => x"76",
          4759 => x"53",
          4760 => x"82",
          4761 => x"80",
          4762 => x"83",
          4763 => x"b4",
          4764 => x"88",
          4765 => x"79",
          4766 => x"84",
          4767 => x"58",
          4768 => x"80",
          4769 => x"9f",
          4770 => x"80",
          4771 => x"88",
          4772 => x"08",
          4773 => x"51",
          4774 => x"82",
          4775 => x"80",
          4776 => x"10",
          4777 => x"74",
          4778 => x"51",
          4779 => x"82",
          4780 => x"83",
          4781 => x"58",
          4782 => x"87",
          4783 => x"08",
          4784 => x"51",
          4785 => x"82",
          4786 => x"9b",
          4787 => x"2b",
          4788 => x"74",
          4789 => x"51",
          4790 => x"82",
          4791 => x"f0",
          4792 => x"83",
          4793 => x"77",
          4794 => x"0c",
          4795 => x"04",
          4796 => x"7a",
          4797 => x"58",
          4798 => x"81",
          4799 => x"9e",
          4800 => x"17",
          4801 => x"96",
          4802 => x"53",
          4803 => x"81",
          4804 => x"79",
          4805 => x"72",
          4806 => x"38",
          4807 => x"72",
          4808 => x"b8",
          4809 => x"39",
          4810 => x"17",
          4811 => x"a4",
          4812 => x"53",
          4813 => x"fb",
          4814 => x"93",
          4815 => x"82",
          4816 => x"81",
          4817 => x"83",
          4818 => x"b4",
          4819 => x"78",
          4820 => x"56",
          4821 => x"76",
          4822 => x"38",
          4823 => x"9f",
          4824 => x"33",
          4825 => x"07",
          4826 => x"74",
          4827 => x"83",
          4828 => x"89",
          4829 => x"08",
          4830 => x"51",
          4831 => x"82",
          4832 => x"59",
          4833 => x"08",
          4834 => x"74",
          4835 => x"16",
          4836 => x"84",
          4837 => x"76",
          4838 => x"88",
          4839 => x"81",
          4840 => x"8f",
          4841 => x"53",
          4842 => x"80",
          4843 => x"88",
          4844 => x"08",
          4845 => x"51",
          4846 => x"82",
          4847 => x"59",
          4848 => x"08",
          4849 => x"77",
          4850 => x"06",
          4851 => x"83",
          4852 => x"05",
          4853 => x"f7",
          4854 => x"39",
          4855 => x"a4",
          4856 => x"52",
          4857 => x"ef",
          4858 => x"84",
          4859 => x"93",
          4860 => x"38",
          4861 => x"06",
          4862 => x"83",
          4863 => x"18",
          4864 => x"54",
          4865 => x"f6",
          4866 => x"93",
          4867 => x"0a",
          4868 => x"52",
          4869 => x"83",
          4870 => x"83",
          4871 => x"82",
          4872 => x"8a",
          4873 => x"f8",
          4874 => x"7c",
          4875 => x"59",
          4876 => x"81",
          4877 => x"38",
          4878 => x"08",
          4879 => x"73",
          4880 => x"38",
          4881 => x"52",
          4882 => x"a4",
          4883 => x"84",
          4884 => x"93",
          4885 => x"f2",
          4886 => x"82",
          4887 => x"39",
          4888 => x"e6",
          4889 => x"84",
          4890 => x"de",
          4891 => x"78",
          4892 => x"3f",
          4893 => x"08",
          4894 => x"84",
          4895 => x"80",
          4896 => x"93",
          4897 => x"2e",
          4898 => x"93",
          4899 => x"2e",
          4900 => x"53",
          4901 => x"51",
          4902 => x"82",
          4903 => x"c5",
          4904 => x"08",
          4905 => x"18",
          4906 => x"57",
          4907 => x"90",
          4908 => x"90",
          4909 => x"16",
          4910 => x"54",
          4911 => x"34",
          4912 => x"78",
          4913 => x"38",
          4914 => x"82",
          4915 => x"8a",
          4916 => x"f6",
          4917 => x"7e",
          4918 => x"5b",
          4919 => x"38",
          4920 => x"58",
          4921 => x"88",
          4922 => x"08",
          4923 => x"38",
          4924 => x"39",
          4925 => x"51",
          4926 => x"81",
          4927 => x"93",
          4928 => x"82",
          4929 => x"93",
          4930 => x"82",
          4931 => x"ff",
          4932 => x"38",
          4933 => x"82",
          4934 => x"26",
          4935 => x"79",
          4936 => x"08",
          4937 => x"73",
          4938 => x"b9",
          4939 => x"2e",
          4940 => x"80",
          4941 => x"1a",
          4942 => x"08",
          4943 => x"38",
          4944 => x"52",
          4945 => x"af",
          4946 => x"82",
          4947 => x"81",
          4948 => x"06",
          4949 => x"93",
          4950 => x"82",
          4951 => x"09",
          4952 => x"72",
          4953 => x"70",
          4954 => x"93",
          4955 => x"51",
          4956 => x"73",
          4957 => x"82",
          4958 => x"80",
          4959 => x"8c",
          4960 => x"81",
          4961 => x"38",
          4962 => x"08",
          4963 => x"73",
          4964 => x"75",
          4965 => x"77",
          4966 => x"56",
          4967 => x"76",
          4968 => x"82",
          4969 => x"26",
          4970 => x"75",
          4971 => x"f8",
          4972 => x"93",
          4973 => x"2e",
          4974 => x"59",
          4975 => x"08",
          4976 => x"81",
          4977 => x"82",
          4978 => x"59",
          4979 => x"08",
          4980 => x"70",
          4981 => x"25",
          4982 => x"51",
          4983 => x"73",
          4984 => x"75",
          4985 => x"81",
          4986 => x"38",
          4987 => x"f5",
          4988 => x"75",
          4989 => x"f9",
          4990 => x"93",
          4991 => x"93",
          4992 => x"70",
          4993 => x"08",
          4994 => x"51",
          4995 => x"80",
          4996 => x"73",
          4997 => x"38",
          4998 => x"52",
          4999 => x"d0",
          5000 => x"84",
          5001 => x"a5",
          5002 => x"18",
          5003 => x"08",
          5004 => x"18",
          5005 => x"74",
          5006 => x"38",
          5007 => x"18",
          5008 => x"33",
          5009 => x"73",
          5010 => x"97",
          5011 => x"74",
          5012 => x"38",
          5013 => x"55",
          5014 => x"93",
          5015 => x"85",
          5016 => x"75",
          5017 => x"93",
          5018 => x"3d",
          5019 => x"3d",
          5020 => x"52",
          5021 => x"3f",
          5022 => x"08",
          5023 => x"82",
          5024 => x"80",
          5025 => x"52",
          5026 => x"c1",
          5027 => x"84",
          5028 => x"84",
          5029 => x"0c",
          5030 => x"53",
          5031 => x"15",
          5032 => x"f2",
          5033 => x"56",
          5034 => x"16",
          5035 => x"22",
          5036 => x"27",
          5037 => x"54",
          5038 => x"76",
          5039 => x"33",
          5040 => x"3f",
          5041 => x"08",
          5042 => x"38",
          5043 => x"76",
          5044 => x"70",
          5045 => x"9f",
          5046 => x"56",
          5047 => x"93",
          5048 => x"3d",
          5049 => x"3d",
          5050 => x"71",
          5051 => x"57",
          5052 => x"0a",
          5053 => x"38",
          5054 => x"53",
          5055 => x"38",
          5056 => x"0c",
          5057 => x"54",
          5058 => x"75",
          5059 => x"73",
          5060 => x"a8",
          5061 => x"73",
          5062 => x"85",
          5063 => x"0b",
          5064 => x"5a",
          5065 => x"27",
          5066 => x"a8",
          5067 => x"18",
          5068 => x"39",
          5069 => x"70",
          5070 => x"58",
          5071 => x"b2",
          5072 => x"76",
          5073 => x"3f",
          5074 => x"08",
          5075 => x"84",
          5076 => x"bd",
          5077 => x"82",
          5078 => x"27",
          5079 => x"16",
          5080 => x"84",
          5081 => x"38",
          5082 => x"39",
          5083 => x"55",
          5084 => x"52",
          5085 => x"d5",
          5086 => x"84",
          5087 => x"0c",
          5088 => x"0c",
          5089 => x"53",
          5090 => x"80",
          5091 => x"85",
          5092 => x"94",
          5093 => x"2a",
          5094 => x"0c",
          5095 => x"06",
          5096 => x"9c",
          5097 => x"58",
          5098 => x"84",
          5099 => x"0d",
          5100 => x"0d",
          5101 => x"90",
          5102 => x"05",
          5103 => x"f0",
          5104 => x"27",
          5105 => x"0b",
          5106 => x"98",
          5107 => x"84",
          5108 => x"2e",
          5109 => x"76",
          5110 => x"58",
          5111 => x"38",
          5112 => x"15",
          5113 => x"08",
          5114 => x"38",
          5115 => x"88",
          5116 => x"53",
          5117 => x"81",
          5118 => x"c0",
          5119 => x"22",
          5120 => x"89",
          5121 => x"72",
          5122 => x"74",
          5123 => x"f3",
          5124 => x"93",
          5125 => x"82",
          5126 => x"82",
          5127 => x"27",
          5128 => x"81",
          5129 => x"84",
          5130 => x"80",
          5131 => x"16",
          5132 => x"84",
          5133 => x"ca",
          5134 => x"38",
          5135 => x"0c",
          5136 => x"dd",
          5137 => x"08",
          5138 => x"f9",
          5139 => x"93",
          5140 => x"87",
          5141 => x"84",
          5142 => x"80",
          5143 => x"55",
          5144 => x"08",
          5145 => x"38",
          5146 => x"93",
          5147 => x"2e",
          5148 => x"93",
          5149 => x"75",
          5150 => x"3f",
          5151 => x"08",
          5152 => x"94",
          5153 => x"52",
          5154 => x"c1",
          5155 => x"84",
          5156 => x"0c",
          5157 => x"0c",
          5158 => x"05",
          5159 => x"80",
          5160 => x"93",
          5161 => x"3d",
          5162 => x"3d",
          5163 => x"71",
          5164 => x"57",
          5165 => x"51",
          5166 => x"82",
          5167 => x"54",
          5168 => x"08",
          5169 => x"82",
          5170 => x"56",
          5171 => x"52",
          5172 => x"83",
          5173 => x"84",
          5174 => x"93",
          5175 => x"d2",
          5176 => x"84",
          5177 => x"08",
          5178 => x"54",
          5179 => x"e5",
          5180 => x"06",
          5181 => x"58",
          5182 => x"08",
          5183 => x"38",
          5184 => x"75",
          5185 => x"80",
          5186 => x"81",
          5187 => x"7a",
          5188 => x"06",
          5189 => x"39",
          5190 => x"08",
          5191 => x"76",
          5192 => x"3f",
          5193 => x"08",
          5194 => x"84",
          5195 => x"ff",
          5196 => x"84",
          5197 => x"06",
          5198 => x"54",
          5199 => x"84",
          5200 => x"0d",
          5201 => x"0d",
          5202 => x"52",
          5203 => x"3f",
          5204 => x"08",
          5205 => x"06",
          5206 => x"51",
          5207 => x"83",
          5208 => x"06",
          5209 => x"14",
          5210 => x"3f",
          5211 => x"08",
          5212 => x"07",
          5213 => x"93",
          5214 => x"3d",
          5215 => x"3d",
          5216 => x"70",
          5217 => x"06",
          5218 => x"53",
          5219 => x"ed",
          5220 => x"33",
          5221 => x"83",
          5222 => x"06",
          5223 => x"90",
          5224 => x"15",
          5225 => x"3f",
          5226 => x"04",
          5227 => x"7b",
          5228 => x"84",
          5229 => x"58",
          5230 => x"80",
          5231 => x"38",
          5232 => x"52",
          5233 => x"8f",
          5234 => x"84",
          5235 => x"93",
          5236 => x"f5",
          5237 => x"08",
          5238 => x"53",
          5239 => x"84",
          5240 => x"39",
          5241 => x"70",
          5242 => x"81",
          5243 => x"51",
          5244 => x"16",
          5245 => x"84",
          5246 => x"81",
          5247 => x"38",
          5248 => x"ae",
          5249 => x"81",
          5250 => x"54",
          5251 => x"2e",
          5252 => x"8f",
          5253 => x"82",
          5254 => x"76",
          5255 => x"54",
          5256 => x"09",
          5257 => x"38",
          5258 => x"7a",
          5259 => x"80",
          5260 => x"fa",
          5261 => x"93",
          5262 => x"82",
          5263 => x"89",
          5264 => x"08",
          5265 => x"86",
          5266 => x"98",
          5267 => x"82",
          5268 => x"8b",
          5269 => x"fb",
          5270 => x"70",
          5271 => x"81",
          5272 => x"fc",
          5273 => x"93",
          5274 => x"82",
          5275 => x"b4",
          5276 => x"08",
          5277 => x"ec",
          5278 => x"93",
          5279 => x"82",
          5280 => x"a0",
          5281 => x"82",
          5282 => x"52",
          5283 => x"51",
          5284 => x"8b",
          5285 => x"52",
          5286 => x"51",
          5287 => x"81",
          5288 => x"34",
          5289 => x"84",
          5290 => x"0d",
          5291 => x"0d",
          5292 => x"98",
          5293 => x"70",
          5294 => x"ec",
          5295 => x"93",
          5296 => x"38",
          5297 => x"53",
          5298 => x"81",
          5299 => x"34",
          5300 => x"04",
          5301 => x"78",
          5302 => x"80",
          5303 => x"34",
          5304 => x"80",
          5305 => x"38",
          5306 => x"18",
          5307 => x"9c",
          5308 => x"70",
          5309 => x"56",
          5310 => x"a0",
          5311 => x"71",
          5312 => x"81",
          5313 => x"81",
          5314 => x"89",
          5315 => x"06",
          5316 => x"73",
          5317 => x"55",
          5318 => x"55",
          5319 => x"81",
          5320 => x"81",
          5321 => x"74",
          5322 => x"75",
          5323 => x"52",
          5324 => x"13",
          5325 => x"08",
          5326 => x"33",
          5327 => x"9c",
          5328 => x"11",
          5329 => x"8a",
          5330 => x"84",
          5331 => x"96",
          5332 => x"e7",
          5333 => x"84",
          5334 => x"23",
          5335 => x"e7",
          5336 => x"93",
          5337 => x"17",
          5338 => x"0d",
          5339 => x"0d",
          5340 => x"5e",
          5341 => x"70",
          5342 => x"55",
          5343 => x"83",
          5344 => x"73",
          5345 => x"91",
          5346 => x"2e",
          5347 => x"1d",
          5348 => x"0c",
          5349 => x"15",
          5350 => x"70",
          5351 => x"56",
          5352 => x"09",
          5353 => x"38",
          5354 => x"80",
          5355 => x"30",
          5356 => x"78",
          5357 => x"54",
          5358 => x"73",
          5359 => x"60",
          5360 => x"54",
          5361 => x"96",
          5362 => x"0b",
          5363 => x"80",
          5364 => x"f6",
          5365 => x"93",
          5366 => x"85",
          5367 => x"3d",
          5368 => x"5c",
          5369 => x"53",
          5370 => x"51",
          5371 => x"80",
          5372 => x"88",
          5373 => x"5c",
          5374 => x"09",
          5375 => x"d4",
          5376 => x"70",
          5377 => x"71",
          5378 => x"30",
          5379 => x"73",
          5380 => x"51",
          5381 => x"57",
          5382 => x"38",
          5383 => x"75",
          5384 => x"17",
          5385 => x"75",
          5386 => x"30",
          5387 => x"51",
          5388 => x"80",
          5389 => x"38",
          5390 => x"87",
          5391 => x"26",
          5392 => x"77",
          5393 => x"a4",
          5394 => x"27",
          5395 => x"a0",
          5396 => x"39",
          5397 => x"33",
          5398 => x"57",
          5399 => x"27",
          5400 => x"75",
          5401 => x"30",
          5402 => x"32",
          5403 => x"80",
          5404 => x"25",
          5405 => x"56",
          5406 => x"80",
          5407 => x"84",
          5408 => x"58",
          5409 => x"70",
          5410 => x"55",
          5411 => x"09",
          5412 => x"38",
          5413 => x"80",
          5414 => x"30",
          5415 => x"77",
          5416 => x"54",
          5417 => x"81",
          5418 => x"ae",
          5419 => x"06",
          5420 => x"54",
          5421 => x"74",
          5422 => x"80",
          5423 => x"7b",
          5424 => x"30",
          5425 => x"70",
          5426 => x"25",
          5427 => x"07",
          5428 => x"51",
          5429 => x"a7",
          5430 => x"8b",
          5431 => x"39",
          5432 => x"54",
          5433 => x"8c",
          5434 => x"ff",
          5435 => x"f0",
          5436 => x"54",
          5437 => x"e1",
          5438 => x"84",
          5439 => x"b2",
          5440 => x"70",
          5441 => x"71",
          5442 => x"54",
          5443 => x"82",
          5444 => x"80",
          5445 => x"38",
          5446 => x"76",
          5447 => x"df",
          5448 => x"54",
          5449 => x"81",
          5450 => x"55",
          5451 => x"34",
          5452 => x"52",
          5453 => x"51",
          5454 => x"82",
          5455 => x"bf",
          5456 => x"16",
          5457 => x"26",
          5458 => x"16",
          5459 => x"06",
          5460 => x"17",
          5461 => x"34",
          5462 => x"fd",
          5463 => x"19",
          5464 => x"80",
          5465 => x"79",
          5466 => x"81",
          5467 => x"81",
          5468 => x"85",
          5469 => x"54",
          5470 => x"8f",
          5471 => x"86",
          5472 => x"39",
          5473 => x"f3",
          5474 => x"73",
          5475 => x"80",
          5476 => x"52",
          5477 => x"ce",
          5478 => x"84",
          5479 => x"93",
          5480 => x"d7",
          5481 => x"08",
          5482 => x"e6",
          5483 => x"93",
          5484 => x"82",
          5485 => x"80",
          5486 => x"1b",
          5487 => x"55",
          5488 => x"2e",
          5489 => x"8b",
          5490 => x"06",
          5491 => x"1c",
          5492 => x"33",
          5493 => x"70",
          5494 => x"55",
          5495 => x"38",
          5496 => x"52",
          5497 => x"9f",
          5498 => x"84",
          5499 => x"8b",
          5500 => x"7a",
          5501 => x"3f",
          5502 => x"75",
          5503 => x"57",
          5504 => x"2e",
          5505 => x"84",
          5506 => x"06",
          5507 => x"75",
          5508 => x"81",
          5509 => x"2a",
          5510 => x"73",
          5511 => x"38",
          5512 => x"54",
          5513 => x"fb",
          5514 => x"80",
          5515 => x"34",
          5516 => x"c1",
          5517 => x"06",
          5518 => x"38",
          5519 => x"39",
          5520 => x"70",
          5521 => x"54",
          5522 => x"86",
          5523 => x"84",
          5524 => x"06",
          5525 => x"73",
          5526 => x"38",
          5527 => x"83",
          5528 => x"b4",
          5529 => x"51",
          5530 => x"82",
          5531 => x"88",
          5532 => x"ea",
          5533 => x"93",
          5534 => x"3d",
          5535 => x"3d",
          5536 => x"ff",
          5537 => x"71",
          5538 => x"5c",
          5539 => x"80",
          5540 => x"38",
          5541 => x"05",
          5542 => x"a0",
          5543 => x"71",
          5544 => x"38",
          5545 => x"71",
          5546 => x"81",
          5547 => x"38",
          5548 => x"11",
          5549 => x"06",
          5550 => x"70",
          5551 => x"38",
          5552 => x"81",
          5553 => x"05",
          5554 => x"76",
          5555 => x"38",
          5556 => x"ff",
          5557 => x"77",
          5558 => x"57",
          5559 => x"05",
          5560 => x"70",
          5561 => x"33",
          5562 => x"53",
          5563 => x"99",
          5564 => x"e0",
          5565 => x"ff",
          5566 => x"ff",
          5567 => x"70",
          5568 => x"38",
          5569 => x"81",
          5570 => x"51",
          5571 => x"9f",
          5572 => x"72",
          5573 => x"81",
          5574 => x"70",
          5575 => x"72",
          5576 => x"32",
          5577 => x"72",
          5578 => x"73",
          5579 => x"53",
          5580 => x"70",
          5581 => x"38",
          5582 => x"19",
          5583 => x"75",
          5584 => x"38",
          5585 => x"83",
          5586 => x"74",
          5587 => x"59",
          5588 => x"39",
          5589 => x"33",
          5590 => x"93",
          5591 => x"3d",
          5592 => x"3d",
          5593 => x"80",
          5594 => x"34",
          5595 => x"17",
          5596 => x"75",
          5597 => x"3f",
          5598 => x"93",
          5599 => x"80",
          5600 => x"16",
          5601 => x"3f",
          5602 => x"08",
          5603 => x"06",
          5604 => x"73",
          5605 => x"2e",
          5606 => x"80",
          5607 => x"0b",
          5608 => x"56",
          5609 => x"e9",
          5610 => x"06",
          5611 => x"57",
          5612 => x"32",
          5613 => x"80",
          5614 => x"51",
          5615 => x"8a",
          5616 => x"e8",
          5617 => x"06",
          5618 => x"53",
          5619 => x"52",
          5620 => x"51",
          5621 => x"82",
          5622 => x"55",
          5623 => x"08",
          5624 => x"38",
          5625 => x"ff",
          5626 => x"86",
          5627 => x"97",
          5628 => x"84",
          5629 => x"93",
          5630 => x"2e",
          5631 => x"55",
          5632 => x"84",
          5633 => x"0d",
          5634 => x"0d",
          5635 => x"05",
          5636 => x"33",
          5637 => x"75",
          5638 => x"fc",
          5639 => x"93",
          5640 => x"8b",
          5641 => x"82",
          5642 => x"24",
          5643 => x"82",
          5644 => x"84",
          5645 => x"b4",
          5646 => x"55",
          5647 => x"73",
          5648 => x"e6",
          5649 => x"0c",
          5650 => x"06",
          5651 => x"57",
          5652 => x"ae",
          5653 => x"33",
          5654 => x"3f",
          5655 => x"08",
          5656 => x"70",
          5657 => x"55",
          5658 => x"76",
          5659 => x"b8",
          5660 => x"2a",
          5661 => x"51",
          5662 => x"72",
          5663 => x"86",
          5664 => x"74",
          5665 => x"15",
          5666 => x"81",
          5667 => x"d7",
          5668 => x"93",
          5669 => x"ff",
          5670 => x"06",
          5671 => x"56",
          5672 => x"38",
          5673 => x"8f",
          5674 => x"2a",
          5675 => x"51",
          5676 => x"72",
          5677 => x"80",
          5678 => x"52",
          5679 => x"3f",
          5680 => x"08",
          5681 => x"57",
          5682 => x"09",
          5683 => x"e2",
          5684 => x"74",
          5685 => x"56",
          5686 => x"33",
          5687 => x"72",
          5688 => x"38",
          5689 => x"51",
          5690 => x"82",
          5691 => x"57",
          5692 => x"84",
          5693 => x"ff",
          5694 => x"56",
          5695 => x"25",
          5696 => x"0b",
          5697 => x"56",
          5698 => x"05",
          5699 => x"83",
          5700 => x"2e",
          5701 => x"52",
          5702 => x"c6",
          5703 => x"84",
          5704 => x"06",
          5705 => x"27",
          5706 => x"16",
          5707 => x"27",
          5708 => x"56",
          5709 => x"84",
          5710 => x"56",
          5711 => x"84",
          5712 => x"14",
          5713 => x"3f",
          5714 => x"08",
          5715 => x"06",
          5716 => x"80",
          5717 => x"06",
          5718 => x"80",
          5719 => x"db",
          5720 => x"93",
          5721 => x"ff",
          5722 => x"77",
          5723 => x"d8",
          5724 => x"de",
          5725 => x"84",
          5726 => x"9c",
          5727 => x"c4",
          5728 => x"15",
          5729 => x"14",
          5730 => x"70",
          5731 => x"51",
          5732 => x"56",
          5733 => x"84",
          5734 => x"81",
          5735 => x"71",
          5736 => x"16",
          5737 => x"53",
          5738 => x"23",
          5739 => x"8b",
          5740 => x"73",
          5741 => x"80",
          5742 => x"8d",
          5743 => x"39",
          5744 => x"51",
          5745 => x"82",
          5746 => x"53",
          5747 => x"08",
          5748 => x"72",
          5749 => x"8d",
          5750 => x"ce",
          5751 => x"14",
          5752 => x"3f",
          5753 => x"08",
          5754 => x"06",
          5755 => x"38",
          5756 => x"51",
          5757 => x"82",
          5758 => x"55",
          5759 => x"51",
          5760 => x"82",
          5761 => x"83",
          5762 => x"53",
          5763 => x"80",
          5764 => x"38",
          5765 => x"78",
          5766 => x"2a",
          5767 => x"78",
          5768 => x"86",
          5769 => x"22",
          5770 => x"31",
          5771 => x"ad",
          5772 => x"84",
          5773 => x"93",
          5774 => x"2e",
          5775 => x"82",
          5776 => x"80",
          5777 => x"f5",
          5778 => x"83",
          5779 => x"ff",
          5780 => x"38",
          5781 => x"9f",
          5782 => x"38",
          5783 => x"39",
          5784 => x"80",
          5785 => x"38",
          5786 => x"98",
          5787 => x"a0",
          5788 => x"1c",
          5789 => x"0c",
          5790 => x"17",
          5791 => x"76",
          5792 => x"81",
          5793 => x"80",
          5794 => x"d9",
          5795 => x"93",
          5796 => x"ff",
          5797 => x"8d",
          5798 => x"8e",
          5799 => x"8a",
          5800 => x"14",
          5801 => x"3f",
          5802 => x"08",
          5803 => x"74",
          5804 => x"a2",
          5805 => x"79",
          5806 => x"ee",
          5807 => x"a8",
          5808 => x"15",
          5809 => x"2e",
          5810 => x"10",
          5811 => x"2a",
          5812 => x"05",
          5813 => x"ff",
          5814 => x"53",
          5815 => x"9c",
          5816 => x"81",
          5817 => x"0b",
          5818 => x"ff",
          5819 => x"0c",
          5820 => x"84",
          5821 => x"83",
          5822 => x"06",
          5823 => x"80",
          5824 => x"d8",
          5825 => x"93",
          5826 => x"ff",
          5827 => x"72",
          5828 => x"81",
          5829 => x"38",
          5830 => x"73",
          5831 => x"3f",
          5832 => x"08",
          5833 => x"82",
          5834 => x"84",
          5835 => x"b2",
          5836 => x"87",
          5837 => x"84",
          5838 => x"ff",
          5839 => x"82",
          5840 => x"09",
          5841 => x"c8",
          5842 => x"51",
          5843 => x"82",
          5844 => x"84",
          5845 => x"d2",
          5846 => x"06",
          5847 => x"98",
          5848 => x"ee",
          5849 => x"84",
          5850 => x"85",
          5851 => x"09",
          5852 => x"38",
          5853 => x"51",
          5854 => x"82",
          5855 => x"90",
          5856 => x"a0",
          5857 => x"ca",
          5858 => x"84",
          5859 => x"0c",
          5860 => x"82",
          5861 => x"81",
          5862 => x"82",
          5863 => x"72",
          5864 => x"80",
          5865 => x"0c",
          5866 => x"82",
          5867 => x"90",
          5868 => x"fb",
          5869 => x"54",
          5870 => x"80",
          5871 => x"73",
          5872 => x"80",
          5873 => x"72",
          5874 => x"80",
          5875 => x"86",
          5876 => x"15",
          5877 => x"71",
          5878 => x"81",
          5879 => x"81",
          5880 => x"d0",
          5881 => x"93",
          5882 => x"06",
          5883 => x"38",
          5884 => x"54",
          5885 => x"80",
          5886 => x"71",
          5887 => x"82",
          5888 => x"87",
          5889 => x"fa",
          5890 => x"ab",
          5891 => x"58",
          5892 => x"05",
          5893 => x"e6",
          5894 => x"80",
          5895 => x"84",
          5896 => x"38",
          5897 => x"08",
          5898 => x"93",
          5899 => x"08",
          5900 => x"80",
          5901 => x"80",
          5902 => x"54",
          5903 => x"84",
          5904 => x"34",
          5905 => x"75",
          5906 => x"2e",
          5907 => x"53",
          5908 => x"53",
          5909 => x"f7",
          5910 => x"93",
          5911 => x"73",
          5912 => x"0c",
          5913 => x"04",
          5914 => x"67",
          5915 => x"80",
          5916 => x"59",
          5917 => x"78",
          5918 => x"c8",
          5919 => x"06",
          5920 => x"3d",
          5921 => x"99",
          5922 => x"52",
          5923 => x"3f",
          5924 => x"08",
          5925 => x"84",
          5926 => x"38",
          5927 => x"52",
          5928 => x"52",
          5929 => x"3f",
          5930 => x"08",
          5931 => x"84",
          5932 => x"02",
          5933 => x"33",
          5934 => x"55",
          5935 => x"25",
          5936 => x"55",
          5937 => x"54",
          5938 => x"81",
          5939 => x"80",
          5940 => x"74",
          5941 => x"81",
          5942 => x"75",
          5943 => x"3f",
          5944 => x"08",
          5945 => x"02",
          5946 => x"91",
          5947 => x"81",
          5948 => x"82",
          5949 => x"06",
          5950 => x"80",
          5951 => x"88",
          5952 => x"39",
          5953 => x"58",
          5954 => x"38",
          5955 => x"70",
          5956 => x"54",
          5957 => x"81",
          5958 => x"52",
          5959 => x"a5",
          5960 => x"84",
          5961 => x"88",
          5962 => x"62",
          5963 => x"d4",
          5964 => x"54",
          5965 => x"15",
          5966 => x"62",
          5967 => x"e8",
          5968 => x"52",
          5969 => x"51",
          5970 => x"7a",
          5971 => x"83",
          5972 => x"80",
          5973 => x"38",
          5974 => x"08",
          5975 => x"53",
          5976 => x"3d",
          5977 => x"dd",
          5978 => x"93",
          5979 => x"82",
          5980 => x"82",
          5981 => x"39",
          5982 => x"38",
          5983 => x"33",
          5984 => x"70",
          5985 => x"55",
          5986 => x"2e",
          5987 => x"55",
          5988 => x"77",
          5989 => x"81",
          5990 => x"73",
          5991 => x"38",
          5992 => x"54",
          5993 => x"a0",
          5994 => x"82",
          5995 => x"52",
          5996 => x"a3",
          5997 => x"84",
          5998 => x"18",
          5999 => x"55",
          6000 => x"84",
          6001 => x"38",
          6002 => x"70",
          6003 => x"54",
          6004 => x"86",
          6005 => x"c0",
          6006 => x"b0",
          6007 => x"1b",
          6008 => x"1b",
          6009 => x"70",
          6010 => x"d9",
          6011 => x"84",
          6012 => x"84",
          6013 => x"0c",
          6014 => x"52",
          6015 => x"3f",
          6016 => x"08",
          6017 => x"08",
          6018 => x"77",
          6019 => x"86",
          6020 => x"1a",
          6021 => x"1a",
          6022 => x"91",
          6023 => x"0b",
          6024 => x"80",
          6025 => x"0c",
          6026 => x"70",
          6027 => x"54",
          6028 => x"81",
          6029 => x"93",
          6030 => x"2e",
          6031 => x"82",
          6032 => x"94",
          6033 => x"17",
          6034 => x"2b",
          6035 => x"57",
          6036 => x"52",
          6037 => x"9f",
          6038 => x"84",
          6039 => x"93",
          6040 => x"26",
          6041 => x"55",
          6042 => x"08",
          6043 => x"81",
          6044 => x"79",
          6045 => x"31",
          6046 => x"70",
          6047 => x"25",
          6048 => x"76",
          6049 => x"81",
          6050 => x"55",
          6051 => x"38",
          6052 => x"0c",
          6053 => x"75",
          6054 => x"54",
          6055 => x"a2",
          6056 => x"7a",
          6057 => x"3f",
          6058 => x"08",
          6059 => x"55",
          6060 => x"89",
          6061 => x"84",
          6062 => x"1a",
          6063 => x"80",
          6064 => x"54",
          6065 => x"84",
          6066 => x"0d",
          6067 => x"0d",
          6068 => x"64",
          6069 => x"59",
          6070 => x"90",
          6071 => x"52",
          6072 => x"cf",
          6073 => x"84",
          6074 => x"93",
          6075 => x"38",
          6076 => x"55",
          6077 => x"86",
          6078 => x"82",
          6079 => x"19",
          6080 => x"55",
          6081 => x"80",
          6082 => x"38",
          6083 => x"0b",
          6084 => x"82",
          6085 => x"39",
          6086 => x"1a",
          6087 => x"82",
          6088 => x"19",
          6089 => x"08",
          6090 => x"7c",
          6091 => x"74",
          6092 => x"2e",
          6093 => x"94",
          6094 => x"83",
          6095 => x"56",
          6096 => x"38",
          6097 => x"22",
          6098 => x"89",
          6099 => x"55",
          6100 => x"75",
          6101 => x"19",
          6102 => x"39",
          6103 => x"52",
          6104 => x"93",
          6105 => x"84",
          6106 => x"75",
          6107 => x"38",
          6108 => x"ff",
          6109 => x"98",
          6110 => x"19",
          6111 => x"51",
          6112 => x"82",
          6113 => x"80",
          6114 => x"38",
          6115 => x"08",
          6116 => x"2a",
          6117 => x"80",
          6118 => x"38",
          6119 => x"8a",
          6120 => x"5c",
          6121 => x"27",
          6122 => x"7a",
          6123 => x"54",
          6124 => x"52",
          6125 => x"51",
          6126 => x"82",
          6127 => x"fe",
          6128 => x"83",
          6129 => x"56",
          6130 => x"9f",
          6131 => x"08",
          6132 => x"74",
          6133 => x"38",
          6134 => x"b4",
          6135 => x"16",
          6136 => x"89",
          6137 => x"51",
          6138 => x"77",
          6139 => x"b9",
          6140 => x"1a",
          6141 => x"08",
          6142 => x"84",
          6143 => x"57",
          6144 => x"27",
          6145 => x"56",
          6146 => x"52",
          6147 => x"c7",
          6148 => x"84",
          6149 => x"38",
          6150 => x"19",
          6151 => x"06",
          6152 => x"52",
          6153 => x"a2",
          6154 => x"31",
          6155 => x"7f",
          6156 => x"94",
          6157 => x"94",
          6158 => x"5c",
          6159 => x"80",
          6160 => x"93",
          6161 => x"3d",
          6162 => x"3d",
          6163 => x"65",
          6164 => x"5d",
          6165 => x"0c",
          6166 => x"05",
          6167 => x"f6",
          6168 => x"93",
          6169 => x"82",
          6170 => x"8a",
          6171 => x"33",
          6172 => x"2e",
          6173 => x"56",
          6174 => x"90",
          6175 => x"81",
          6176 => x"06",
          6177 => x"87",
          6178 => x"2e",
          6179 => x"95",
          6180 => x"91",
          6181 => x"56",
          6182 => x"81",
          6183 => x"34",
          6184 => x"8e",
          6185 => x"08",
          6186 => x"56",
          6187 => x"84",
          6188 => x"5c",
          6189 => x"82",
          6190 => x"18",
          6191 => x"ff",
          6192 => x"74",
          6193 => x"7e",
          6194 => x"ff",
          6195 => x"2a",
          6196 => x"7a",
          6197 => x"8c",
          6198 => x"08",
          6199 => x"38",
          6200 => x"39",
          6201 => x"52",
          6202 => x"e7",
          6203 => x"84",
          6204 => x"93",
          6205 => x"2e",
          6206 => x"74",
          6207 => x"91",
          6208 => x"2e",
          6209 => x"74",
          6210 => x"88",
          6211 => x"38",
          6212 => x"0c",
          6213 => x"15",
          6214 => x"08",
          6215 => x"06",
          6216 => x"51",
          6217 => x"82",
          6218 => x"fe",
          6219 => x"18",
          6220 => x"51",
          6221 => x"82",
          6222 => x"80",
          6223 => x"38",
          6224 => x"08",
          6225 => x"2a",
          6226 => x"80",
          6227 => x"38",
          6228 => x"8a",
          6229 => x"5b",
          6230 => x"27",
          6231 => x"7b",
          6232 => x"54",
          6233 => x"52",
          6234 => x"51",
          6235 => x"82",
          6236 => x"fe",
          6237 => x"b0",
          6238 => x"31",
          6239 => x"79",
          6240 => x"84",
          6241 => x"16",
          6242 => x"89",
          6243 => x"52",
          6244 => x"cc",
          6245 => x"55",
          6246 => x"16",
          6247 => x"2b",
          6248 => x"39",
          6249 => x"94",
          6250 => x"93",
          6251 => x"cd",
          6252 => x"93",
          6253 => x"e3",
          6254 => x"b0",
          6255 => x"76",
          6256 => x"94",
          6257 => x"ff",
          6258 => x"71",
          6259 => x"7b",
          6260 => x"38",
          6261 => x"18",
          6262 => x"51",
          6263 => x"82",
          6264 => x"fd",
          6265 => x"53",
          6266 => x"18",
          6267 => x"06",
          6268 => x"51",
          6269 => x"7e",
          6270 => x"83",
          6271 => x"76",
          6272 => x"17",
          6273 => x"1e",
          6274 => x"18",
          6275 => x"0c",
          6276 => x"58",
          6277 => x"74",
          6278 => x"38",
          6279 => x"8c",
          6280 => x"90",
          6281 => x"33",
          6282 => x"55",
          6283 => x"34",
          6284 => x"82",
          6285 => x"90",
          6286 => x"f8",
          6287 => x"8b",
          6288 => x"53",
          6289 => x"f2",
          6290 => x"93",
          6291 => x"82",
          6292 => x"80",
          6293 => x"16",
          6294 => x"2a",
          6295 => x"51",
          6296 => x"80",
          6297 => x"38",
          6298 => x"52",
          6299 => x"e7",
          6300 => x"84",
          6301 => x"93",
          6302 => x"d4",
          6303 => x"08",
          6304 => x"a0",
          6305 => x"73",
          6306 => x"88",
          6307 => x"74",
          6308 => x"51",
          6309 => x"8c",
          6310 => x"9c",
          6311 => x"fb",
          6312 => x"b2",
          6313 => x"15",
          6314 => x"3f",
          6315 => x"15",
          6316 => x"3f",
          6317 => x"0b",
          6318 => x"78",
          6319 => x"3f",
          6320 => x"08",
          6321 => x"81",
          6322 => x"57",
          6323 => x"34",
          6324 => x"84",
          6325 => x"0d",
          6326 => x"0d",
          6327 => x"54",
          6328 => x"82",
          6329 => x"53",
          6330 => x"08",
          6331 => x"3d",
          6332 => x"73",
          6333 => x"3f",
          6334 => x"08",
          6335 => x"84",
          6336 => x"82",
          6337 => x"74",
          6338 => x"93",
          6339 => x"3d",
          6340 => x"3d",
          6341 => x"51",
          6342 => x"8b",
          6343 => x"82",
          6344 => x"24",
          6345 => x"93",
          6346 => x"93",
          6347 => x"52",
          6348 => x"84",
          6349 => x"0d",
          6350 => x"0d",
          6351 => x"3d",
          6352 => x"94",
          6353 => x"c1",
          6354 => x"84",
          6355 => x"93",
          6356 => x"e0",
          6357 => x"63",
          6358 => x"d4",
          6359 => x"8d",
          6360 => x"84",
          6361 => x"93",
          6362 => x"38",
          6363 => x"05",
          6364 => x"2b",
          6365 => x"80",
          6366 => x"76",
          6367 => x"0c",
          6368 => x"02",
          6369 => x"70",
          6370 => x"81",
          6371 => x"56",
          6372 => x"9e",
          6373 => x"53",
          6374 => x"db",
          6375 => x"93",
          6376 => x"15",
          6377 => x"82",
          6378 => x"84",
          6379 => x"06",
          6380 => x"55",
          6381 => x"84",
          6382 => x"0d",
          6383 => x"0d",
          6384 => x"5b",
          6385 => x"80",
          6386 => x"ff",
          6387 => x"9f",
          6388 => x"b5",
          6389 => x"84",
          6390 => x"93",
          6391 => x"fc",
          6392 => x"7a",
          6393 => x"08",
          6394 => x"64",
          6395 => x"2e",
          6396 => x"a0",
          6397 => x"70",
          6398 => x"ea",
          6399 => x"84",
          6400 => x"93",
          6401 => x"d4",
          6402 => x"7b",
          6403 => x"3f",
          6404 => x"08",
          6405 => x"84",
          6406 => x"38",
          6407 => x"51",
          6408 => x"82",
          6409 => x"45",
          6410 => x"51",
          6411 => x"82",
          6412 => x"57",
          6413 => x"08",
          6414 => x"80",
          6415 => x"da",
          6416 => x"93",
          6417 => x"82",
          6418 => x"a4",
          6419 => x"7b",
          6420 => x"3f",
          6421 => x"84",
          6422 => x"38",
          6423 => x"51",
          6424 => x"82",
          6425 => x"57",
          6426 => x"08",
          6427 => x"38",
          6428 => x"09",
          6429 => x"38",
          6430 => x"e0",
          6431 => x"dc",
          6432 => x"ff",
          6433 => x"74",
          6434 => x"3f",
          6435 => x"78",
          6436 => x"33",
          6437 => x"56",
          6438 => x"91",
          6439 => x"05",
          6440 => x"81",
          6441 => x"56",
          6442 => x"f5",
          6443 => x"54",
          6444 => x"81",
          6445 => x"80",
          6446 => x"78",
          6447 => x"55",
          6448 => x"11",
          6449 => x"18",
          6450 => x"58",
          6451 => x"34",
          6452 => x"ff",
          6453 => x"55",
          6454 => x"34",
          6455 => x"77",
          6456 => x"81",
          6457 => x"ff",
          6458 => x"55",
          6459 => x"34",
          6460 => x"93",
          6461 => x"84",
          6462 => x"e0",
          6463 => x"70",
          6464 => x"56",
          6465 => x"76",
          6466 => x"81",
          6467 => x"70",
          6468 => x"56",
          6469 => x"82",
          6470 => x"78",
          6471 => x"80",
          6472 => x"27",
          6473 => x"19",
          6474 => x"7a",
          6475 => x"5c",
          6476 => x"55",
          6477 => x"7a",
          6478 => x"5c",
          6479 => x"2e",
          6480 => x"85",
          6481 => x"94",
          6482 => x"81",
          6483 => x"73",
          6484 => x"81",
          6485 => x"7a",
          6486 => x"38",
          6487 => x"76",
          6488 => x"0c",
          6489 => x"04",
          6490 => x"7b",
          6491 => x"fc",
          6492 => x"53",
          6493 => x"bb",
          6494 => x"84",
          6495 => x"93",
          6496 => x"fa",
          6497 => x"33",
          6498 => x"f2",
          6499 => x"08",
          6500 => x"27",
          6501 => x"15",
          6502 => x"2a",
          6503 => x"51",
          6504 => x"83",
          6505 => x"94",
          6506 => x"80",
          6507 => x"0c",
          6508 => x"2e",
          6509 => x"79",
          6510 => x"70",
          6511 => x"51",
          6512 => x"2e",
          6513 => x"52",
          6514 => x"fe",
          6515 => x"82",
          6516 => x"ff",
          6517 => x"70",
          6518 => x"fe",
          6519 => x"82",
          6520 => x"73",
          6521 => x"76",
          6522 => x"06",
          6523 => x"0c",
          6524 => x"98",
          6525 => x"58",
          6526 => x"39",
          6527 => x"54",
          6528 => x"73",
          6529 => x"cd",
          6530 => x"93",
          6531 => x"82",
          6532 => x"81",
          6533 => x"38",
          6534 => x"08",
          6535 => x"9b",
          6536 => x"84",
          6537 => x"0c",
          6538 => x"0c",
          6539 => x"81",
          6540 => x"76",
          6541 => x"38",
          6542 => x"94",
          6543 => x"94",
          6544 => x"16",
          6545 => x"2a",
          6546 => x"51",
          6547 => x"72",
          6548 => x"38",
          6549 => x"51",
          6550 => x"82",
          6551 => x"54",
          6552 => x"08",
          6553 => x"93",
          6554 => x"a7",
          6555 => x"74",
          6556 => x"3f",
          6557 => x"08",
          6558 => x"2e",
          6559 => x"74",
          6560 => x"79",
          6561 => x"14",
          6562 => x"38",
          6563 => x"0c",
          6564 => x"94",
          6565 => x"94",
          6566 => x"83",
          6567 => x"72",
          6568 => x"38",
          6569 => x"51",
          6570 => x"82",
          6571 => x"94",
          6572 => x"91",
          6573 => x"53",
          6574 => x"81",
          6575 => x"34",
          6576 => x"39",
          6577 => x"82",
          6578 => x"05",
          6579 => x"08",
          6580 => x"08",
          6581 => x"38",
          6582 => x"0c",
          6583 => x"80",
          6584 => x"72",
          6585 => x"73",
          6586 => x"53",
          6587 => x"8c",
          6588 => x"16",
          6589 => x"38",
          6590 => x"0c",
          6591 => x"82",
          6592 => x"8b",
          6593 => x"f9",
          6594 => x"56",
          6595 => x"80",
          6596 => x"38",
          6597 => x"3d",
          6598 => x"8a",
          6599 => x"51",
          6600 => x"82",
          6601 => x"55",
          6602 => x"08",
          6603 => x"77",
          6604 => x"52",
          6605 => x"b5",
          6606 => x"84",
          6607 => x"93",
          6608 => x"c3",
          6609 => x"33",
          6610 => x"55",
          6611 => x"24",
          6612 => x"16",
          6613 => x"2a",
          6614 => x"51",
          6615 => x"80",
          6616 => x"9c",
          6617 => x"77",
          6618 => x"3f",
          6619 => x"08",
          6620 => x"77",
          6621 => x"22",
          6622 => x"74",
          6623 => x"ce",
          6624 => x"93",
          6625 => x"74",
          6626 => x"81",
          6627 => x"85",
          6628 => x"74",
          6629 => x"38",
          6630 => x"74",
          6631 => x"93",
          6632 => x"3d",
          6633 => x"3d",
          6634 => x"3d",
          6635 => x"70",
          6636 => x"ff",
          6637 => x"84",
          6638 => x"82",
          6639 => x"73",
          6640 => x"0d",
          6641 => x"0d",
          6642 => x"3d",
          6643 => x"71",
          6644 => x"e7",
          6645 => x"93",
          6646 => x"82",
          6647 => x"80",
          6648 => x"93",
          6649 => x"84",
          6650 => x"51",
          6651 => x"82",
          6652 => x"53",
          6653 => x"82",
          6654 => x"52",
          6655 => x"ac",
          6656 => x"84",
          6657 => x"93",
          6658 => x"2e",
          6659 => x"85",
          6660 => x"87",
          6661 => x"84",
          6662 => x"74",
          6663 => x"d5",
          6664 => x"52",
          6665 => x"89",
          6666 => x"84",
          6667 => x"70",
          6668 => x"07",
          6669 => x"82",
          6670 => x"06",
          6671 => x"54",
          6672 => x"84",
          6673 => x"0d",
          6674 => x"0d",
          6675 => x"53",
          6676 => x"53",
          6677 => x"56",
          6678 => x"82",
          6679 => x"55",
          6680 => x"08",
          6681 => x"52",
          6682 => x"81",
          6683 => x"84",
          6684 => x"93",
          6685 => x"38",
          6686 => x"05",
          6687 => x"2b",
          6688 => x"80",
          6689 => x"86",
          6690 => x"76",
          6691 => x"38",
          6692 => x"51",
          6693 => x"74",
          6694 => x"0c",
          6695 => x"04",
          6696 => x"63",
          6697 => x"80",
          6698 => x"ec",
          6699 => x"3d",
          6700 => x"3f",
          6701 => x"08",
          6702 => x"84",
          6703 => x"38",
          6704 => x"73",
          6705 => x"08",
          6706 => x"13",
          6707 => x"58",
          6708 => x"26",
          6709 => x"7c",
          6710 => x"39",
          6711 => x"cc",
          6712 => x"81",
          6713 => x"93",
          6714 => x"33",
          6715 => x"81",
          6716 => x"06",
          6717 => x"75",
          6718 => x"52",
          6719 => x"05",
          6720 => x"3f",
          6721 => x"08",
          6722 => x"38",
          6723 => x"08",
          6724 => x"38",
          6725 => x"08",
          6726 => x"93",
          6727 => x"80",
          6728 => x"81",
          6729 => x"59",
          6730 => x"14",
          6731 => x"ca",
          6732 => x"39",
          6733 => x"82",
          6734 => x"57",
          6735 => x"38",
          6736 => x"18",
          6737 => x"ff",
          6738 => x"82",
          6739 => x"5b",
          6740 => x"08",
          6741 => x"7c",
          6742 => x"12",
          6743 => x"52",
          6744 => x"82",
          6745 => x"06",
          6746 => x"14",
          6747 => x"cb",
          6748 => x"84",
          6749 => x"ff",
          6750 => x"70",
          6751 => x"82",
          6752 => x"51",
          6753 => x"b4",
          6754 => x"bb",
          6755 => x"93",
          6756 => x"0a",
          6757 => x"70",
          6758 => x"84",
          6759 => x"51",
          6760 => x"ff",
          6761 => x"56",
          6762 => x"38",
          6763 => x"7c",
          6764 => x"0c",
          6765 => x"81",
          6766 => x"74",
          6767 => x"7a",
          6768 => x"0c",
          6769 => x"04",
          6770 => x"79",
          6771 => x"05",
          6772 => x"57",
          6773 => x"82",
          6774 => x"56",
          6775 => x"08",
          6776 => x"91",
          6777 => x"75",
          6778 => x"90",
          6779 => x"81",
          6780 => x"06",
          6781 => x"87",
          6782 => x"2e",
          6783 => x"94",
          6784 => x"73",
          6785 => x"27",
          6786 => x"73",
          6787 => x"93",
          6788 => x"88",
          6789 => x"76",
          6790 => x"3f",
          6791 => x"08",
          6792 => x"0c",
          6793 => x"39",
          6794 => x"52",
          6795 => x"bf",
          6796 => x"93",
          6797 => x"2e",
          6798 => x"83",
          6799 => x"82",
          6800 => x"81",
          6801 => x"06",
          6802 => x"56",
          6803 => x"a0",
          6804 => x"82",
          6805 => x"98",
          6806 => x"94",
          6807 => x"08",
          6808 => x"84",
          6809 => x"51",
          6810 => x"82",
          6811 => x"56",
          6812 => x"8c",
          6813 => x"17",
          6814 => x"07",
          6815 => x"18",
          6816 => x"2e",
          6817 => x"91",
          6818 => x"55",
          6819 => x"84",
          6820 => x"0d",
          6821 => x"0d",
          6822 => x"3d",
          6823 => x"52",
          6824 => x"da",
          6825 => x"93",
          6826 => x"82",
          6827 => x"81",
          6828 => x"45",
          6829 => x"52",
          6830 => x"52",
          6831 => x"3f",
          6832 => x"08",
          6833 => x"84",
          6834 => x"38",
          6835 => x"05",
          6836 => x"2a",
          6837 => x"51",
          6838 => x"55",
          6839 => x"38",
          6840 => x"54",
          6841 => x"81",
          6842 => x"80",
          6843 => x"70",
          6844 => x"54",
          6845 => x"81",
          6846 => x"52",
          6847 => x"c5",
          6848 => x"84",
          6849 => x"2a",
          6850 => x"51",
          6851 => x"80",
          6852 => x"38",
          6853 => x"93",
          6854 => x"15",
          6855 => x"86",
          6856 => x"82",
          6857 => x"5c",
          6858 => x"3d",
          6859 => x"c7",
          6860 => x"93",
          6861 => x"82",
          6862 => x"80",
          6863 => x"93",
          6864 => x"73",
          6865 => x"3f",
          6866 => x"08",
          6867 => x"84",
          6868 => x"87",
          6869 => x"39",
          6870 => x"08",
          6871 => x"38",
          6872 => x"08",
          6873 => x"77",
          6874 => x"3f",
          6875 => x"08",
          6876 => x"08",
          6877 => x"93",
          6878 => x"80",
          6879 => x"55",
          6880 => x"94",
          6881 => x"2e",
          6882 => x"53",
          6883 => x"51",
          6884 => x"82",
          6885 => x"55",
          6886 => x"78",
          6887 => x"fe",
          6888 => x"84",
          6889 => x"82",
          6890 => x"a0",
          6891 => x"e9",
          6892 => x"53",
          6893 => x"05",
          6894 => x"51",
          6895 => x"82",
          6896 => x"54",
          6897 => x"08",
          6898 => x"78",
          6899 => x"8e",
          6900 => x"58",
          6901 => x"82",
          6902 => x"54",
          6903 => x"08",
          6904 => x"54",
          6905 => x"82",
          6906 => x"84",
          6907 => x"06",
          6908 => x"02",
          6909 => x"33",
          6910 => x"81",
          6911 => x"86",
          6912 => x"f6",
          6913 => x"74",
          6914 => x"70",
          6915 => x"c3",
          6916 => x"84",
          6917 => x"56",
          6918 => x"08",
          6919 => x"54",
          6920 => x"08",
          6921 => x"81",
          6922 => x"82",
          6923 => x"84",
          6924 => x"09",
          6925 => x"38",
          6926 => x"b4",
          6927 => x"b0",
          6928 => x"84",
          6929 => x"51",
          6930 => x"82",
          6931 => x"54",
          6932 => x"08",
          6933 => x"8b",
          6934 => x"b4",
          6935 => x"b7",
          6936 => x"54",
          6937 => x"15",
          6938 => x"90",
          6939 => x"34",
          6940 => x"0a",
          6941 => x"19",
          6942 => x"9f",
          6943 => x"78",
          6944 => x"51",
          6945 => x"a0",
          6946 => x"11",
          6947 => x"05",
          6948 => x"b6",
          6949 => x"ae",
          6950 => x"15",
          6951 => x"78",
          6952 => x"53",
          6953 => x"3f",
          6954 => x"0b",
          6955 => x"77",
          6956 => x"3f",
          6957 => x"08",
          6958 => x"84",
          6959 => x"82",
          6960 => x"52",
          6961 => x"51",
          6962 => x"3f",
          6963 => x"52",
          6964 => x"aa",
          6965 => x"90",
          6966 => x"34",
          6967 => x"0b",
          6968 => x"78",
          6969 => x"b6",
          6970 => x"84",
          6971 => x"39",
          6972 => x"52",
          6973 => x"be",
          6974 => x"82",
          6975 => x"99",
          6976 => x"da",
          6977 => x"3d",
          6978 => x"d2",
          6979 => x"53",
          6980 => x"84",
          6981 => x"3d",
          6982 => x"3f",
          6983 => x"08",
          6984 => x"84",
          6985 => x"38",
          6986 => x"3d",
          6987 => x"3d",
          6988 => x"cc",
          6989 => x"93",
          6990 => x"82",
          6991 => x"82",
          6992 => x"81",
          6993 => x"81",
          6994 => x"86",
          6995 => x"aa",
          6996 => x"a4",
          6997 => x"a8",
          6998 => x"05",
          6999 => x"ea",
          7000 => x"77",
          7001 => x"70",
          7002 => x"b4",
          7003 => x"3d",
          7004 => x"51",
          7005 => x"82",
          7006 => x"55",
          7007 => x"08",
          7008 => x"6f",
          7009 => x"06",
          7010 => x"a2",
          7011 => x"92",
          7012 => x"81",
          7013 => x"93",
          7014 => x"2e",
          7015 => x"81",
          7016 => x"51",
          7017 => x"82",
          7018 => x"55",
          7019 => x"08",
          7020 => x"68",
          7021 => x"a8",
          7022 => x"05",
          7023 => x"51",
          7024 => x"3f",
          7025 => x"33",
          7026 => x"8b",
          7027 => x"84",
          7028 => x"06",
          7029 => x"73",
          7030 => x"a0",
          7031 => x"8b",
          7032 => x"54",
          7033 => x"15",
          7034 => x"33",
          7035 => x"70",
          7036 => x"55",
          7037 => x"2e",
          7038 => x"6e",
          7039 => x"df",
          7040 => x"78",
          7041 => x"3f",
          7042 => x"08",
          7043 => x"ff",
          7044 => x"82",
          7045 => x"84",
          7046 => x"80",
          7047 => x"93",
          7048 => x"78",
          7049 => x"af",
          7050 => x"84",
          7051 => x"d4",
          7052 => x"55",
          7053 => x"08",
          7054 => x"81",
          7055 => x"73",
          7056 => x"81",
          7057 => x"63",
          7058 => x"76",
          7059 => x"3f",
          7060 => x"0b",
          7061 => x"87",
          7062 => x"84",
          7063 => x"77",
          7064 => x"3f",
          7065 => x"08",
          7066 => x"84",
          7067 => x"78",
          7068 => x"aa",
          7069 => x"84",
          7070 => x"82",
          7071 => x"a8",
          7072 => x"ed",
          7073 => x"80",
          7074 => x"02",
          7075 => x"df",
          7076 => x"57",
          7077 => x"3d",
          7078 => x"96",
          7079 => x"e9",
          7080 => x"84",
          7081 => x"93",
          7082 => x"cf",
          7083 => x"65",
          7084 => x"d4",
          7085 => x"b5",
          7086 => x"84",
          7087 => x"93",
          7088 => x"38",
          7089 => x"05",
          7090 => x"06",
          7091 => x"73",
          7092 => x"a7",
          7093 => x"09",
          7094 => x"71",
          7095 => x"06",
          7096 => x"55",
          7097 => x"15",
          7098 => x"81",
          7099 => x"34",
          7100 => x"b4",
          7101 => x"93",
          7102 => x"74",
          7103 => x"0c",
          7104 => x"04",
          7105 => x"64",
          7106 => x"93",
          7107 => x"52",
          7108 => x"d1",
          7109 => x"93",
          7110 => x"82",
          7111 => x"80",
          7112 => x"58",
          7113 => x"3d",
          7114 => x"c8",
          7115 => x"93",
          7116 => x"82",
          7117 => x"b4",
          7118 => x"c7",
          7119 => x"a0",
          7120 => x"55",
          7121 => x"84",
          7122 => x"17",
          7123 => x"2b",
          7124 => x"96",
          7125 => x"b0",
          7126 => x"54",
          7127 => x"15",
          7128 => x"ff",
          7129 => x"82",
          7130 => x"55",
          7131 => x"84",
          7132 => x"0d",
          7133 => x"0d",
          7134 => x"5a",
          7135 => x"3d",
          7136 => x"99",
          7137 => x"81",
          7138 => x"84",
          7139 => x"84",
          7140 => x"82",
          7141 => x"07",
          7142 => x"55",
          7143 => x"2e",
          7144 => x"81",
          7145 => x"55",
          7146 => x"2e",
          7147 => x"7b",
          7148 => x"80",
          7149 => x"70",
          7150 => x"be",
          7151 => x"93",
          7152 => x"82",
          7153 => x"80",
          7154 => x"52",
          7155 => x"dc",
          7156 => x"84",
          7157 => x"93",
          7158 => x"38",
          7159 => x"08",
          7160 => x"08",
          7161 => x"56",
          7162 => x"19",
          7163 => x"59",
          7164 => x"74",
          7165 => x"56",
          7166 => x"ec",
          7167 => x"75",
          7168 => x"74",
          7169 => x"2e",
          7170 => x"16",
          7171 => x"33",
          7172 => x"73",
          7173 => x"38",
          7174 => x"84",
          7175 => x"06",
          7176 => x"7a",
          7177 => x"76",
          7178 => x"07",
          7179 => x"54",
          7180 => x"80",
          7181 => x"80",
          7182 => x"7b",
          7183 => x"53",
          7184 => x"93",
          7185 => x"84",
          7186 => x"93",
          7187 => x"38",
          7188 => x"55",
          7189 => x"56",
          7190 => x"8b",
          7191 => x"56",
          7192 => x"83",
          7193 => x"75",
          7194 => x"51",
          7195 => x"3f",
          7196 => x"08",
          7197 => x"82",
          7198 => x"98",
          7199 => x"e6",
          7200 => x"53",
          7201 => x"b8",
          7202 => x"3d",
          7203 => x"3f",
          7204 => x"08",
          7205 => x"08",
          7206 => x"93",
          7207 => x"98",
          7208 => x"a0",
          7209 => x"70",
          7210 => x"ae",
          7211 => x"6d",
          7212 => x"81",
          7213 => x"57",
          7214 => x"74",
          7215 => x"38",
          7216 => x"81",
          7217 => x"81",
          7218 => x"52",
          7219 => x"89",
          7220 => x"84",
          7221 => x"a5",
          7222 => x"33",
          7223 => x"54",
          7224 => x"3f",
          7225 => x"08",
          7226 => x"38",
          7227 => x"76",
          7228 => x"05",
          7229 => x"39",
          7230 => x"08",
          7231 => x"15",
          7232 => x"ff",
          7233 => x"73",
          7234 => x"38",
          7235 => x"83",
          7236 => x"56",
          7237 => x"75",
          7238 => x"81",
          7239 => x"33",
          7240 => x"2e",
          7241 => x"52",
          7242 => x"51",
          7243 => x"3f",
          7244 => x"08",
          7245 => x"ff",
          7246 => x"38",
          7247 => x"88",
          7248 => x"8a",
          7249 => x"38",
          7250 => x"ec",
          7251 => x"75",
          7252 => x"74",
          7253 => x"73",
          7254 => x"05",
          7255 => x"17",
          7256 => x"70",
          7257 => x"34",
          7258 => x"70",
          7259 => x"ff",
          7260 => x"55",
          7261 => x"26",
          7262 => x"8b",
          7263 => x"86",
          7264 => x"e5",
          7265 => x"38",
          7266 => x"99",
          7267 => x"05",
          7268 => x"70",
          7269 => x"73",
          7270 => x"81",
          7271 => x"ff",
          7272 => x"ed",
          7273 => x"80",
          7274 => x"91",
          7275 => x"55",
          7276 => x"3f",
          7277 => x"08",
          7278 => x"84",
          7279 => x"38",
          7280 => x"51",
          7281 => x"3f",
          7282 => x"08",
          7283 => x"84",
          7284 => x"76",
          7285 => x"67",
          7286 => x"34",
          7287 => x"82",
          7288 => x"84",
          7289 => x"06",
          7290 => x"80",
          7291 => x"2e",
          7292 => x"81",
          7293 => x"ff",
          7294 => x"82",
          7295 => x"54",
          7296 => x"08",
          7297 => x"53",
          7298 => x"08",
          7299 => x"ff",
          7300 => x"67",
          7301 => x"8b",
          7302 => x"53",
          7303 => x"51",
          7304 => x"3f",
          7305 => x"0b",
          7306 => x"79",
          7307 => x"ee",
          7308 => x"84",
          7309 => x"55",
          7310 => x"84",
          7311 => x"0d",
          7312 => x"0d",
          7313 => x"88",
          7314 => x"05",
          7315 => x"fc",
          7316 => x"54",
          7317 => x"d2",
          7318 => x"93",
          7319 => x"82",
          7320 => x"82",
          7321 => x"1a",
          7322 => x"82",
          7323 => x"80",
          7324 => x"8c",
          7325 => x"78",
          7326 => x"1a",
          7327 => x"2a",
          7328 => x"51",
          7329 => x"90",
          7330 => x"82",
          7331 => x"58",
          7332 => x"81",
          7333 => x"39",
          7334 => x"22",
          7335 => x"70",
          7336 => x"56",
          7337 => x"e5",
          7338 => x"14",
          7339 => x"30",
          7340 => x"9f",
          7341 => x"84",
          7342 => x"19",
          7343 => x"5a",
          7344 => x"81",
          7345 => x"38",
          7346 => x"77",
          7347 => x"82",
          7348 => x"56",
          7349 => x"74",
          7350 => x"ff",
          7351 => x"81",
          7352 => x"55",
          7353 => x"75",
          7354 => x"82",
          7355 => x"84",
          7356 => x"ff",
          7357 => x"93",
          7358 => x"2e",
          7359 => x"82",
          7360 => x"8e",
          7361 => x"56",
          7362 => x"09",
          7363 => x"38",
          7364 => x"59",
          7365 => x"77",
          7366 => x"06",
          7367 => x"87",
          7368 => x"39",
          7369 => x"ba",
          7370 => x"55",
          7371 => x"2e",
          7372 => x"15",
          7373 => x"2e",
          7374 => x"83",
          7375 => x"75",
          7376 => x"7e",
          7377 => x"a8",
          7378 => x"84",
          7379 => x"93",
          7380 => x"ce",
          7381 => x"16",
          7382 => x"56",
          7383 => x"38",
          7384 => x"19",
          7385 => x"8c",
          7386 => x"7d",
          7387 => x"38",
          7388 => x"0c",
          7389 => x"0c",
          7390 => x"80",
          7391 => x"73",
          7392 => x"98",
          7393 => x"05",
          7394 => x"57",
          7395 => x"26",
          7396 => x"7b",
          7397 => x"0c",
          7398 => x"81",
          7399 => x"84",
          7400 => x"54",
          7401 => x"84",
          7402 => x"0d",
          7403 => x"0d",
          7404 => x"88",
          7405 => x"05",
          7406 => x"54",
          7407 => x"c5",
          7408 => x"56",
          7409 => x"93",
          7410 => x"8b",
          7411 => x"93",
          7412 => x"29",
          7413 => x"05",
          7414 => x"55",
          7415 => x"84",
          7416 => x"34",
          7417 => x"08",
          7418 => x"5f",
          7419 => x"51",
          7420 => x"3f",
          7421 => x"08",
          7422 => x"70",
          7423 => x"57",
          7424 => x"8b",
          7425 => x"82",
          7426 => x"06",
          7427 => x"56",
          7428 => x"38",
          7429 => x"05",
          7430 => x"7e",
          7431 => x"f0",
          7432 => x"84",
          7433 => x"67",
          7434 => x"2e",
          7435 => x"82",
          7436 => x"8b",
          7437 => x"75",
          7438 => x"80",
          7439 => x"81",
          7440 => x"2e",
          7441 => x"80",
          7442 => x"38",
          7443 => x"0a",
          7444 => x"ff",
          7445 => x"55",
          7446 => x"86",
          7447 => x"8a",
          7448 => x"89",
          7449 => x"2a",
          7450 => x"77",
          7451 => x"59",
          7452 => x"81",
          7453 => x"70",
          7454 => x"07",
          7455 => x"56",
          7456 => x"38",
          7457 => x"05",
          7458 => x"7e",
          7459 => x"80",
          7460 => x"82",
          7461 => x"8a",
          7462 => x"83",
          7463 => x"06",
          7464 => x"08",
          7465 => x"74",
          7466 => x"41",
          7467 => x"56",
          7468 => x"8a",
          7469 => x"61",
          7470 => x"55",
          7471 => x"27",
          7472 => x"93",
          7473 => x"80",
          7474 => x"38",
          7475 => x"70",
          7476 => x"43",
          7477 => x"95",
          7478 => x"06",
          7479 => x"2e",
          7480 => x"77",
          7481 => x"74",
          7482 => x"83",
          7483 => x"06",
          7484 => x"82",
          7485 => x"2e",
          7486 => x"78",
          7487 => x"2e",
          7488 => x"80",
          7489 => x"ae",
          7490 => x"2a",
          7491 => x"82",
          7492 => x"56",
          7493 => x"2e",
          7494 => x"77",
          7495 => x"82",
          7496 => x"79",
          7497 => x"70",
          7498 => x"5a",
          7499 => x"86",
          7500 => x"27",
          7501 => x"52",
          7502 => x"e0",
          7503 => x"93",
          7504 => x"29",
          7505 => x"70",
          7506 => x"55",
          7507 => x"0b",
          7508 => x"08",
          7509 => x"05",
          7510 => x"ff",
          7511 => x"27",
          7512 => x"88",
          7513 => x"ae",
          7514 => x"2a",
          7515 => x"82",
          7516 => x"56",
          7517 => x"2e",
          7518 => x"77",
          7519 => x"82",
          7520 => x"79",
          7521 => x"70",
          7522 => x"5a",
          7523 => x"86",
          7524 => x"27",
          7525 => x"52",
          7526 => x"df",
          7527 => x"93",
          7528 => x"84",
          7529 => x"93",
          7530 => x"f5",
          7531 => x"81",
          7532 => x"84",
          7533 => x"93",
          7534 => x"71",
          7535 => x"83",
          7536 => x"5e",
          7537 => x"89",
          7538 => x"5c",
          7539 => x"1c",
          7540 => x"05",
          7541 => x"ff",
          7542 => x"70",
          7543 => x"31",
          7544 => x"57",
          7545 => x"83",
          7546 => x"06",
          7547 => x"1c",
          7548 => x"5c",
          7549 => x"1d",
          7550 => x"29",
          7551 => x"31",
          7552 => x"55",
          7553 => x"87",
          7554 => x"7c",
          7555 => x"7a",
          7556 => x"31",
          7557 => x"de",
          7558 => x"93",
          7559 => x"7d",
          7560 => x"81",
          7561 => x"82",
          7562 => x"83",
          7563 => x"80",
          7564 => x"87",
          7565 => x"81",
          7566 => x"fd",
          7567 => x"f8",
          7568 => x"2e",
          7569 => x"80",
          7570 => x"ff",
          7571 => x"93",
          7572 => x"a0",
          7573 => x"38",
          7574 => x"74",
          7575 => x"86",
          7576 => x"fd",
          7577 => x"81",
          7578 => x"80",
          7579 => x"83",
          7580 => x"39",
          7581 => x"08",
          7582 => x"92",
          7583 => x"b8",
          7584 => x"59",
          7585 => x"27",
          7586 => x"86",
          7587 => x"55",
          7588 => x"09",
          7589 => x"38",
          7590 => x"f5",
          7591 => x"38",
          7592 => x"55",
          7593 => x"86",
          7594 => x"80",
          7595 => x"7a",
          7596 => x"b9",
          7597 => x"81",
          7598 => x"7a",
          7599 => x"8a",
          7600 => x"52",
          7601 => x"ff",
          7602 => x"79",
          7603 => x"7b",
          7604 => x"06",
          7605 => x"51",
          7606 => x"3f",
          7607 => x"1c",
          7608 => x"32",
          7609 => x"96",
          7610 => x"06",
          7611 => x"91",
          7612 => x"a1",
          7613 => x"55",
          7614 => x"ff",
          7615 => x"74",
          7616 => x"06",
          7617 => x"51",
          7618 => x"3f",
          7619 => x"52",
          7620 => x"ff",
          7621 => x"f8",
          7622 => x"34",
          7623 => x"1b",
          7624 => x"d9",
          7625 => x"52",
          7626 => x"ff",
          7627 => x"60",
          7628 => x"51",
          7629 => x"3f",
          7630 => x"09",
          7631 => x"cb",
          7632 => x"b2",
          7633 => x"c3",
          7634 => x"a0",
          7635 => x"52",
          7636 => x"ff",
          7637 => x"82",
          7638 => x"51",
          7639 => x"3f",
          7640 => x"1b",
          7641 => x"95",
          7642 => x"b2",
          7643 => x"a0",
          7644 => x"80",
          7645 => x"1c",
          7646 => x"80",
          7647 => x"93",
          7648 => x"b8",
          7649 => x"1b",
          7650 => x"82",
          7651 => x"52",
          7652 => x"ff",
          7653 => x"7c",
          7654 => x"06",
          7655 => x"51",
          7656 => x"3f",
          7657 => x"a4",
          7658 => x"0b",
          7659 => x"93",
          7660 => x"cc",
          7661 => x"51",
          7662 => x"3f",
          7663 => x"52",
          7664 => x"70",
          7665 => x"9f",
          7666 => x"54",
          7667 => x"52",
          7668 => x"9b",
          7669 => x"56",
          7670 => x"08",
          7671 => x"7d",
          7672 => x"81",
          7673 => x"38",
          7674 => x"86",
          7675 => x"52",
          7676 => x"9b",
          7677 => x"80",
          7678 => x"7a",
          7679 => x"ed",
          7680 => x"85",
          7681 => x"7a",
          7682 => x"8f",
          7683 => x"85",
          7684 => x"83",
          7685 => x"ff",
          7686 => x"ff",
          7687 => x"e8",
          7688 => x"9e",
          7689 => x"52",
          7690 => x"51",
          7691 => x"3f",
          7692 => x"52",
          7693 => x"9e",
          7694 => x"54",
          7695 => x"53",
          7696 => x"51",
          7697 => x"3f",
          7698 => x"16",
          7699 => x"7e",
          7700 => x"d8",
          7701 => x"80",
          7702 => x"ff",
          7703 => x"7f",
          7704 => x"7d",
          7705 => x"81",
          7706 => x"f8",
          7707 => x"ff",
          7708 => x"ff",
          7709 => x"51",
          7710 => x"3f",
          7711 => x"88",
          7712 => x"39",
          7713 => x"f8",
          7714 => x"2e",
          7715 => x"55",
          7716 => x"51",
          7717 => x"3f",
          7718 => x"57",
          7719 => x"83",
          7720 => x"76",
          7721 => x"7a",
          7722 => x"ff",
          7723 => x"82",
          7724 => x"82",
          7725 => x"80",
          7726 => x"84",
          7727 => x"51",
          7728 => x"3f",
          7729 => x"78",
          7730 => x"74",
          7731 => x"18",
          7732 => x"2e",
          7733 => x"79",
          7734 => x"2e",
          7735 => x"55",
          7736 => x"62",
          7737 => x"74",
          7738 => x"75",
          7739 => x"7e",
          7740 => x"b8",
          7741 => x"84",
          7742 => x"38",
          7743 => x"78",
          7744 => x"74",
          7745 => x"56",
          7746 => x"93",
          7747 => x"66",
          7748 => x"26",
          7749 => x"56",
          7750 => x"83",
          7751 => x"64",
          7752 => x"77",
          7753 => x"84",
          7754 => x"52",
          7755 => x"9d",
          7756 => x"d4",
          7757 => x"51",
          7758 => x"3f",
          7759 => x"55",
          7760 => x"81",
          7761 => x"34",
          7762 => x"16",
          7763 => x"16",
          7764 => x"16",
          7765 => x"05",
          7766 => x"c1",
          7767 => x"fe",
          7768 => x"fe",
          7769 => x"34",
          7770 => x"08",
          7771 => x"07",
          7772 => x"16",
          7773 => x"84",
          7774 => x"34",
          7775 => x"c6",
          7776 => x"9c",
          7777 => x"52",
          7778 => x"51",
          7779 => x"3f",
          7780 => x"53",
          7781 => x"51",
          7782 => x"3f",
          7783 => x"93",
          7784 => x"38",
          7785 => x"52",
          7786 => x"99",
          7787 => x"56",
          7788 => x"08",
          7789 => x"39",
          7790 => x"39",
          7791 => x"39",
          7792 => x"08",
          7793 => x"93",
          7794 => x"3d",
          7795 => x"3d",
          7796 => x"5b",
          7797 => x"60",
          7798 => x"57",
          7799 => x"25",
          7800 => x"3d",
          7801 => x"55",
          7802 => x"15",
          7803 => x"c9",
          7804 => x"81",
          7805 => x"06",
          7806 => x"3d",
          7807 => x"8d",
          7808 => x"74",
          7809 => x"05",
          7810 => x"17",
          7811 => x"2e",
          7812 => x"c9",
          7813 => x"34",
          7814 => x"83",
          7815 => x"74",
          7816 => x"0c",
          7817 => x"04",
          7818 => x"7b",
          7819 => x"b3",
          7820 => x"57",
          7821 => x"09",
          7822 => x"38",
          7823 => x"51",
          7824 => x"17",
          7825 => x"76",
          7826 => x"88",
          7827 => x"17",
          7828 => x"59",
          7829 => x"81",
          7830 => x"76",
          7831 => x"8b",
          7832 => x"54",
          7833 => x"17",
          7834 => x"51",
          7835 => x"79",
          7836 => x"30",
          7837 => x"9f",
          7838 => x"53",
          7839 => x"75",
          7840 => x"81",
          7841 => x"0c",
          7842 => x"04",
          7843 => x"79",
          7844 => x"56",
          7845 => x"24",
          7846 => x"3d",
          7847 => x"74",
          7848 => x"52",
          7849 => x"cb",
          7850 => x"93",
          7851 => x"38",
          7852 => x"78",
          7853 => x"06",
          7854 => x"16",
          7855 => x"39",
          7856 => x"82",
          7857 => x"89",
          7858 => x"fd",
          7859 => x"54",
          7860 => x"80",
          7861 => x"ff",
          7862 => x"76",
          7863 => x"3d",
          7864 => x"3d",
          7865 => x"e3",
          7866 => x"53",
          7867 => x"53",
          7868 => x"3f",
          7869 => x"51",
          7870 => x"72",
          7871 => x"3f",
          7872 => x"04",
          7873 => x"7a",
          7874 => x"56",
          7875 => x"80",
          7876 => x"38",
          7877 => x"15",
          7878 => x"16",
          7879 => x"d4",
          7880 => x"54",
          7881 => x"09",
          7882 => x"38",
          7883 => x"f1",
          7884 => x"76",
          7885 => x"8f",
          7886 => x"08",
          7887 => x"da",
          7888 => x"93",
          7889 => x"93",
          7890 => x"75",
          7891 => x"52",
          7892 => x"fd",
          7893 => x"84",
          7894 => x"84",
          7895 => x"73",
          7896 => x"b2",
          7897 => x"70",
          7898 => x"58",
          7899 => x"27",
          7900 => x"54",
          7901 => x"84",
          7902 => x"0d",
          7903 => x"0d",
          7904 => x"93",
          7905 => x"38",
          7906 => x"81",
          7907 => x"52",
          7908 => x"82",
          7909 => x"81",
          7910 => x"82",
          7911 => x"f9",
          7912 => x"ec",
          7913 => x"39",
          7914 => x"51",
          7915 => x"82",
          7916 => x"80",
          7917 => x"83",
          7918 => x"dd",
          7919 => x"b4",
          7920 => x"39",
          7921 => x"51",
          7922 => x"82",
          7923 => x"80",
          7924 => x"83",
          7925 => x"c1",
          7926 => x"8c",
          7927 => x"82",
          7928 => x"b5",
          7929 => x"bc",
          7930 => x"82",
          7931 => x"a9",
          7932 => x"fc",
          7933 => x"82",
          7934 => x"9d",
          7935 => x"b0",
          7936 => x"82",
          7937 => x"91",
          7938 => x"e0",
          7939 => x"82",
          7940 => x"85",
          7941 => x"84",
          7942 => x"ae",
          7943 => x"0d",
          7944 => x"0d",
          7945 => x"56",
          7946 => x"26",
          7947 => x"52",
          7948 => x"29",
          7949 => x"87",
          7950 => x"51",
          7951 => x"3f",
          7952 => x"08",
          7953 => x"fe",
          7954 => x"82",
          7955 => x"54",
          7956 => x"52",
          7957 => x"51",
          7958 => x"3f",
          7959 => x"04",
          7960 => x"66",
          7961 => x"80",
          7962 => x"5b",
          7963 => x"78",
          7964 => x"07",
          7965 => x"57",
          7966 => x"56",
          7967 => x"26",
          7968 => x"56",
          7969 => x"70",
          7970 => x"51",
          7971 => x"74",
          7972 => x"81",
          7973 => x"8c",
          7974 => x"56",
          7975 => x"3f",
          7976 => x"08",
          7977 => x"84",
          7978 => x"82",
          7979 => x"87",
          7980 => x"0c",
          7981 => x"08",
          7982 => x"d4",
          7983 => x"80",
          7984 => x"75",
          7985 => x"3f",
          7986 => x"08",
          7987 => x"84",
          7988 => x"7a",
          7989 => x"2e",
          7990 => x"19",
          7991 => x"59",
          7992 => x"3d",
          7993 => x"cb",
          7994 => x"30",
          7995 => x"80",
          7996 => x"70",
          7997 => x"06",
          7998 => x"56",
          7999 => x"90",
          8000 => x"b8",
          8001 => x"98",
          8002 => x"78",
          8003 => x"3f",
          8004 => x"82",
          8005 => x"96",
          8006 => x"f9",
          8007 => x"02",
          8008 => x"05",
          8009 => x"ff",
          8010 => x"7a",
          8011 => x"fe",
          8012 => x"93",
          8013 => x"38",
          8014 => x"88",
          8015 => x"2e",
          8016 => x"39",
          8017 => x"54",
          8018 => x"53",
          8019 => x"51",
          8020 => x"93",
          8021 => x"83",
          8022 => x"76",
          8023 => x"0c",
          8024 => x"04",
          8025 => x"7f",
          8026 => x"8c",
          8027 => x"05",
          8028 => x"15",
          8029 => x"5c",
          8030 => x"5e",
          8031 => x"86",
          8032 => x"f5",
          8033 => x"86",
          8034 => x"ef",
          8035 => x"55",
          8036 => x"80",
          8037 => x"90",
          8038 => x"7b",
          8039 => x"38",
          8040 => x"74",
          8041 => x"7a",
          8042 => x"72",
          8043 => x"86",
          8044 => x"f4",
          8045 => x"39",
          8046 => x"51",
          8047 => x"3f",
          8048 => x"80",
          8049 => x"18",
          8050 => x"27",
          8051 => x"08",
          8052 => x"c0",
          8053 => x"d6",
          8054 => x"82",
          8055 => x"fe",
          8056 => x"84",
          8057 => x"39",
          8058 => x"72",
          8059 => x"38",
          8060 => x"82",
          8061 => x"fe",
          8062 => x"89",
          8063 => x"e8",
          8064 => x"c6",
          8065 => x"55",
          8066 => x"ed",
          8067 => x"80",
          8068 => x"ec",
          8069 => x"b2",
          8070 => x"74",
          8071 => x"38",
          8072 => x"33",
          8073 => x"56",
          8074 => x"83",
          8075 => x"80",
          8076 => x"27",
          8077 => x"53",
          8078 => x"70",
          8079 => x"51",
          8080 => x"2e",
          8081 => x"80",
          8082 => x"38",
          8083 => x"39",
          8084 => x"ed",
          8085 => x"15",
          8086 => x"82",
          8087 => x"fe",
          8088 => x"78",
          8089 => x"5c",
          8090 => x"94",
          8091 => x"84",
          8092 => x"70",
          8093 => x"57",
          8094 => x"09",
          8095 => x"38",
          8096 => x"3f",
          8097 => x"08",
          8098 => x"98",
          8099 => x"32",
          8100 => x"9b",
          8101 => x"70",
          8102 => x"75",
          8103 => x"58",
          8104 => x"51",
          8105 => x"24",
          8106 => x"9b",
          8107 => x"06",
          8108 => x"53",
          8109 => x"1e",
          8110 => x"26",
          8111 => x"ff",
          8112 => x"93",
          8113 => x"3d",
          8114 => x"3d",
          8115 => x"05",
          8116 => x"f4",
          8117 => x"fc",
          8118 => x"f2",
          8119 => x"8e",
          8120 => x"fe",
          8121 => x"82",
          8122 => x"82",
          8123 => x"82",
          8124 => x"52",
          8125 => x"51",
          8126 => x"3f",
          8127 => x"85",
          8128 => x"a0",
          8129 => x"0d",
          8130 => x"0d",
          8131 => x"80",
          8132 => x"e7",
          8133 => x"51",
          8134 => x"3f",
          8135 => x"51",
          8136 => x"3f",
          8137 => x"d8",
          8138 => x"81",
          8139 => x"06",
          8140 => x"80",
          8141 => x"81",
          8142 => x"d8",
          8143 => x"d4",
          8144 => x"d0",
          8145 => x"fe",
          8146 => x"72",
          8147 => x"81",
          8148 => x"71",
          8149 => x"38",
          8150 => x"d8",
          8151 => x"87",
          8152 => x"da",
          8153 => x"51",
          8154 => x"3f",
          8155 => x"70",
          8156 => x"52",
          8157 => x"95",
          8158 => x"fe",
          8159 => x"82",
          8160 => x"fe",
          8161 => x"80",
          8162 => x"88",
          8163 => x"2a",
          8164 => x"51",
          8165 => x"2e",
          8166 => x"51",
          8167 => x"3f",
          8168 => x"51",
          8169 => x"3f",
          8170 => x"d7",
          8171 => x"85",
          8172 => x"06",
          8173 => x"80",
          8174 => x"81",
          8175 => x"d4",
          8176 => x"a0",
          8177 => x"cc",
          8178 => x"fe",
          8179 => x"72",
          8180 => x"81",
          8181 => x"71",
          8182 => x"38",
          8183 => x"d7",
          8184 => x"88",
          8185 => x"d9",
          8186 => x"51",
          8187 => x"3f",
          8188 => x"70",
          8189 => x"52",
          8190 => x"95",
          8191 => x"fe",
          8192 => x"82",
          8193 => x"fe",
          8194 => x"80",
          8195 => x"84",
          8196 => x"2a",
          8197 => x"51",
          8198 => x"2e",
          8199 => x"51",
          8200 => x"3f",
          8201 => x"51",
          8202 => x"3f",
          8203 => x"d6",
          8204 => x"e5",
          8205 => x"3d",
          8206 => x"3d",
          8207 => x"84",
          8208 => x"33",
          8209 => x"56",
          8210 => x"51",
          8211 => x"3f",
          8212 => x"33",
          8213 => x"38",
          8214 => x"89",
          8215 => x"aa",
          8216 => x"b8",
          8217 => x"93",
          8218 => x"70",
          8219 => x"08",
          8220 => x"82",
          8221 => x"51",
          8222 => x"8f",
          8223 => x"8f",
          8224 => x"73",
          8225 => x"81",
          8226 => x"82",
          8227 => x"74",
          8228 => x"f2",
          8229 => x"93",
          8230 => x"2e",
          8231 => x"93",
          8232 => x"fe",
          8233 => x"8e",
          8234 => x"9c",
          8235 => x"3f",
          8236 => x"8f",
          8237 => x"8f",
          8238 => x"73",
          8239 => x"81",
          8240 => x"74",
          8241 => x"fe",
          8242 => x"80",
          8243 => x"84",
          8244 => x"0d",
          8245 => x"0d",
          8246 => x"82",
          8247 => x"5f",
          8248 => x"7c",
          8249 => x"db",
          8250 => x"84",
          8251 => x"06",
          8252 => x"2e",
          8253 => x"a2",
          8254 => x"ac",
          8255 => x"70",
          8256 => x"ee",
          8257 => x"53",
          8258 => x"94",
          8259 => x"b5",
          8260 => x"93",
          8261 => x"2e",
          8262 => x"89",
          8263 => x"fe",
          8264 => x"5f",
          8265 => x"e8",
          8266 => x"9e",
          8267 => x"70",
          8268 => x"f8",
          8269 => x"fe",
          8270 => x"3d",
          8271 => x"51",
          8272 => x"82",
          8273 => x"90",
          8274 => x"2c",
          8275 => x"80",
          8276 => x"f1",
          8277 => x"c1",
          8278 => x"38",
          8279 => x"83",
          8280 => x"ab",
          8281 => x"78",
          8282 => x"b3",
          8283 => x"24",
          8284 => x"80",
          8285 => x"38",
          8286 => x"78",
          8287 => x"86",
          8288 => x"2e",
          8289 => x"8f",
          8290 => x"bd",
          8291 => x"38",
          8292 => x"90",
          8293 => x"2e",
          8294 => x"78",
          8295 => x"91",
          8296 => x"39",
          8297 => x"85",
          8298 => x"80",
          8299 => x"d2",
          8300 => x"39",
          8301 => x"2e",
          8302 => x"78",
          8303 => x"b0",
          8304 => x"d0",
          8305 => x"38",
          8306 => x"24",
          8307 => x"80",
          8308 => x"99",
          8309 => x"c3",
          8310 => x"38",
          8311 => x"78",
          8312 => x"8c",
          8313 => x"80",
          8314 => x"f3",
          8315 => x"39",
          8316 => x"2e",
          8317 => x"78",
          8318 => x"92",
          8319 => x"f8",
          8320 => x"38",
          8321 => x"2e",
          8322 => x"8e",
          8323 => x"81",
          8324 => x"f7",
          8325 => x"85",
          8326 => x"38",
          8327 => x"b4",
          8328 => x"11",
          8329 => x"05",
          8330 => x"f7",
          8331 => x"84",
          8332 => x"82",
          8333 => x"8f",
          8334 => x"3d",
          8335 => x"53",
          8336 => x"51",
          8337 => x"3f",
          8338 => x"08",
          8339 => x"38",
          8340 => x"83",
          8341 => x"02",
          8342 => x"33",
          8343 => x"cf",
          8344 => x"ff",
          8345 => x"82",
          8346 => x"81",
          8347 => x"78",
          8348 => x"89",
          8349 => x"e5",
          8350 => x"5e",
          8351 => x"82",
          8352 => x"87",
          8353 => x"3d",
          8354 => x"53",
          8355 => x"51",
          8356 => x"3f",
          8357 => x"08",
          8358 => x"89",
          8359 => x"80",
          8360 => x"cf",
          8361 => x"ff",
          8362 => x"82",
          8363 => x"52",
          8364 => x"51",
          8365 => x"b4",
          8366 => x"11",
          8367 => x"05",
          8368 => x"df",
          8369 => x"84",
          8370 => x"87",
          8371 => x"26",
          8372 => x"b4",
          8373 => x"11",
          8374 => x"05",
          8375 => x"c3",
          8376 => x"84",
          8377 => x"82",
          8378 => x"43",
          8379 => x"8a",
          8380 => x"51",
          8381 => x"3f",
          8382 => x"05",
          8383 => x"52",
          8384 => x"29",
          8385 => x"05",
          8386 => x"fb",
          8387 => x"84",
          8388 => x"38",
          8389 => x"51",
          8390 => x"3f",
          8391 => x"85",
          8392 => x"ff",
          8393 => x"fe",
          8394 => x"82",
          8395 => x"b5",
          8396 => x"05",
          8397 => x"cd",
          8398 => x"53",
          8399 => x"08",
          8400 => x"f2",
          8401 => x"d5",
          8402 => x"ff",
          8403 => x"fe",
          8404 => x"82",
          8405 => x"b5",
          8406 => x"05",
          8407 => x"cd",
          8408 => x"93",
          8409 => x"3d",
          8410 => x"52",
          8411 => x"b7",
          8412 => x"84",
          8413 => x"ff",
          8414 => x"59",
          8415 => x"3f",
          8416 => x"58",
          8417 => x"57",
          8418 => x"55",
          8419 => x"08",
          8420 => x"54",
          8421 => x"52",
          8422 => x"ff",
          8423 => x"84",
          8424 => x"fb",
          8425 => x"93",
          8426 => x"ef",
          8427 => x"f5",
          8428 => x"ff",
          8429 => x"ff",
          8430 => x"fe",
          8431 => x"82",
          8432 => x"80",
          8433 => x"38",
          8434 => x"fc",
          8435 => x"84",
          8436 => x"ea",
          8437 => x"93",
          8438 => x"2e",
          8439 => x"b4",
          8440 => x"11",
          8441 => x"05",
          8442 => x"b7",
          8443 => x"84",
          8444 => x"82",
          8445 => x"42",
          8446 => x"51",
          8447 => x"3f",
          8448 => x"5a",
          8449 => x"81",
          8450 => x"59",
          8451 => x"84",
          8452 => x"7a",
          8453 => x"38",
          8454 => x"b4",
          8455 => x"11",
          8456 => x"05",
          8457 => x"fb",
          8458 => x"84",
          8459 => x"f9",
          8460 => x"3d",
          8461 => x"53",
          8462 => x"51",
          8463 => x"3f",
          8464 => x"08",
          8465 => x"dd",
          8466 => x"fe",
          8467 => x"ff",
          8468 => x"fe",
          8469 => x"82",
          8470 => x"80",
          8471 => x"38",
          8472 => x"51",
          8473 => x"3f",
          8474 => x"63",
          8475 => x"38",
          8476 => x"70",
          8477 => x"33",
          8478 => x"81",
          8479 => x"39",
          8480 => x"80",
          8481 => x"84",
          8482 => x"e9",
          8483 => x"93",
          8484 => x"2e",
          8485 => x"b4",
          8486 => x"11",
          8487 => x"05",
          8488 => x"ff",
          8489 => x"84",
          8490 => x"f8",
          8491 => x"3d",
          8492 => x"53",
          8493 => x"51",
          8494 => x"3f",
          8495 => x"08",
          8496 => x"e1",
          8497 => x"cc",
          8498 => x"fe",
          8499 => x"79",
          8500 => x"38",
          8501 => x"7b",
          8502 => x"5b",
          8503 => x"92",
          8504 => x"7a",
          8505 => x"53",
          8506 => x"8a",
          8507 => x"e6",
          8508 => x"1a",
          8509 => x"43",
          8510 => x"82",
          8511 => x"82",
          8512 => x"3d",
          8513 => x"53",
          8514 => x"51",
          8515 => x"3f",
          8516 => x"08",
          8517 => x"82",
          8518 => x"59",
          8519 => x"89",
          8520 => x"80",
          8521 => x"cd",
          8522 => x"c9",
          8523 => x"80",
          8524 => x"82",
          8525 => x"44",
          8526 => x"8e",
          8527 => x"78",
          8528 => x"38",
          8529 => x"08",
          8530 => x"82",
          8531 => x"59",
          8532 => x"88",
          8533 => x"98",
          8534 => x"39",
          8535 => x"33",
          8536 => x"2e",
          8537 => x"8e",
          8538 => x"89",
          8539 => x"b0",
          8540 => x"05",
          8541 => x"fe",
          8542 => x"ff",
          8543 => x"fe",
          8544 => x"82",
          8545 => x"80",
          8546 => x"8e",
          8547 => x"78",
          8548 => x"38",
          8549 => x"08",
          8550 => x"39",
          8551 => x"33",
          8552 => x"2e",
          8553 => x"8e",
          8554 => x"bb",
          8555 => x"ca",
          8556 => x"80",
          8557 => x"82",
          8558 => x"43",
          8559 => x"8e",
          8560 => x"78",
          8561 => x"38",
          8562 => x"08",
          8563 => x"82",
          8564 => x"59",
          8565 => x"88",
          8566 => x"a4",
          8567 => x"39",
          8568 => x"08",
          8569 => x"b4",
          8570 => x"11",
          8571 => x"05",
          8572 => x"af",
          8573 => x"84",
          8574 => x"a7",
          8575 => x"5c",
          8576 => x"2e",
          8577 => x"5c",
          8578 => x"70",
          8579 => x"07",
          8580 => x"7f",
          8581 => x"5a",
          8582 => x"2e",
          8583 => x"a0",
          8584 => x"88",
          8585 => x"f8",
          8586 => x"9e",
          8587 => x"63",
          8588 => x"62",
          8589 => x"ee",
          8590 => x"8b",
          8591 => x"de",
          8592 => x"e1",
          8593 => x"ff",
          8594 => x"ff",
          8595 => x"fe",
          8596 => x"82",
          8597 => x"80",
          8598 => x"38",
          8599 => x"fc",
          8600 => x"84",
          8601 => x"e5",
          8602 => x"93",
          8603 => x"2e",
          8604 => x"59",
          8605 => x"05",
          8606 => x"63",
          8607 => x"b4",
          8608 => x"11",
          8609 => x"05",
          8610 => x"97",
          8611 => x"84",
          8612 => x"f5",
          8613 => x"70",
          8614 => x"82",
          8615 => x"fe",
          8616 => x"80",
          8617 => x"51",
          8618 => x"3f",
          8619 => x"33",
          8620 => x"2e",
          8621 => x"9f",
          8622 => x"38",
          8623 => x"fc",
          8624 => x"84",
          8625 => x"e4",
          8626 => x"93",
          8627 => x"2e",
          8628 => x"59",
          8629 => x"05",
          8630 => x"63",
          8631 => x"ff",
          8632 => x"8b",
          8633 => x"dc",
          8634 => x"aa",
          8635 => x"fe",
          8636 => x"ff",
          8637 => x"fe",
          8638 => x"82",
          8639 => x"80",
          8640 => x"38",
          8641 => x"f0",
          8642 => x"84",
          8643 => x"e6",
          8644 => x"93",
          8645 => x"2e",
          8646 => x"59",
          8647 => x"22",
          8648 => x"05",
          8649 => x"41",
          8650 => x"f0",
          8651 => x"84",
          8652 => x"e5",
          8653 => x"93",
          8654 => x"38",
          8655 => x"60",
          8656 => x"52",
          8657 => x"51",
          8658 => x"3f",
          8659 => x"79",
          8660 => x"b4",
          8661 => x"79",
          8662 => x"ae",
          8663 => x"38",
          8664 => x"87",
          8665 => x"05",
          8666 => x"b4",
          8667 => x"11",
          8668 => x"05",
          8669 => x"9d",
          8670 => x"84",
          8671 => x"92",
          8672 => x"02",
          8673 => x"79",
          8674 => x"5b",
          8675 => x"ff",
          8676 => x"8b",
          8677 => x"db",
          8678 => x"a3",
          8679 => x"fe",
          8680 => x"ff",
          8681 => x"fe",
          8682 => x"82",
          8683 => x"80",
          8684 => x"38",
          8685 => x"f0",
          8686 => x"84",
          8687 => x"e4",
          8688 => x"93",
          8689 => x"2e",
          8690 => x"60",
          8691 => x"60",
          8692 => x"b4",
          8693 => x"11",
          8694 => x"05",
          8695 => x"b5",
          8696 => x"84",
          8697 => x"f2",
          8698 => x"70",
          8699 => x"82",
          8700 => x"fe",
          8701 => x"80",
          8702 => x"51",
          8703 => x"3f",
          8704 => x"33",
          8705 => x"2e",
          8706 => x"9f",
          8707 => x"38",
          8708 => x"f0",
          8709 => x"84",
          8710 => x"e3",
          8711 => x"93",
          8712 => x"2e",
          8713 => x"60",
          8714 => x"60",
          8715 => x"ff",
          8716 => x"8b",
          8717 => x"da",
          8718 => x"ae",
          8719 => x"c0",
          8720 => x"86",
          8721 => x"fe",
          8722 => x"f1",
          8723 => x"8b",
          8724 => x"d9",
          8725 => x"51",
          8726 => x"3f",
          8727 => x"82",
          8728 => x"fe",
          8729 => x"84",
          8730 => x"87",
          8731 => x"0c",
          8732 => x"0b",
          8733 => x"94",
          8734 => x"39",
          8735 => x"51",
          8736 => x"3f",
          8737 => x"0b",
          8738 => x"84",
          8739 => x"83",
          8740 => x"94",
          8741 => x"8d",
          8742 => x"ff",
          8743 => x"ff",
          8744 => x"fe",
          8745 => x"82",
          8746 => x"80",
          8747 => x"38",
          8748 => x"8c",
          8749 => x"de",
          8750 => x"59",
          8751 => x"3d",
          8752 => x"53",
          8753 => x"51",
          8754 => x"3f",
          8755 => x"08",
          8756 => x"d1",
          8757 => x"82",
          8758 => x"fe",
          8759 => x"63",
          8760 => x"82",
          8761 => x"80",
          8762 => x"38",
          8763 => x"08",
          8764 => x"d0",
          8765 => x"b6",
          8766 => x"39",
          8767 => x"51",
          8768 => x"3f",
          8769 => x"3f",
          8770 => x"82",
          8771 => x"fe",
          8772 => x"80",
          8773 => x"39",
          8774 => x"3f",
          8775 => x"79",
          8776 => x"59",
          8777 => x"ef",
          8778 => x"7d",
          8779 => x"80",
          8780 => x"38",
          8781 => x"84",
          8782 => x"c1",
          8783 => x"93",
          8784 => x"81",
          8785 => x"2e",
          8786 => x"82",
          8787 => x"7b",
          8788 => x"38",
          8789 => x"7b",
          8790 => x"38",
          8791 => x"82",
          8792 => x"7a",
          8793 => x"a0",
          8794 => x"82",
          8795 => x"b4",
          8796 => x"05",
          8797 => x"cc",
          8798 => x"82",
          8799 => x"b4",
          8800 => x"05",
          8801 => x"bc",
          8802 => x"7a",
          8803 => x"a0",
          8804 => x"82",
          8805 => x"b4",
          8806 => x"05",
          8807 => x"a4",
          8808 => x"7a",
          8809 => x"82",
          8810 => x"b4",
          8811 => x"05",
          8812 => x"90",
          8813 => x"80",
          8814 => x"cc",
          8815 => x"64",
          8816 => x"83",
          8817 => x"83",
          8818 => x"b4",
          8819 => x"05",
          8820 => x"3f",
          8821 => x"08",
          8822 => x"08",
          8823 => x"70",
          8824 => x"25",
          8825 => x"5f",
          8826 => x"83",
          8827 => x"81",
          8828 => x"06",
          8829 => x"2e",
          8830 => x"1c",
          8831 => x"06",
          8832 => x"fe",
          8833 => x"81",
          8834 => x"32",
          8835 => x"8a",
          8836 => x"2e",
          8837 => x"ee",
          8838 => x"8d",
          8839 => x"dc",
          8840 => x"81",
          8841 => x"0d",
          8842 => x"93",
          8843 => x"c0",
          8844 => x"08",
          8845 => x"84",
          8846 => x"51",
          8847 => x"3f",
          8848 => x"08",
          8849 => x"08",
          8850 => x"84",
          8851 => x"51",
          8852 => x"3f",
          8853 => x"84",
          8854 => x"0c",
          8855 => x"9c",
          8856 => x"55",
          8857 => x"52",
          8858 => x"b5",
          8859 => x"93",
          8860 => x"2b",
          8861 => x"53",
          8862 => x"52",
          8863 => x"b5",
          8864 => x"82",
          8865 => x"07",
          8866 => x"80",
          8867 => x"c0",
          8868 => x"8c",
          8869 => x"87",
          8870 => x"0c",
          8871 => x"82",
          8872 => x"ba",
          8873 => x"93",
          8874 => x"c6",
          8875 => x"d0",
          8876 => x"8d",
          8877 => x"d5",
          8878 => x"8d",
          8879 => x"d5",
          8880 => x"de",
          8881 => x"cf",
          8882 => x"51",
          8883 => x"ec",
          8884 => x"04",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"64",
          8923 => x"2f",
          8924 => x"25",
          8925 => x"64",
          8926 => x"2e",
          8927 => x"64",
          8928 => x"6f",
          8929 => x"6f",
          8930 => x"67",
          8931 => x"74",
          8932 => x"00",
          8933 => x"28",
          8934 => x"6d",
          8935 => x"43",
          8936 => x"6e",
          8937 => x"29",
          8938 => x"0a",
          8939 => x"69",
          8940 => x"20",
          8941 => x"6c",
          8942 => x"6e",
          8943 => x"3a",
          8944 => x"20",
          8945 => x"42",
          8946 => x"52",
          8947 => x"20",
          8948 => x"38",
          8949 => x"30",
          8950 => x"2e",
          8951 => x"20",
          8952 => x"44",
          8953 => x"20",
          8954 => x"20",
          8955 => x"38",
          8956 => x"30",
          8957 => x"2e",
          8958 => x"20",
          8959 => x"4e",
          8960 => x"42",
          8961 => x"20",
          8962 => x"38",
          8963 => x"30",
          8964 => x"2e",
          8965 => x"20",
          8966 => x"52",
          8967 => x"20",
          8968 => x"20",
          8969 => x"38",
          8970 => x"30",
          8971 => x"2e",
          8972 => x"20",
          8973 => x"41",
          8974 => x"20",
          8975 => x"20",
          8976 => x"38",
          8977 => x"30",
          8978 => x"2e",
          8979 => x"20",
          8980 => x"44",
          8981 => x"52",
          8982 => x"20",
          8983 => x"76",
          8984 => x"73",
          8985 => x"30",
          8986 => x"2e",
          8987 => x"20",
          8988 => x"49",
          8989 => x"31",
          8990 => x"20",
          8991 => x"6d",
          8992 => x"20",
          8993 => x"30",
          8994 => x"2e",
          8995 => x"20",
          8996 => x"4e",
          8997 => x"43",
          8998 => x"20",
          8999 => x"61",
          9000 => x"6c",
          9001 => x"30",
          9002 => x"2e",
          9003 => x"20",
          9004 => x"49",
          9005 => x"4f",
          9006 => x"42",
          9007 => x"00",
          9008 => x"20",
          9009 => x"42",
          9010 => x"43",
          9011 => x"20",
          9012 => x"4f",
          9013 => x"0a",
          9014 => x"20",
          9015 => x"53",
          9016 => x"00",
          9017 => x"20",
          9018 => x"50",
          9019 => x"00",
          9020 => x"64",
          9021 => x"73",
          9022 => x"3a",
          9023 => x"20",
          9024 => x"50",
          9025 => x"65",
          9026 => x"20",
          9027 => x"74",
          9028 => x"41",
          9029 => x"65",
          9030 => x"3d",
          9031 => x"38",
          9032 => x"00",
          9033 => x"20",
          9034 => x"50",
          9035 => x"65",
          9036 => x"79",
          9037 => x"61",
          9038 => x"41",
          9039 => x"65",
          9040 => x"3d",
          9041 => x"38",
          9042 => x"00",
          9043 => x"20",
          9044 => x"74",
          9045 => x"20",
          9046 => x"72",
          9047 => x"64",
          9048 => x"73",
          9049 => x"20",
          9050 => x"3d",
          9051 => x"38",
          9052 => x"00",
          9053 => x"69",
          9054 => x"0a",
          9055 => x"20",
          9056 => x"50",
          9057 => x"64",
          9058 => x"20",
          9059 => x"20",
          9060 => x"20",
          9061 => x"20",
          9062 => x"3d",
          9063 => x"34",
          9064 => x"00",
          9065 => x"20",
          9066 => x"79",
          9067 => x"6d",
          9068 => x"6f",
          9069 => x"46",
          9070 => x"20",
          9071 => x"20",
          9072 => x"3d",
          9073 => x"2e",
          9074 => x"64",
          9075 => x"0a",
          9076 => x"20",
          9077 => x"44",
          9078 => x"20",
          9079 => x"63",
          9080 => x"72",
          9081 => x"20",
          9082 => x"20",
          9083 => x"3d",
          9084 => x"2e",
          9085 => x"64",
          9086 => x"0a",
          9087 => x"20",
          9088 => x"69",
          9089 => x"6f",
          9090 => x"53",
          9091 => x"4d",
          9092 => x"6f",
          9093 => x"46",
          9094 => x"3d",
          9095 => x"2e",
          9096 => x"64",
          9097 => x"0a",
          9098 => x"6d",
          9099 => x"00",
          9100 => x"65",
          9101 => x"6d",
          9102 => x"6c",
          9103 => x"00",
          9104 => x"56",
          9105 => x"56",
          9106 => x"6e",
          9107 => x"6e",
          9108 => x"77",
          9109 => x"69",
          9110 => x"72",
          9111 => x"78",
          9112 => x"69",
          9113 => x"72",
          9114 => x"69",
          9115 => x"00",
          9116 => x"00",
          9117 => x"30",
          9118 => x"20",
          9119 => x"00",
          9120 => x"61",
          9121 => x"64",
          9122 => x"20",
          9123 => x"65",
          9124 => x"68",
          9125 => x"69",
          9126 => x"72",
          9127 => x"69",
          9128 => x"74",
          9129 => x"4f",
          9130 => x"00",
          9131 => x"61",
          9132 => x"74",
          9133 => x"65",
          9134 => x"72",
          9135 => x"65",
          9136 => x"73",
          9137 => x"79",
          9138 => x"6c",
          9139 => x"64",
          9140 => x"62",
          9141 => x"67",
          9142 => x"00",
          9143 => x"00",
          9144 => x"00",
          9145 => x"00",
          9146 => x"00",
          9147 => x"00",
          9148 => x"00",
          9149 => x"00",
          9150 => x"00",
          9151 => x"00",
          9152 => x"00",
          9153 => x"00",
          9154 => x"00",
          9155 => x"00",
          9156 => x"00",
          9157 => x"00",
          9158 => x"00",
          9159 => x"00",
          9160 => x"00",
          9161 => x"00",
          9162 => x"00",
          9163 => x"00",
          9164 => x"00",
          9165 => x"00",
          9166 => x"00",
          9167 => x"00",
          9168 => x"00",
          9169 => x"00",
          9170 => x"00",
          9171 => x"00",
          9172 => x"00",
          9173 => x"00",
          9174 => x"00",
          9175 => x"00",
          9176 => x"5b",
          9177 => x"5b",
          9178 => x"5b",
          9179 => x"5b",
          9180 => x"5b",
          9181 => x"5b",
          9182 => x"5b",
          9183 => x"5b",
          9184 => x"5b",
          9185 => x"00",
          9186 => x"00",
          9187 => x"44",
          9188 => x"2a",
          9189 => x"3b",
          9190 => x"3f",
          9191 => x"7f",
          9192 => x"41",
          9193 => x"41",
          9194 => x"00",
          9195 => x"fe",
          9196 => x"44",
          9197 => x"2e",
          9198 => x"4f",
          9199 => x"4d",
          9200 => x"20",
          9201 => x"54",
          9202 => x"20",
          9203 => x"4f",
          9204 => x"4d",
          9205 => x"20",
          9206 => x"54",
          9207 => x"20",
          9208 => x"00",
          9209 => x"00",
          9210 => x"00",
          9211 => x"00",
          9212 => x"9a",
          9213 => x"41",
          9214 => x"45",
          9215 => x"49",
          9216 => x"92",
          9217 => x"4f",
          9218 => x"99",
          9219 => x"9d",
          9220 => x"49",
          9221 => x"a5",
          9222 => x"a9",
          9223 => x"ad",
          9224 => x"b1",
          9225 => x"b5",
          9226 => x"b9",
          9227 => x"bd",
          9228 => x"c1",
          9229 => x"c5",
          9230 => x"c9",
          9231 => x"cd",
          9232 => x"d1",
          9233 => x"d5",
          9234 => x"d9",
          9235 => x"dd",
          9236 => x"e1",
          9237 => x"e5",
          9238 => x"e9",
          9239 => x"ed",
          9240 => x"f1",
          9241 => x"f5",
          9242 => x"f9",
          9243 => x"fd",
          9244 => x"2e",
          9245 => x"5b",
          9246 => x"22",
          9247 => x"3e",
          9248 => x"00",
          9249 => x"01",
          9250 => x"10",
          9251 => x"00",
          9252 => x"00",
          9253 => x"01",
          9254 => x"04",
          9255 => x"10",
          9256 => x"00",
          9257 => x"69",
          9258 => x"00",
          9259 => x"69",
          9260 => x"6c",
          9261 => x"69",
          9262 => x"00",
          9263 => x"6c",
          9264 => x"00",
          9265 => x"65",
          9266 => x"00",
          9267 => x"63",
          9268 => x"72",
          9269 => x"63",
          9270 => x"00",
          9271 => x"64",
          9272 => x"00",
          9273 => x"64",
          9274 => x"00",
          9275 => x"65",
          9276 => x"65",
          9277 => x"65",
          9278 => x"69",
          9279 => x"69",
          9280 => x"66",
          9281 => x"66",
          9282 => x"61",
          9283 => x"00",
          9284 => x"6d",
          9285 => x"65",
          9286 => x"72",
          9287 => x"65",
          9288 => x"00",
          9289 => x"6e",
          9290 => x"00",
          9291 => x"65",
          9292 => x"00",
          9293 => x"62",
          9294 => x"63",
          9295 => x"62",
          9296 => x"63",
          9297 => x"69",
          9298 => x"00",
          9299 => x"69",
          9300 => x"45",
          9301 => x"72",
          9302 => x"6e",
          9303 => x"6e",
          9304 => x"65",
          9305 => x"72",
          9306 => x"00",
          9307 => x"69",
          9308 => x"6e",
          9309 => x"72",
          9310 => x"79",
          9311 => x"00",
          9312 => x"6f",
          9313 => x"6c",
          9314 => x"6f",
          9315 => x"2e",
          9316 => x"6f",
          9317 => x"74",
          9318 => x"6f",
          9319 => x"2e",
          9320 => x"6e",
          9321 => x"69",
          9322 => x"69",
          9323 => x"61",
          9324 => x"0a",
          9325 => x"63",
          9326 => x"73",
          9327 => x"6e",
          9328 => x"2e",
          9329 => x"69",
          9330 => x"61",
          9331 => x"61",
          9332 => x"65",
          9333 => x"74",
          9334 => x"00",
          9335 => x"69",
          9336 => x"68",
          9337 => x"6c",
          9338 => x"6e",
          9339 => x"69",
          9340 => x"00",
          9341 => x"44",
          9342 => x"20",
          9343 => x"74",
          9344 => x"72",
          9345 => x"63",
          9346 => x"2e",
          9347 => x"72",
          9348 => x"20",
          9349 => x"62",
          9350 => x"69",
          9351 => x"6e",
          9352 => x"69",
          9353 => x"00",
          9354 => x"69",
          9355 => x"6e",
          9356 => x"65",
          9357 => x"6c",
          9358 => x"0a",
          9359 => x"6f",
          9360 => x"6d",
          9361 => x"69",
          9362 => x"20",
          9363 => x"65",
          9364 => x"74",
          9365 => x"66",
          9366 => x"64",
          9367 => x"20",
          9368 => x"6b",
          9369 => x"00",
          9370 => x"6f",
          9371 => x"74",
          9372 => x"6f",
          9373 => x"64",
          9374 => x"00",
          9375 => x"69",
          9376 => x"75",
          9377 => x"6f",
          9378 => x"61",
          9379 => x"6e",
          9380 => x"6e",
          9381 => x"6c",
          9382 => x"0a",
          9383 => x"69",
          9384 => x"69",
          9385 => x"6f",
          9386 => x"64",
          9387 => x"00",
          9388 => x"6e",
          9389 => x"66",
          9390 => x"65",
          9391 => x"6d",
          9392 => x"72",
          9393 => x"00",
          9394 => x"6f",
          9395 => x"61",
          9396 => x"6f",
          9397 => x"20",
          9398 => x"65",
          9399 => x"00",
          9400 => x"61",
          9401 => x"65",
          9402 => x"73",
          9403 => x"63",
          9404 => x"65",
          9405 => x"0a",
          9406 => x"75",
          9407 => x"73",
          9408 => x"00",
          9409 => x"6e",
          9410 => x"77",
          9411 => x"72",
          9412 => x"2e",
          9413 => x"25",
          9414 => x"62",
          9415 => x"73",
          9416 => x"20",
          9417 => x"25",
          9418 => x"62",
          9419 => x"73",
          9420 => x"63",
          9421 => x"00",
          9422 => x"65",
          9423 => x"00",
          9424 => x"30",
          9425 => x"00",
          9426 => x"20",
          9427 => x"30",
          9428 => x"00",
          9429 => x"20",
          9430 => x"20",
          9431 => x"00",
          9432 => x"30",
          9433 => x"00",
          9434 => x"20",
          9435 => x"7c",
          9436 => x"0d",
          9437 => x"50",
          9438 => x"00",
          9439 => x"2a",
          9440 => x"73",
          9441 => x"00",
          9442 => x"31",
          9443 => x"2f",
          9444 => x"30",
          9445 => x"31",
          9446 => x"00",
          9447 => x"5a",
          9448 => x"20",
          9449 => x"20",
          9450 => x"78",
          9451 => x"73",
          9452 => x"20",
          9453 => x"0a",
          9454 => x"50",
          9455 => x"20",
          9456 => x"65",
          9457 => x"70",
          9458 => x"61",
          9459 => x"65",
          9460 => x"00",
          9461 => x"69",
          9462 => x"20",
          9463 => x"65",
          9464 => x"70",
          9465 => x"00",
          9466 => x"53",
          9467 => x"6e",
          9468 => x"72",
          9469 => x"0a",
          9470 => x"4f",
          9471 => x"20",
          9472 => x"69",
          9473 => x"72",
          9474 => x"74",
          9475 => x"4f",
          9476 => x"20",
          9477 => x"69",
          9478 => x"72",
          9479 => x"74",
          9480 => x"41",
          9481 => x"20",
          9482 => x"69",
          9483 => x"72",
          9484 => x"74",
          9485 => x"41",
          9486 => x"20",
          9487 => x"69",
          9488 => x"72",
          9489 => x"74",
          9490 => x"41",
          9491 => x"20",
          9492 => x"69",
          9493 => x"72",
          9494 => x"74",
          9495 => x"41",
          9496 => x"20",
          9497 => x"69",
          9498 => x"72",
          9499 => x"74",
          9500 => x"65",
          9501 => x"6e",
          9502 => x"70",
          9503 => x"6d",
          9504 => x"2e",
          9505 => x"00",
          9506 => x"6e",
          9507 => x"69",
          9508 => x"74",
          9509 => x"72",
          9510 => x"0a",
          9511 => x"75",
          9512 => x"78",
          9513 => x"62",
          9514 => x"00",
          9515 => x"3a",
          9516 => x"61",
          9517 => x"64",
          9518 => x"20",
          9519 => x"74",
          9520 => x"69",
          9521 => x"73",
          9522 => x"61",
          9523 => x"30",
          9524 => x"6c",
          9525 => x"65",
          9526 => x"69",
          9527 => x"61",
          9528 => x"6c",
          9529 => x"0a",
          9530 => x"20",
          9531 => x"61",
          9532 => x"69",
          9533 => x"69",
          9534 => x"00",
          9535 => x"6e",
          9536 => x"61",
          9537 => x"65",
          9538 => x"00",
          9539 => x"61",
          9540 => x"64",
          9541 => x"20",
          9542 => x"74",
          9543 => x"69",
          9544 => x"0a",
          9545 => x"63",
          9546 => x"0a",
          9547 => x"75",
          9548 => x"6c",
          9549 => x"69",
          9550 => x"2e",
          9551 => x"00",
          9552 => x"6f",
          9553 => x"6e",
          9554 => x"2e",
          9555 => x"6f",
          9556 => x"72",
          9557 => x"2e",
          9558 => x"00",
          9559 => x"30",
          9560 => x"28",
          9561 => x"78",
          9562 => x"25",
          9563 => x"78",
          9564 => x"38",
          9565 => x"00",
          9566 => x"75",
          9567 => x"4d",
          9568 => x"72",
          9569 => x"00",
          9570 => x"43",
          9571 => x"6c",
          9572 => x"2e",
          9573 => x"30",
          9574 => x"25",
          9575 => x"2d",
          9576 => x"3f",
          9577 => x"00",
          9578 => x"30",
          9579 => x"25",
          9580 => x"2d",
          9581 => x"30",
          9582 => x"25",
          9583 => x"2d",
          9584 => x"69",
          9585 => x"6c",
          9586 => x"20",
          9587 => x"65",
          9588 => x"70",
          9589 => x"00",
          9590 => x"6e",
          9591 => x"69",
          9592 => x"69",
          9593 => x"72",
          9594 => x"74",
          9595 => x"00",
          9596 => x"69",
          9597 => x"6c",
          9598 => x"75",
          9599 => x"20",
          9600 => x"6f",
          9601 => x"6e",
          9602 => x"69",
          9603 => x"75",
          9604 => x"20",
          9605 => x"6f",
          9606 => x"78",
          9607 => x"74",
          9608 => x"20",
          9609 => x"65",
          9610 => x"25",
          9611 => x"20",
          9612 => x"0a",
          9613 => x"61",
          9614 => x"6e",
          9615 => x"6f",
          9616 => x"40",
          9617 => x"38",
          9618 => x"2e",
          9619 => x"00",
          9620 => x"61",
          9621 => x"72",
          9622 => x"72",
          9623 => x"20",
          9624 => x"65",
          9625 => x"64",
          9626 => x"00",
          9627 => x"65",
          9628 => x"72",
          9629 => x"67",
          9630 => x"70",
          9631 => x"61",
          9632 => x"6e",
          9633 => x"0a",
          9634 => x"6f",
          9635 => x"72",
          9636 => x"6f",
          9637 => x"67",
          9638 => x"0a",
          9639 => x"50",
          9640 => x"69",
          9641 => x"64",
          9642 => x"73",
          9643 => x"2e",
          9644 => x"00",
          9645 => x"64",
          9646 => x"73",
          9647 => x"00",
          9648 => x"64",
          9649 => x"73",
          9650 => x"61",
          9651 => x"6f",
          9652 => x"6e",
          9653 => x"00",
          9654 => x"75",
          9655 => x"6e",
          9656 => x"2e",
          9657 => x"6e",
          9658 => x"69",
          9659 => x"69",
          9660 => x"72",
          9661 => x"74",
          9662 => x"2e",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"01",
          9669 => x"00",
          9670 => x"01",
          9671 => x"81",
          9672 => x"00",
          9673 => x"7f",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"f5",
          9679 => x"f5",
          9680 => x"f5",
          9681 => x"00",
          9682 => x"01",
          9683 => x"01",
          9684 => x"01",
          9685 => x"00",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"00",
          9719 => x"00",
          9720 => x"00",
          9721 => x"00",
          9722 => x"00",
          9723 => x"00",
          9724 => x"00",
          9725 => x"00",
          9726 => x"02",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"04",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"14",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"2b",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"30",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"3c",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"3d",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"3f",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"40",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"41",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"42",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"43",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"50",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"51",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"54",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"55",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"79",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"78",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"82",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"83",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"85",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"87",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"8c",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"8d",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"8e",
          9823 => x"00",
          9824 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"e0",
             2 => x"00",
             3 => x"00",
             4 => x"00",
             5 => x"00",
             6 => x"00",
             7 => x"00",
             8 => x"88",
             9 => x"90",
            10 => x"0b",
            11 => x"2d",
            12 => x"0c",
            13 => x"00",
            14 => x"00",
            15 => x"00",
            16 => x"71",
            17 => x"72",
            18 => x"81",
            19 => x"83",
            20 => x"ff",
            21 => x"04",
            22 => x"00",
            23 => x"00",
            24 => x"71",
            25 => x"83",
            26 => x"83",
            27 => x"05",
            28 => x"2b",
            29 => x"73",
            30 => x"0b",
            31 => x"83",
            32 => x"72",
            33 => x"72",
            34 => x"09",
            35 => x"73",
            36 => x"07",
            37 => x"53",
            38 => x"00",
            39 => x"00",
            40 => x"72",
            41 => x"73",
            42 => x"51",
            43 => x"00",
            44 => x"00",
            45 => x"00",
            46 => x"00",
            47 => x"00",
            48 => x"71",
            49 => x"71",
            50 => x"09",
            51 => x"0a",
            52 => x"0a",
            53 => x"05",
            54 => x"51",
            55 => x"04",
            56 => x"72",
            57 => x"73",
            58 => x"51",
            59 => x"00",
            60 => x"00",
            61 => x"00",
            62 => x"00",
            63 => x"00",
            64 => x"00",
            65 => x"00",
            66 => x"00",
            67 => x"00",
            68 => x"00",
            69 => x"00",
            70 => x"00",
            71 => x"00",
            72 => x"0b",
            73 => x"c4",
            74 => x"00",
            75 => x"00",
            76 => x"00",
            77 => x"00",
            78 => x"00",
            79 => x"00",
            80 => x"72",
            81 => x"0a",
            82 => x"00",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"72",
            89 => x"09",
            90 => x"0b",
            91 => x"05",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"72",
            97 => x"73",
            98 => x"09",
            99 => x"81",
           100 => x"06",
           101 => x"04",
           102 => x"00",
           103 => x"00",
           104 => x"71",
           105 => x"04",
           106 => x"06",
           107 => x"82",
           108 => x"0b",
           109 => x"fc",
           110 => x"51",
           111 => x"00",
           112 => x"72",
           113 => x"72",
           114 => x"81",
           115 => x"0a",
           116 => x"51",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"72",
           121 => x"72",
           122 => x"81",
           123 => x"0a",
           124 => x"53",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"71",
           129 => x"52",
           130 => x"00",
           131 => x"00",
           132 => x"00",
           133 => x"00",
           134 => x"00",
           135 => x"00",
           136 => x"72",
           137 => x"05",
           138 => x"04",
           139 => x"00",
           140 => x"00",
           141 => x"00",
           142 => x"00",
           143 => x"00",
           144 => x"72",
           145 => x"73",
           146 => x"07",
           147 => x"00",
           148 => x"00",
           149 => x"00",
           150 => x"00",
           151 => x"00",
           152 => x"71",
           153 => x"72",
           154 => x"81",
           155 => x"10",
           156 => x"81",
           157 => x"04",
           158 => x"00",
           159 => x"00",
           160 => x"71",
           161 => x"0b",
           162 => x"d0",
           163 => x"10",
           164 => x"06",
           165 => x"88",
           166 => x"00",
           167 => x"00",
           168 => x"88",
           169 => x"90",
           170 => x"0b",
           171 => x"cf",
           172 => x"88",
           173 => x"0c",
           174 => x"0c",
           175 => x"00",
           176 => x"88",
           177 => x"90",
           178 => x"0b",
           179 => x"81",
           180 => x"88",
           181 => x"0c",
           182 => x"0c",
           183 => x"00",
           184 => x"72",
           185 => x"05",
           186 => x"81",
           187 => x"70",
           188 => x"73",
           189 => x"05",
           190 => x"07",
           191 => x"04",
           192 => x"72",
           193 => x"05",
           194 => x"09",
           195 => x"05",
           196 => x"06",
           197 => x"74",
           198 => x"06",
           199 => x"51",
           200 => x"05",
           201 => x"00",
           202 => x"00",
           203 => x"00",
           204 => x"00",
           205 => x"00",
           206 => x"00",
           207 => x"00",
           208 => x"04",
           209 => x"00",
           210 => x"00",
           211 => x"00",
           212 => x"00",
           213 => x"00",
           214 => x"00",
           215 => x"00",
           216 => x"71",
           217 => x"04",
           218 => x"00",
           219 => x"00",
           220 => x"00",
           221 => x"00",
           222 => x"00",
           223 => x"00",
           224 => x"04",
           225 => x"00",
           226 => x"00",
           227 => x"00",
           228 => x"00",
           229 => x"00",
           230 => x"00",
           231 => x"00",
           232 => x"02",
           233 => x"10",
           234 => x"04",
           235 => x"00",
           236 => x"00",
           237 => x"00",
           238 => x"00",
           239 => x"00",
           240 => x"00",
           241 => x"00",
           242 => x"00",
           243 => x"00",
           244 => x"00",
           245 => x"00",
           246 => x"00",
           247 => x"00",
           248 => x"71",
           249 => x"05",
           250 => x"02",
           251 => x"00",
           252 => x"00",
           253 => x"00",
           254 => x"00",
           255 => x"00",
           256 => x"00",
           257 => x"04",
           258 => x"10",
           259 => x"10",
           260 => x"10",
           261 => x"10",
           262 => x"10",
           263 => x"10",
           264 => x"10",
           265 => x"10",
           266 => x"51",
           267 => x"73",
           268 => x"73",
           269 => x"81",
           270 => x"10",
           271 => x"07",
           272 => x"0c",
           273 => x"72",
           274 => x"81",
           275 => x"09",
           276 => x"71",
           277 => x"0a",
           278 => x"72",
           279 => x"51",
           280 => x"9f",
           281 => x"a4",
           282 => x"80",
           283 => x"05",
           284 => x"0b",
           285 => x"04",
           286 => x"9e",
           287 => x"80",
           288 => x"fe",
           289 => x"00",
           290 => x"94",
           291 => x"0d",
           292 => x"08",
           293 => x"52",
           294 => x"05",
           295 => x"de",
           296 => x"70",
           297 => x"85",
           298 => x"0c",
           299 => x"02",
           300 => x"3d",
           301 => x"94",
           302 => x"08",
           303 => x"88",
           304 => x"82",
           305 => x"08",
           306 => x"54",
           307 => x"94",
           308 => x"08",
           309 => x"f9",
           310 => x"0b",
           311 => x"05",
           312 => x"88",
           313 => x"25",
           314 => x"08",
           315 => x"30",
           316 => x"05",
           317 => x"94",
           318 => x"0c",
           319 => x"05",
           320 => x"81",
           321 => x"f4",
           322 => x"08",
           323 => x"94",
           324 => x"0c",
           325 => x"05",
           326 => x"ab",
           327 => x"8c",
           328 => x"94",
           329 => x"0c",
           330 => x"08",
           331 => x"94",
           332 => x"08",
           333 => x"0b",
           334 => x"05",
           335 => x"f0",
           336 => x"08",
           337 => x"80",
           338 => x"8c",
           339 => x"94",
           340 => x"08",
           341 => x"3f",
           342 => x"94",
           343 => x"0c",
           344 => x"fc",
           345 => x"2e",
           346 => x"08",
           347 => x"30",
           348 => x"05",
           349 => x"f8",
           350 => x"88",
           351 => x"3d",
           352 => x"04",
           353 => x"94",
           354 => x"0d",
           355 => x"08",
           356 => x"94",
           357 => x"08",
           358 => x"38",
           359 => x"05",
           360 => x"08",
           361 => x"81",
           362 => x"fc",
           363 => x"08",
           364 => x"80",
           365 => x"94",
           366 => x"08",
           367 => x"8c",
           368 => x"53",
           369 => x"05",
           370 => x"08",
           371 => x"51",
           372 => x"08",
           373 => x"f8",
           374 => x"94",
           375 => x"08",
           376 => x"38",
           377 => x"05",
           378 => x"08",
           379 => x"94",
           380 => x"08",
           381 => x"54",
           382 => x"94",
           383 => x"08",
           384 => x"fd",
           385 => x"0b",
           386 => x"05",
           387 => x"94",
           388 => x"0c",
           389 => x"05",
           390 => x"88",
           391 => x"ac",
           392 => x"fc",
           393 => x"2e",
           394 => x"0b",
           395 => x"05",
           396 => x"38",
           397 => x"05",
           398 => x"08",
           399 => x"94",
           400 => x"08",
           401 => x"fc",
           402 => x"39",
           403 => x"05",
           404 => x"80",
           405 => x"08",
           406 => x"94",
           407 => x"08",
           408 => x"94",
           409 => x"08",
           410 => x"05",
           411 => x"08",
           412 => x"94",
           413 => x"08",
           414 => x"05",
           415 => x"08",
           416 => x"94",
           417 => x"08",
           418 => x"08",
           419 => x"94",
           420 => x"08",
           421 => x"08",
           422 => x"ff",
           423 => x"08",
           424 => x"80",
           425 => x"94",
           426 => x"08",
           427 => x"f4",
           428 => x"8d",
           429 => x"f8",
           430 => x"94",
           431 => x"0c",
           432 => x"f4",
           433 => x"0c",
           434 => x"94",
           435 => x"3d",
           436 => x"0b",
           437 => x"8c",
           438 => x"87",
           439 => x"0c",
           440 => x"c0",
           441 => x"87",
           442 => x"08",
           443 => x"51",
           444 => x"2e",
           445 => x"c0",
           446 => x"51",
           447 => x"87",
           448 => x"08",
           449 => x"06",
           450 => x"38",
           451 => x"8c",
           452 => x"80",
           453 => x"71",
           454 => x"9f",
           455 => x"0b",
           456 => x"33",
           457 => x"3d",
           458 => x"3d",
           459 => x"7d",
           460 => x"80",
           461 => x"0b",
           462 => x"81",
           463 => x"82",
           464 => x"2e",
           465 => x"81",
           466 => x"0b",
           467 => x"8c",
           468 => x"c0",
           469 => x"84",
           470 => x"92",
           471 => x"c0",
           472 => x"70",
           473 => x"81",
           474 => x"53",
           475 => x"a7",
           476 => x"92",
           477 => x"81",
           478 => x"79",
           479 => x"51",
           480 => x"90",
           481 => x"2e",
           482 => x"76",
           483 => x"58",
           484 => x"54",
           485 => x"72",
           486 => x"70",
           487 => x"38",
           488 => x"8c",
           489 => x"ff",
           490 => x"c0",
           491 => x"51",
           492 => x"81",
           493 => x"92",
           494 => x"c0",
           495 => x"70",
           496 => x"51",
           497 => x"80",
           498 => x"80",
           499 => x"70",
           500 => x"81",
           501 => x"87",
           502 => x"08",
           503 => x"2e",
           504 => x"83",
           505 => x"71",
           506 => x"3d",
           507 => x"3d",
           508 => x"11",
           509 => x"71",
           510 => x"88",
           511 => x"84",
           512 => x"fd",
           513 => x"83",
           514 => x"12",
           515 => x"2b",
           516 => x"07",
           517 => x"70",
           518 => x"2b",
           519 => x"07",
           520 => x"53",
           521 => x"52",
           522 => x"04",
           523 => x"79",
           524 => x"9f",
           525 => x"57",
           526 => x"80",
           527 => x"88",
           528 => x"80",
           529 => x"33",
           530 => x"2e",
           531 => x"83",
           532 => x"80",
           533 => x"54",
           534 => x"fe",
           535 => x"88",
           536 => x"08",
           537 => x"3d",
           538 => x"fd",
           539 => x"08",
           540 => x"51",
           541 => x"88",
           542 => x"ff",
           543 => x"39",
           544 => x"82",
           545 => x"06",
           546 => x"2a",
           547 => x"05",
           548 => x"70",
           549 => x"92",
           550 => x"8e",
           551 => x"fe",
           552 => x"08",
           553 => x"55",
           554 => x"55",
           555 => x"89",
           556 => x"fb",
           557 => x"0b",
           558 => x"08",
           559 => x"12",
           560 => x"55",
           561 => x"56",
           562 => x"8d",
           563 => x"33",
           564 => x"94",
           565 => x"57",
           566 => x"0c",
           567 => x"04",
           568 => x"75",
           569 => x"0b",
           570 => x"f4",
           571 => x"51",
           572 => x"83",
           573 => x"06",
           574 => x"14",
           575 => x"3f",
           576 => x"2b",
           577 => x"51",
           578 => x"88",
           579 => x"ff",
           580 => x"88",
           581 => x"0d",
           582 => x"0d",
           583 => x"0b",
           584 => x"55",
           585 => x"23",
           586 => x"53",
           587 => x"88",
           588 => x"08",
           589 => x"38",
           590 => x"39",
           591 => x"73",
           592 => x"83",
           593 => x"06",
           594 => x"14",
           595 => x"8c",
           596 => x"80",
           597 => x"72",
           598 => x"3f",
           599 => x"85",
           600 => x"08",
           601 => x"16",
           602 => x"71",
           603 => x"3d",
           604 => x"3d",
           605 => x"0b",
           606 => x"08",
           607 => x"05",
           608 => x"ff",
           609 => x"57",
           610 => x"2e",
           611 => x"15",
           612 => x"86",
           613 => x"80",
           614 => x"8f",
           615 => x"80",
           616 => x"13",
           617 => x"8c",
           618 => x"72",
           619 => x"0b",
           620 => x"57",
           621 => x"27",
           622 => x"39",
           623 => x"ff",
           624 => x"2a",
           625 => x"a8",
           626 => x"fc",
           627 => x"52",
           628 => x"27",
           629 => x"52",
           630 => x"17",
           631 => x"38",
           632 => x"16",
           633 => x"51",
           634 => x"88",
           635 => x"0c",
           636 => x"80",
           637 => x"0c",
           638 => x"04",
           639 => x"60",
           640 => x"5e",
           641 => x"55",
           642 => x"09",
           643 => x"38",
           644 => x"44",
           645 => x"62",
           646 => x"56",
           647 => x"09",
           648 => x"38",
           649 => x"80",
           650 => x"0c",
           651 => x"51",
           652 => x"26",
           653 => x"51",
           654 => x"88",
           655 => x"7d",
           656 => x"39",
           657 => x"1d",
           658 => x"5a",
           659 => x"a0",
           660 => x"05",
           661 => x"15",
           662 => x"2e",
           663 => x"ef",
           664 => x"59",
           665 => x"08",
           666 => x"81",
           667 => x"ff",
           668 => x"70",
           669 => x"32",
           670 => x"73",
           671 => x"25",
           672 => x"52",
           673 => x"57",
           674 => x"c7",
           675 => x"2e",
           676 => x"83",
           677 => x"77",
           678 => x"07",
           679 => x"2e",
           680 => x"88",
           681 => x"78",
           682 => x"30",
           683 => x"9f",
           684 => x"57",
           685 => x"9b",
           686 => x"8b",
           687 => x"39",
           688 => x"70",
           689 => x"72",
           690 => x"57",
           691 => x"34",
           692 => x"7a",
           693 => x"80",
           694 => x"26",
           695 => x"55",
           696 => x"34",
           697 => x"b1",
           698 => x"80",
           699 => x"54",
           700 => x"85",
           701 => x"06",
           702 => x"1c",
           703 => x"51",
           704 => x"88",
           705 => x"08",
           706 => x"7c",
           707 => x"80",
           708 => x"38",
           709 => x"70",
           710 => x"81",
           711 => x"56",
           712 => x"8b",
           713 => x"08",
           714 => x"5b",
           715 => x"18",
           716 => x"2e",
           717 => x"70",
           718 => x"33",
           719 => x"05",
           720 => x"71",
           721 => x"56",
           722 => x"e2",
           723 => x"75",
           724 => x"38",
           725 => x"9a",
           726 => x"39",
           727 => x"88",
           728 => x"83",
           729 => x"84",
           730 => x"11",
           731 => x"74",
           732 => x"1d",
           733 => x"2a",
           734 => x"51",
           735 => x"89",
           736 => x"92",
           737 => x"8e",
           738 => x"fa",
           739 => x"08",
           740 => x"fd",
           741 => x"88",
           742 => x"0d",
           743 => x"0d",
           744 => x"57",
           745 => x"fe",
           746 => x"76",
           747 => x"3f",
           748 => x"08",
           749 => x"76",
           750 => x"3f",
           751 => x"ff",
           752 => x"82",
           753 => x"d4",
           754 => x"81",
           755 => x"38",
           756 => x"53",
           757 => x"51",
           758 => x"88",
           759 => x"08",
           760 => x"51",
           761 => x"88",
           762 => x"ff",
           763 => x"81",
           764 => x"a9",
           765 => x"80",
           766 => x"52",
           767 => x"aa",
           768 => x"56",
           769 => x"38",
           770 => x"e2",
           771 => x"83",
           772 => x"55",
           773 => x"c6",
           774 => x"81",
           775 => x"0c",
           776 => x"04",
           777 => x"65",
           778 => x"0b",
           779 => x"f4",
           780 => x"3f",
           781 => x"06",
           782 => x"74",
           783 => x"74",
           784 => x"3d",
           785 => x"5a",
           786 => x"88",
           787 => x"06",
           788 => x"2e",
           789 => x"b3",
           790 => x"83",
           791 => x"52",
           792 => x"c6",
           793 => x"ab",
           794 => x"33",
           795 => x"2e",
           796 => x"3d",
           797 => x"f7",
           798 => x"08",
           799 => x"76",
           800 => x"99",
           801 => x"81",
           802 => x"76",
           803 => x"81",
           804 => x"81",
           805 => x"39",
           806 => x"86",
           807 => x"82",
           808 => x"54",
           809 => x"52",
           810 => x"fe",
           811 => x"88",
           812 => x"38",
           813 => x"05",
           814 => x"3f",
           815 => x"ff",
           816 => x"77",
           817 => x"3d",
           818 => x"f6",
           819 => x"08",
           820 => x"05",
           821 => x"29",
           822 => x"ad",
           823 => x"52",
           824 => x"8a",
           825 => x"83",
           826 => x"7a",
           827 => x"0c",
           828 => x"82",
           829 => x"3d",
           830 => x"f5",
           831 => x"08",
           832 => x"95",
           833 => x"51",
           834 => x"88",
           835 => x"ff",
           836 => x"8c",
           837 => x"ef",
           838 => x"e7",
           839 => x"56",
           840 => x"ca",
           841 => x"83",
           842 => x"76",
           843 => x"31",
           844 => x"70",
           845 => x"1d",
           846 => x"71",
           847 => x"5c",
           848 => x"c4",
           849 => x"82",
           850 => x"1b",
           851 => x"e0",
           852 => x"56",
           853 => x"fe",
           854 => x"82",
           855 => x"f6",
           856 => x"38",
           857 => x"39",
           858 => x"80",
           859 => x"38",
           860 => x"76",
           861 => x"81",
           862 => x"95",
           863 => x"51",
           864 => x"88",
           865 => x"0c",
           866 => x"19",
           867 => x"1a",
           868 => x"ff",
           869 => x"1a",
           870 => x"84",
           871 => x"1b",
           872 => x"0b",
           873 => x"78",
           874 => x"9f",
           875 => x"56",
           876 => x"95",
           877 => x"ea",
           878 => x"0b",
           879 => x"08",
           880 => x"74",
           881 => x"df",
           882 => x"81",
           883 => x"3d",
           884 => x"69",
           885 => x"70",
           886 => x"05",
           887 => x"3f",
           888 => x"88",
           889 => x"38",
           890 => x"54",
           891 => x"93",
           892 => x"05",
           893 => x"2a",
           894 => x"51",
           895 => x"80",
           896 => x"83",
           897 => x"75",
           898 => x"3f",
           899 => x"16",
           900 => x"dc",
           901 => x"eb",
           902 => x"9c",
           903 => x"98",
           904 => x"0b",
           905 => x"73",
           906 => x"3d",
           907 => x"3d",
           908 => x"7e",
           909 => x"9f",
           910 => x"5b",
           911 => x"7b",
           912 => x"75",
           913 => x"d1",
           914 => x"33",
           915 => x"84",
           916 => x"2e",
           917 => x"91",
           918 => x"17",
           919 => x"80",
           920 => x"34",
           921 => x"b1",
           922 => x"08",
           923 => x"31",
           924 => x"27",
           925 => x"58",
           926 => x"81",
           927 => x"16",
           928 => x"ff",
           929 => x"74",
           930 => x"82",
           931 => x"05",
           932 => x"06",
           933 => x"06",
           934 => x"9e",
           935 => x"38",
           936 => x"55",
           937 => x"16",
           938 => x"80",
           939 => x"55",
           940 => x"ff",
           941 => x"a4",
           942 => x"16",
           943 => x"f3",
           944 => x"55",
           945 => x"2e",
           946 => x"88",
           947 => x"17",
           948 => x"08",
           949 => x"84",
           950 => x"51",
           951 => x"27",
           952 => x"55",
           953 => x"16",
           954 => x"06",
           955 => x"08",
           956 => x"f0",
           957 => x"08",
           958 => x"98",
           959 => x"98",
           960 => x"75",
           961 => x"16",
           962 => x"78",
           963 => x"e8",
           964 => x"59",
           965 => x"80",
           966 => x"0c",
           967 => x"04",
           968 => x"87",
           969 => x"08",
           970 => x"80",
           971 => x"ea",
           972 => x"08",
           973 => x"c0",
           974 => x"56",
           975 => x"80",
           976 => x"ea",
           977 => x"88",
           978 => x"c0",
           979 => x"87",
           980 => x"08",
           981 => x"80",
           982 => x"ea",
           983 => x"08",
           984 => x"c0",
           985 => x"56",
           986 => x"80",
           987 => x"ea",
           988 => x"88",
           989 => x"c0",
           990 => x"8c",
           991 => x"87",
           992 => x"0c",
           993 => x"0b",
           994 => x"94",
           995 => x"51",
           996 => x"88",
           997 => x"9f",
           998 => x"9b",
           999 => x"ae",
          1000 => x"0b",
          1001 => x"c0",
          1002 => x"55",
          1003 => x"05",
          1004 => x"52",
          1005 => x"f6",
          1006 => x"8d",
          1007 => x"73",
          1008 => x"38",
          1009 => x"e4",
          1010 => x"54",
          1011 => x"54",
          1012 => x"00",
          1013 => x"ff",
          1014 => x"ff",
          1015 => x"ff",
          1016 => x"42",
          1017 => x"54",
          1018 => x"2e",
          1019 => x"00",
          1020 => x"01",
          2048 => x"0b",
          2049 => x"80",
          2050 => x"0b",
          2051 => x"ff",
          2052 => x"ff",
          2053 => x"ff",
          2054 => x"ff",
          2055 => x"ff",
          2056 => x"0b",
          2057 => x"80",
          2058 => x"0b",
          2059 => x"0b",
          2060 => x"93",
          2061 => x"0b",
          2062 => x"0b",
          2063 => x"b3",
          2064 => x"0b",
          2065 => x"0b",
          2066 => x"d3",
          2067 => x"0b",
          2068 => x"0b",
          2069 => x"f3",
          2070 => x"0b",
          2071 => x"0b",
          2072 => x"93",
          2073 => x"0b",
          2074 => x"0b",
          2075 => x"b3",
          2076 => x"0b",
          2077 => x"0b",
          2078 => x"d3",
          2079 => x"0b",
          2080 => x"0b",
          2081 => x"f1",
          2082 => x"0b",
          2083 => x"0b",
          2084 => x"8f",
          2085 => x"0b",
          2086 => x"0b",
          2087 => x"ae",
          2088 => x"0b",
          2089 => x"0b",
          2090 => x"ce",
          2091 => x"0b",
          2092 => x"0b",
          2093 => x"ee",
          2094 => x"0b",
          2095 => x"0b",
          2096 => x"8e",
          2097 => x"0b",
          2098 => x"0b",
          2099 => x"ae",
          2100 => x"0b",
          2101 => x"0b",
          2102 => x"ce",
          2103 => x"0b",
          2104 => x"0b",
          2105 => x"ee",
          2106 => x"0b",
          2107 => x"0b",
          2108 => x"8e",
          2109 => x"0b",
          2110 => x"0b",
          2111 => x"ae",
          2112 => x"0b",
          2113 => x"0b",
          2114 => x"ce",
          2115 => x"0b",
          2116 => x"0b",
          2117 => x"ee",
          2118 => x"0b",
          2119 => x"0b",
          2120 => x"8e",
          2121 => x"0b",
          2122 => x"0b",
          2123 => x"ae",
          2124 => x"0b",
          2125 => x"0b",
          2126 => x"ce",
          2127 => x"0b",
          2128 => x"0b",
          2129 => x"ee",
          2130 => x"0b",
          2131 => x"0b",
          2132 => x"8d",
          2133 => x"0b",
          2134 => x"0b",
          2135 => x"ab",
          2136 => x"00",
          2137 => x"00",
          2138 => x"00",
          2139 => x"00",
          2140 => x"00",
          2141 => x"00",
          2142 => x"00",
          2143 => x"00",
          2144 => x"00",
          2145 => x"00",
          2146 => x"00",
          2147 => x"00",
          2148 => x"00",
          2149 => x"00",
          2150 => x"00",
          2151 => x"00",
          2152 => x"00",
          2153 => x"00",
          2154 => x"00",
          2155 => x"00",
          2156 => x"00",
          2157 => x"00",
          2158 => x"00",
          2159 => x"00",
          2160 => x"00",
          2161 => x"00",
          2162 => x"00",
          2163 => x"00",
          2164 => x"00",
          2165 => x"00",
          2166 => x"00",
          2167 => x"00",
          2168 => x"00",
          2169 => x"00",
          2170 => x"00",
          2171 => x"00",
          2172 => x"00",
          2173 => x"00",
          2174 => x"00",
          2175 => x"00",
          2176 => x"00",
          2177 => x"82",
          2178 => x"b8",
          2179 => x"93",
          2180 => x"80",
          2181 => x"93",
          2182 => x"c9",
          2183 => x"93",
          2184 => x"80",
          2185 => x"93",
          2186 => x"ca",
          2187 => x"93",
          2188 => x"80",
          2189 => x"93",
          2190 => x"ca",
          2191 => x"93",
          2192 => x"80",
          2193 => x"93",
          2194 => x"d1",
          2195 => x"93",
          2196 => x"80",
          2197 => x"93",
          2198 => x"d2",
          2199 => x"93",
          2200 => x"80",
          2201 => x"93",
          2202 => x"ca",
          2203 => x"93",
          2204 => x"80",
          2205 => x"93",
          2206 => x"d2",
          2207 => x"93",
          2208 => x"80",
          2209 => x"93",
          2210 => x"d4",
          2211 => x"93",
          2212 => x"80",
          2213 => x"93",
          2214 => x"d0",
          2215 => x"93",
          2216 => x"80",
          2217 => x"93",
          2218 => x"cb",
          2219 => x"93",
          2220 => x"80",
          2221 => x"93",
          2222 => x"d0",
          2223 => x"93",
          2224 => x"80",
          2225 => x"93",
          2226 => x"d0",
          2227 => x"93",
          2228 => x"80",
          2229 => x"93",
          2230 => x"ad",
          2231 => x"90",
          2232 => x"90",
          2233 => x"90",
          2234 => x"2d",
          2235 => x"08",
          2236 => x"04",
          2237 => x"0c",
          2238 => x"82",
          2239 => x"83",
          2240 => x"82",
          2241 => x"b4",
          2242 => x"93",
          2243 => x"80",
          2244 => x"93",
          2245 => x"82",
          2246 => x"90",
          2247 => x"90",
          2248 => x"90",
          2249 => x"e6",
          2250 => x"90",
          2251 => x"90",
          2252 => x"90",
          2253 => x"d7",
          2254 => x"90",
          2255 => x"90",
          2256 => x"90",
          2257 => x"cb",
          2258 => x"90",
          2259 => x"90",
          2260 => x"90",
          2261 => x"c8",
          2262 => x"90",
          2263 => x"90",
          2264 => x"90",
          2265 => x"e6",
          2266 => x"90",
          2267 => x"90",
          2268 => x"90",
          2269 => x"c6",
          2270 => x"90",
          2271 => x"90",
          2272 => x"90",
          2273 => x"b9",
          2274 => x"90",
          2275 => x"90",
          2276 => x"90",
          2277 => x"85",
          2278 => x"90",
          2279 => x"90",
          2280 => x"90",
          2281 => x"a4",
          2282 => x"90",
          2283 => x"90",
          2284 => x"90",
          2285 => x"c3",
          2286 => x"90",
          2287 => x"90",
          2288 => x"90",
          2289 => x"ad",
          2290 => x"90",
          2291 => x"90",
          2292 => x"90",
          2293 => x"93",
          2294 => x"90",
          2295 => x"90",
          2296 => x"90",
          2297 => x"81",
          2298 => x"90",
          2299 => x"90",
          2300 => x"90",
          2301 => x"c7",
          2302 => x"90",
          2303 => x"90",
          2304 => x"90",
          2305 => x"81",
          2306 => x"90",
          2307 => x"90",
          2308 => x"90",
          2309 => x"82",
          2310 => x"90",
          2311 => x"90",
          2312 => x"90",
          2313 => x"b7",
          2314 => x"90",
          2315 => x"90",
          2316 => x"90",
          2317 => x"90",
          2318 => x"90",
          2319 => x"90",
          2320 => x"90",
          2321 => x"bb",
          2322 => x"90",
          2323 => x"90",
          2324 => x"90",
          2325 => x"9e",
          2326 => x"90",
          2327 => x"90",
          2328 => x"90",
          2329 => x"f3",
          2330 => x"90",
          2331 => x"90",
          2332 => x"90",
          2333 => x"fd",
          2334 => x"90",
          2335 => x"90",
          2336 => x"90",
          2337 => x"bf",
          2338 => x"90",
          2339 => x"90",
          2340 => x"90",
          2341 => x"85",
          2342 => x"90",
          2343 => x"90",
          2344 => x"90",
          2345 => x"ab",
          2346 => x"90",
          2347 => x"90",
          2348 => x"90",
          2349 => x"e0",
          2350 => x"90",
          2351 => x"90",
          2352 => x"90",
          2353 => x"cc",
          2354 => x"90",
          2355 => x"90",
          2356 => x"90",
          2357 => x"c0",
          2358 => x"90",
          2359 => x"90",
          2360 => x"90",
          2361 => x"aa",
          2362 => x"90",
          2363 => x"90",
          2364 => x"90",
          2365 => x"8e",
          2366 => x"90",
          2367 => x"90",
          2368 => x"90",
          2369 => x"2d",
          2370 => x"08",
          2371 => x"04",
          2372 => x"0c",
          2373 => x"82",
          2374 => x"83",
          2375 => x"82",
          2376 => x"b7",
          2377 => x"93",
          2378 => x"80",
          2379 => x"93",
          2380 => x"d6",
          2381 => x"93",
          2382 => x"80",
          2383 => x"93",
          2384 => x"aa",
          2385 => x"38",
          2386 => x"84",
          2387 => x"0b",
          2388 => x"be",
          2389 => x"51",
          2390 => x"04",
          2391 => x"93",
          2392 => x"82",
          2393 => x"fd",
          2394 => x"53",
          2395 => x"08",
          2396 => x"52",
          2397 => x"08",
          2398 => x"51",
          2399 => x"82",
          2400 => x"70",
          2401 => x"0c",
          2402 => x"0d",
          2403 => x"0c",
          2404 => x"90",
          2405 => x"93",
          2406 => x"3d",
          2407 => x"82",
          2408 => x"8c",
          2409 => x"82",
          2410 => x"88",
          2411 => x"93",
          2412 => x"84",
          2413 => x"93",
          2414 => x"85",
          2415 => x"93",
          2416 => x"82",
          2417 => x"02",
          2418 => x"0c",
          2419 => x"81",
          2420 => x"90",
          2421 => x"0c",
          2422 => x"93",
          2423 => x"05",
          2424 => x"90",
          2425 => x"08",
          2426 => x"08",
          2427 => x"27",
          2428 => x"93",
          2429 => x"05",
          2430 => x"ae",
          2431 => x"82",
          2432 => x"8c",
          2433 => x"a2",
          2434 => x"90",
          2435 => x"08",
          2436 => x"90",
          2437 => x"0c",
          2438 => x"08",
          2439 => x"10",
          2440 => x"08",
          2441 => x"ff",
          2442 => x"93",
          2443 => x"05",
          2444 => x"80",
          2445 => x"93",
          2446 => x"05",
          2447 => x"90",
          2448 => x"08",
          2449 => x"82",
          2450 => x"88",
          2451 => x"93",
          2452 => x"05",
          2453 => x"93",
          2454 => x"05",
          2455 => x"90",
          2456 => x"08",
          2457 => x"08",
          2458 => x"07",
          2459 => x"08",
          2460 => x"82",
          2461 => x"fc",
          2462 => x"2a",
          2463 => x"08",
          2464 => x"82",
          2465 => x"8c",
          2466 => x"2a",
          2467 => x"08",
          2468 => x"ff",
          2469 => x"93",
          2470 => x"05",
          2471 => x"93",
          2472 => x"90",
          2473 => x"08",
          2474 => x"90",
          2475 => x"0c",
          2476 => x"82",
          2477 => x"f8",
          2478 => x"82",
          2479 => x"f4",
          2480 => x"82",
          2481 => x"f4",
          2482 => x"93",
          2483 => x"3d",
          2484 => x"90",
          2485 => x"3d",
          2486 => x"79",
          2487 => x"55",
          2488 => x"27",
          2489 => x"75",
          2490 => x"51",
          2491 => x"a9",
          2492 => x"52",
          2493 => x"98",
          2494 => x"81",
          2495 => x"74",
          2496 => x"56",
          2497 => x"52",
          2498 => x"09",
          2499 => x"38",
          2500 => x"84",
          2501 => x"0d",
          2502 => x"72",
          2503 => x"54",
          2504 => x"84",
          2505 => x"72",
          2506 => x"54",
          2507 => x"84",
          2508 => x"72",
          2509 => x"54",
          2510 => x"84",
          2511 => x"72",
          2512 => x"54",
          2513 => x"84",
          2514 => x"f0",
          2515 => x"8f",
          2516 => x"83",
          2517 => x"38",
          2518 => x"05",
          2519 => x"70",
          2520 => x"0c",
          2521 => x"71",
          2522 => x"38",
          2523 => x"81",
          2524 => x"0d",
          2525 => x"02",
          2526 => x"05",
          2527 => x"53",
          2528 => x"27",
          2529 => x"83",
          2530 => x"80",
          2531 => x"ff",
          2532 => x"ff",
          2533 => x"73",
          2534 => x"05",
          2535 => x"12",
          2536 => x"2e",
          2537 => x"ef",
          2538 => x"93",
          2539 => x"3d",
          2540 => x"74",
          2541 => x"07",
          2542 => x"2b",
          2543 => x"51",
          2544 => x"a5",
          2545 => x"70",
          2546 => x"0c",
          2547 => x"84",
          2548 => x"72",
          2549 => x"05",
          2550 => x"71",
          2551 => x"53",
          2552 => x"52",
          2553 => x"dd",
          2554 => x"27",
          2555 => x"71",
          2556 => x"53",
          2557 => x"52",
          2558 => x"f2",
          2559 => x"ff",
          2560 => x"3d",
          2561 => x"79",
          2562 => x"83",
          2563 => x"54",
          2564 => x"c3",
          2565 => x"08",
          2566 => x"f7",
          2567 => x"13",
          2568 => x"84",
          2569 => x"06",
          2570 => x"53",
          2571 => x"38",
          2572 => x"74",
          2573 => x"56",
          2574 => x"70",
          2575 => x"fb",
          2576 => x"06",
          2577 => x"82",
          2578 => x"51",
          2579 => x"54",
          2580 => x"dc",
          2581 => x"71",
          2582 => x"53",
          2583 => x"73",
          2584 => x"55",
          2585 => x"38",
          2586 => x"84",
          2587 => x"0d",
          2588 => x"0d",
          2589 => x"83",
          2590 => x"52",
          2591 => x"71",
          2592 => x"09",
          2593 => x"ff",
          2594 => x"f8",
          2595 => x"80",
          2596 => x"52",
          2597 => x"38",
          2598 => x"08",
          2599 => x"fb",
          2600 => x"06",
          2601 => x"82",
          2602 => x"51",
          2603 => x"70",
          2604 => x"38",
          2605 => x"33",
          2606 => x"2e",
          2607 => x"12",
          2608 => x"52",
          2609 => x"71",
          2610 => x"93",
          2611 => x"3d",
          2612 => x"3d",
          2613 => x"7c",
          2614 => x"55",
          2615 => x"2e",
          2616 => x"71",
          2617 => x"06",
          2618 => x"2e",
          2619 => x"ff",
          2620 => x"ff",
          2621 => x"71",
          2622 => x"56",
          2623 => x"2e",
          2624 => x"a9",
          2625 => x"2e",
          2626 => x"70",
          2627 => x"51",
          2628 => x"80",
          2629 => x"12",
          2630 => x"15",
          2631 => x"72",
          2632 => x"81",
          2633 => x"71",
          2634 => x"56",
          2635 => x"ff",
          2636 => x"ff",
          2637 => x"31",
          2638 => x"70",
          2639 => x"0c",
          2640 => x"04",
          2641 => x"55",
          2642 => x"88",
          2643 => x"74",
          2644 => x"38",
          2645 => x"52",
          2646 => x"fc",
          2647 => x"80",
          2648 => x"74",
          2649 => x"f7",
          2650 => x"12",
          2651 => x"84",
          2652 => x"06",
          2653 => x"70",
          2654 => x"15",
          2655 => x"55",
          2656 => x"d0",
          2657 => x"76",
          2658 => x"38",
          2659 => x"52",
          2660 => x"80",
          2661 => x"84",
          2662 => x"0d",
          2663 => x"0d",
          2664 => x"53",
          2665 => x"52",
          2666 => x"82",
          2667 => x"81",
          2668 => x"07",
          2669 => x"52",
          2670 => x"e8",
          2671 => x"93",
          2672 => x"3d",
          2673 => x"3d",
          2674 => x"08",
          2675 => x"56",
          2676 => x"80",
          2677 => x"33",
          2678 => x"2e",
          2679 => x"86",
          2680 => x"52",
          2681 => x"53",
          2682 => x"13",
          2683 => x"33",
          2684 => x"06",
          2685 => x"70",
          2686 => x"38",
          2687 => x"80",
          2688 => x"74",
          2689 => x"81",
          2690 => x"70",
          2691 => x"81",
          2692 => x"80",
          2693 => x"05",
          2694 => x"76",
          2695 => x"70",
          2696 => x"0c",
          2697 => x"04",
          2698 => x"76",
          2699 => x"80",
          2700 => x"86",
          2701 => x"52",
          2702 => x"da",
          2703 => x"84",
          2704 => x"80",
          2705 => x"74",
          2706 => x"93",
          2707 => x"3d",
          2708 => x"3d",
          2709 => x"11",
          2710 => x"52",
          2711 => x"70",
          2712 => x"98",
          2713 => x"33",
          2714 => x"82",
          2715 => x"26",
          2716 => x"84",
          2717 => x"83",
          2718 => x"26",
          2719 => x"85",
          2720 => x"84",
          2721 => x"26",
          2722 => x"86",
          2723 => x"85",
          2724 => x"26",
          2725 => x"88",
          2726 => x"86",
          2727 => x"e7",
          2728 => x"38",
          2729 => x"54",
          2730 => x"87",
          2731 => x"cc",
          2732 => x"87",
          2733 => x"0c",
          2734 => x"c0",
          2735 => x"82",
          2736 => x"c0",
          2737 => x"83",
          2738 => x"c0",
          2739 => x"84",
          2740 => x"c0",
          2741 => x"85",
          2742 => x"c0",
          2743 => x"86",
          2744 => x"c0",
          2745 => x"74",
          2746 => x"a4",
          2747 => x"c0",
          2748 => x"80",
          2749 => x"98",
          2750 => x"52",
          2751 => x"84",
          2752 => x"0d",
          2753 => x"0d",
          2754 => x"c0",
          2755 => x"81",
          2756 => x"c0",
          2757 => x"5e",
          2758 => x"87",
          2759 => x"08",
          2760 => x"1c",
          2761 => x"98",
          2762 => x"79",
          2763 => x"87",
          2764 => x"08",
          2765 => x"1c",
          2766 => x"98",
          2767 => x"79",
          2768 => x"87",
          2769 => x"08",
          2770 => x"1c",
          2771 => x"98",
          2772 => x"7b",
          2773 => x"87",
          2774 => x"08",
          2775 => x"1c",
          2776 => x"0c",
          2777 => x"ff",
          2778 => x"83",
          2779 => x"58",
          2780 => x"57",
          2781 => x"56",
          2782 => x"55",
          2783 => x"54",
          2784 => x"53",
          2785 => x"ff",
          2786 => x"f6",
          2787 => x"9f",
          2788 => x"0d",
          2789 => x"0d",
          2790 => x"33",
          2791 => x"9f",
          2792 => x"52",
          2793 => x"82",
          2794 => x"83",
          2795 => x"fb",
          2796 => x"0b",
          2797 => x"fc",
          2798 => x"ff",
          2799 => x"56",
          2800 => x"84",
          2801 => x"2e",
          2802 => x"c0",
          2803 => x"70",
          2804 => x"2a",
          2805 => x"53",
          2806 => x"80",
          2807 => x"71",
          2808 => x"81",
          2809 => x"70",
          2810 => x"81",
          2811 => x"06",
          2812 => x"80",
          2813 => x"71",
          2814 => x"81",
          2815 => x"70",
          2816 => x"73",
          2817 => x"51",
          2818 => x"80",
          2819 => x"2e",
          2820 => x"c0",
          2821 => x"75",
          2822 => x"82",
          2823 => x"87",
          2824 => x"fb",
          2825 => x"9f",
          2826 => x"0b",
          2827 => x"33",
          2828 => x"06",
          2829 => x"87",
          2830 => x"51",
          2831 => x"86",
          2832 => x"94",
          2833 => x"08",
          2834 => x"70",
          2835 => x"54",
          2836 => x"2e",
          2837 => x"91",
          2838 => x"06",
          2839 => x"d7",
          2840 => x"32",
          2841 => x"51",
          2842 => x"2e",
          2843 => x"93",
          2844 => x"06",
          2845 => x"ff",
          2846 => x"81",
          2847 => x"87",
          2848 => x"52",
          2849 => x"86",
          2850 => x"94",
          2851 => x"72",
          2852 => x"0d",
          2853 => x"0d",
          2854 => x"74",
          2855 => x"ff",
          2856 => x"57",
          2857 => x"80",
          2858 => x"81",
          2859 => x"15",
          2860 => x"8d",
          2861 => x"81",
          2862 => x"57",
          2863 => x"c0",
          2864 => x"75",
          2865 => x"38",
          2866 => x"94",
          2867 => x"70",
          2868 => x"81",
          2869 => x"52",
          2870 => x"8c",
          2871 => x"2a",
          2872 => x"51",
          2873 => x"38",
          2874 => x"70",
          2875 => x"51",
          2876 => x"8d",
          2877 => x"2a",
          2878 => x"51",
          2879 => x"be",
          2880 => x"ff",
          2881 => x"c0",
          2882 => x"70",
          2883 => x"38",
          2884 => x"90",
          2885 => x"0c",
          2886 => x"33",
          2887 => x"06",
          2888 => x"70",
          2889 => x"76",
          2890 => x"0c",
          2891 => x"04",
          2892 => x"0b",
          2893 => x"fc",
          2894 => x"ff",
          2895 => x"87",
          2896 => x"51",
          2897 => x"86",
          2898 => x"94",
          2899 => x"08",
          2900 => x"70",
          2901 => x"51",
          2902 => x"2e",
          2903 => x"81",
          2904 => x"87",
          2905 => x"52",
          2906 => x"86",
          2907 => x"94",
          2908 => x"08",
          2909 => x"06",
          2910 => x"0c",
          2911 => x"0d",
          2912 => x"0d",
          2913 => x"8d",
          2914 => x"81",
          2915 => x"53",
          2916 => x"84",
          2917 => x"2e",
          2918 => x"c0",
          2919 => x"71",
          2920 => x"2a",
          2921 => x"51",
          2922 => x"52",
          2923 => x"a0",
          2924 => x"ff",
          2925 => x"c0",
          2926 => x"70",
          2927 => x"38",
          2928 => x"90",
          2929 => x"70",
          2930 => x"98",
          2931 => x"51",
          2932 => x"84",
          2933 => x"0d",
          2934 => x"0d",
          2935 => x"80",
          2936 => x"2a",
          2937 => x"51",
          2938 => x"84",
          2939 => x"c0",
          2940 => x"82",
          2941 => x"87",
          2942 => x"08",
          2943 => x"0c",
          2944 => x"94",
          2945 => x"88",
          2946 => x"9e",
          2947 => x"8e",
          2948 => x"c0",
          2949 => x"82",
          2950 => x"87",
          2951 => x"08",
          2952 => x"0c",
          2953 => x"ac",
          2954 => x"98",
          2955 => x"9e",
          2956 => x"8e",
          2957 => x"c0",
          2958 => x"82",
          2959 => x"87",
          2960 => x"08",
          2961 => x"0c",
          2962 => x"bc",
          2963 => x"a8",
          2964 => x"9e",
          2965 => x"8e",
          2966 => x"c0",
          2967 => x"82",
          2968 => x"87",
          2969 => x"08",
          2970 => x"8e",
          2971 => x"c0",
          2972 => x"82",
          2973 => x"87",
          2974 => x"08",
          2975 => x"0c",
          2976 => x"8c",
          2977 => x"c0",
          2978 => x"82",
          2979 => x"80",
          2980 => x"9e",
          2981 => x"84",
          2982 => x"51",
          2983 => x"80",
          2984 => x"81",
          2985 => x"8e",
          2986 => x"0b",
          2987 => x"90",
          2988 => x"80",
          2989 => x"52",
          2990 => x"2e",
          2991 => x"52",
          2992 => x"c6",
          2993 => x"87",
          2994 => x"08",
          2995 => x"0a",
          2996 => x"52",
          2997 => x"83",
          2998 => x"71",
          2999 => x"34",
          3000 => x"c0",
          3001 => x"70",
          3002 => x"06",
          3003 => x"70",
          3004 => x"38",
          3005 => x"82",
          3006 => x"80",
          3007 => x"9e",
          3008 => x"a0",
          3009 => x"51",
          3010 => x"80",
          3011 => x"81",
          3012 => x"8e",
          3013 => x"0b",
          3014 => x"90",
          3015 => x"80",
          3016 => x"52",
          3017 => x"2e",
          3018 => x"52",
          3019 => x"ca",
          3020 => x"87",
          3021 => x"08",
          3022 => x"80",
          3023 => x"52",
          3024 => x"83",
          3025 => x"71",
          3026 => x"34",
          3027 => x"c0",
          3028 => x"70",
          3029 => x"06",
          3030 => x"70",
          3031 => x"38",
          3032 => x"82",
          3033 => x"80",
          3034 => x"9e",
          3035 => x"81",
          3036 => x"51",
          3037 => x"80",
          3038 => x"81",
          3039 => x"8e",
          3040 => x"0b",
          3041 => x"90",
          3042 => x"c0",
          3043 => x"52",
          3044 => x"2e",
          3045 => x"52",
          3046 => x"ce",
          3047 => x"87",
          3048 => x"08",
          3049 => x"06",
          3050 => x"70",
          3051 => x"38",
          3052 => x"82",
          3053 => x"87",
          3054 => x"08",
          3055 => x"06",
          3056 => x"51",
          3057 => x"82",
          3058 => x"80",
          3059 => x"9e",
          3060 => x"84",
          3061 => x"52",
          3062 => x"2e",
          3063 => x"52",
          3064 => x"d1",
          3065 => x"9e",
          3066 => x"83",
          3067 => x"84",
          3068 => x"51",
          3069 => x"d2",
          3070 => x"87",
          3071 => x"08",
          3072 => x"51",
          3073 => x"80",
          3074 => x"81",
          3075 => x"8e",
          3076 => x"c0",
          3077 => x"70",
          3078 => x"51",
          3079 => x"d4",
          3080 => x"0d",
          3081 => x"0d",
          3082 => x"51",
          3083 => x"82",
          3084 => x"54",
          3085 => x"88",
          3086 => x"94",
          3087 => x"3f",
          3088 => x"51",
          3089 => x"82",
          3090 => x"54",
          3091 => x"93",
          3092 => x"a0",
          3093 => x"a4",
          3094 => x"52",
          3095 => x"51",
          3096 => x"82",
          3097 => x"54",
          3098 => x"93",
          3099 => x"98",
          3100 => x"9c",
          3101 => x"52",
          3102 => x"51",
          3103 => x"82",
          3104 => x"54",
          3105 => x"93",
          3106 => x"80",
          3107 => x"84",
          3108 => x"52",
          3109 => x"51",
          3110 => x"82",
          3111 => x"54",
          3112 => x"93",
          3113 => x"88",
          3114 => x"8c",
          3115 => x"52",
          3116 => x"51",
          3117 => x"82",
          3118 => x"54",
          3119 => x"93",
          3120 => x"90",
          3121 => x"94",
          3122 => x"52",
          3123 => x"51",
          3124 => x"82",
          3125 => x"54",
          3126 => x"8d",
          3127 => x"d0",
          3128 => x"f8",
          3129 => x"c7",
          3130 => x"d3",
          3131 => x"80",
          3132 => x"82",
          3133 => x"52",
          3134 => x"51",
          3135 => x"82",
          3136 => x"54",
          3137 => x"8d",
          3138 => x"d2",
          3139 => x"f9",
          3140 => x"9b",
          3141 => x"c5",
          3142 => x"80",
          3143 => x"81",
          3144 => x"88",
          3145 => x"8e",
          3146 => x"73",
          3147 => x"38",
          3148 => x"51",
          3149 => x"82",
          3150 => x"54",
          3151 => x"88",
          3152 => x"cc",
          3153 => x"3f",
          3154 => x"33",
          3155 => x"2e",
          3156 => x"f9",
          3157 => x"f3",
          3158 => x"ce",
          3159 => x"80",
          3160 => x"81",
          3161 => x"87",
          3162 => x"f9",
          3163 => x"db",
          3164 => x"a8",
          3165 => x"f9",
          3166 => x"b3",
          3167 => x"ac",
          3168 => x"fa",
          3169 => x"a7",
          3170 => x"b0",
          3171 => x"fa",
          3172 => x"9b",
          3173 => x"f4",
          3174 => x"3f",
          3175 => x"22",
          3176 => x"fc",
          3177 => x"3f",
          3178 => x"08",
          3179 => x"c0",
          3180 => x"e7",
          3181 => x"93",
          3182 => x"84",
          3183 => x"71",
          3184 => x"82",
          3185 => x"52",
          3186 => x"51",
          3187 => x"82",
          3188 => x"54",
          3189 => x"a8",
          3190 => x"bc",
          3191 => x"84",
          3192 => x"51",
          3193 => x"82",
          3194 => x"bd",
          3195 => x"76",
          3196 => x"54",
          3197 => x"08",
          3198 => x"d0",
          3199 => x"3f",
          3200 => x"33",
          3201 => x"2e",
          3202 => x"8e",
          3203 => x"bd",
          3204 => x"75",
          3205 => x"3f",
          3206 => x"08",
          3207 => x"29",
          3208 => x"54",
          3209 => x"84",
          3210 => x"fb",
          3211 => x"ff",
          3212 => x"f8",
          3213 => x"3f",
          3214 => x"04",
          3215 => x"02",
          3216 => x"ff",
          3217 => x"84",
          3218 => x"71",
          3219 => x"0b",
          3220 => x"05",
          3221 => x"04",
          3222 => x"51",
          3223 => x"fc",
          3224 => x"39",
          3225 => x"51",
          3226 => x"fc",
          3227 => x"39",
          3228 => x"51",
          3229 => x"fc",
          3230 => x"cf",
          3231 => x"0d",
          3232 => x"80",
          3233 => x"3d",
          3234 => x"96",
          3235 => x"52",
          3236 => x"0c",
          3237 => x"70",
          3238 => x"0c",
          3239 => x"3d",
          3240 => x"3d",
          3241 => x"96",
          3242 => x"82",
          3243 => x"52",
          3244 => x"73",
          3245 => x"8e",
          3246 => x"70",
          3247 => x"0c",
          3248 => x"83",
          3249 => x"80",
          3250 => x"96",
          3251 => x"82",
          3252 => x"87",
          3253 => x"0c",
          3254 => x"0d",
          3255 => x"08",
          3256 => x"aa",
          3257 => x"93",
          3258 => x"93",
          3259 => x"11",
          3260 => x"53",
          3261 => x"f8",
          3262 => x"70",
          3263 => x"0c",
          3264 => x"82",
          3265 => x"84",
          3266 => x"f9",
          3267 => x"7b",
          3268 => x"a0",
          3269 => x"08",
          3270 => x"90",
          3271 => x"58",
          3272 => x"53",
          3273 => x"ba",
          3274 => x"88",
          3275 => x"51",
          3276 => x"76",
          3277 => x"12",
          3278 => x"0c",
          3279 => x"0c",
          3280 => x"0c",
          3281 => x"0c",
          3282 => x"0c",
          3283 => x"0c",
          3284 => x"0c",
          3285 => x"0c",
          3286 => x"0c",
          3287 => x"0c",
          3288 => x"73",
          3289 => x"16",
          3290 => x"15",
          3291 => x"93",
          3292 => x"3d",
          3293 => x"3d",
          3294 => x"11",
          3295 => x"08",
          3296 => x"71",
          3297 => x"09",
          3298 => x"38",
          3299 => x"70",
          3300 => x"70",
          3301 => x"81",
          3302 => x"84",
          3303 => x"84",
          3304 => x"88",
          3305 => x"8c",
          3306 => x"53",
          3307 => x"73",
          3308 => x"ec",
          3309 => x"0c",
          3310 => x"0b",
          3311 => x"72",
          3312 => x"0c",
          3313 => x"73",
          3314 => x"51",
          3315 => x"2e",
          3316 => x"b3",
          3317 => x"08",
          3318 => x"52",
          3319 => x"09",
          3320 => x"38",
          3321 => x"12",
          3322 => x"94",
          3323 => x"15",
          3324 => x"13",
          3325 => x"12",
          3326 => x"08",
          3327 => x"70",
          3328 => x"52",
          3329 => x"72",
          3330 => x"0c",
          3331 => x"04",
          3332 => x"79",
          3333 => x"76",
          3334 => x"b5",
          3335 => x"f0",
          3336 => x"ec",
          3337 => x"75",
          3338 => x"8f",
          3339 => x"08",
          3340 => x"c7",
          3341 => x"08",
          3342 => x"83",
          3343 => x"fc",
          3344 => x"70",
          3345 => x"91",
          3346 => x"84",
          3347 => x"84",
          3348 => x"82",
          3349 => x"07",
          3350 => x"93",
          3351 => x"70",
          3352 => x"07",
          3353 => x"07",
          3354 => x"51",
          3355 => x"54",
          3356 => x"09",
          3357 => x"d9",
          3358 => x"76",
          3359 => x"80",
          3360 => x"0b",
          3361 => x"08",
          3362 => x"93",
          3363 => x"05",
          3364 => x"e8",
          3365 => x"08",
          3366 => x"38",
          3367 => x"87",
          3368 => x"08",
          3369 => x"88",
          3370 => x"17",
          3371 => x"17",
          3372 => x"14",
          3373 => x"08",
          3374 => x"0c",
          3375 => x"fd",
          3376 => x"52",
          3377 => x"08",
          3378 => x"3f",
          3379 => x"08",
          3380 => x"93",
          3381 => x"3d",
          3382 => x"3d",
          3383 => x"71",
          3384 => x"38",
          3385 => x"fd",
          3386 => x"3d",
          3387 => x"3d",
          3388 => x"05",
          3389 => x"8a",
          3390 => x"06",
          3391 => x"51",
          3392 => x"93",
          3393 => x"71",
          3394 => x"38",
          3395 => x"82",
          3396 => x"81",
          3397 => x"a0",
          3398 => x"82",
          3399 => x"52",
          3400 => x"85",
          3401 => x"71",
          3402 => x"0d",
          3403 => x"0d",
          3404 => x"33",
          3405 => x"08",
          3406 => x"98",
          3407 => x"ff",
          3408 => x"82",
          3409 => x"84",
          3410 => x"fd",
          3411 => x"54",
          3412 => x"81",
          3413 => x"53",
          3414 => x"8e",
          3415 => x"ff",
          3416 => x"14",
          3417 => x"3f",
          3418 => x"3d",
          3419 => x"3d",
          3420 => x"93",
          3421 => x"82",
          3422 => x"56",
          3423 => x"70",
          3424 => x"53",
          3425 => x"2e",
          3426 => x"81",
          3427 => x"81",
          3428 => x"da",
          3429 => x"74",
          3430 => x"0c",
          3431 => x"04",
          3432 => x"66",
          3433 => x"78",
          3434 => x"5a",
          3435 => x"80",
          3436 => x"38",
          3437 => x"09",
          3438 => x"de",
          3439 => x"7a",
          3440 => x"5c",
          3441 => x"5b",
          3442 => x"09",
          3443 => x"38",
          3444 => x"39",
          3445 => x"09",
          3446 => x"38",
          3447 => x"70",
          3448 => x"33",
          3449 => x"2e",
          3450 => x"92",
          3451 => x"19",
          3452 => x"70",
          3453 => x"33",
          3454 => x"53",
          3455 => x"16",
          3456 => x"26",
          3457 => x"88",
          3458 => x"05",
          3459 => x"05",
          3460 => x"05",
          3461 => x"5b",
          3462 => x"80",
          3463 => x"30",
          3464 => x"80",
          3465 => x"cc",
          3466 => x"70",
          3467 => x"25",
          3468 => x"54",
          3469 => x"53",
          3470 => x"8c",
          3471 => x"07",
          3472 => x"05",
          3473 => x"5a",
          3474 => x"83",
          3475 => x"54",
          3476 => x"27",
          3477 => x"16",
          3478 => x"06",
          3479 => x"80",
          3480 => x"aa",
          3481 => x"cf",
          3482 => x"73",
          3483 => x"81",
          3484 => x"80",
          3485 => x"38",
          3486 => x"2e",
          3487 => x"81",
          3488 => x"80",
          3489 => x"8a",
          3490 => x"39",
          3491 => x"2e",
          3492 => x"73",
          3493 => x"8a",
          3494 => x"d3",
          3495 => x"80",
          3496 => x"80",
          3497 => x"ee",
          3498 => x"39",
          3499 => x"71",
          3500 => x"53",
          3501 => x"54",
          3502 => x"2e",
          3503 => x"15",
          3504 => x"33",
          3505 => x"72",
          3506 => x"81",
          3507 => x"39",
          3508 => x"56",
          3509 => x"27",
          3510 => x"51",
          3511 => x"75",
          3512 => x"72",
          3513 => x"38",
          3514 => x"df",
          3515 => x"16",
          3516 => x"7b",
          3517 => x"38",
          3518 => x"f2",
          3519 => x"77",
          3520 => x"12",
          3521 => x"53",
          3522 => x"5c",
          3523 => x"5c",
          3524 => x"5c",
          3525 => x"5c",
          3526 => x"51",
          3527 => x"fd",
          3528 => x"82",
          3529 => x"06",
          3530 => x"80",
          3531 => x"77",
          3532 => x"53",
          3533 => x"18",
          3534 => x"72",
          3535 => x"c4",
          3536 => x"70",
          3537 => x"25",
          3538 => x"55",
          3539 => x"8d",
          3540 => x"2e",
          3541 => x"30",
          3542 => x"5b",
          3543 => x"8f",
          3544 => x"7b",
          3545 => x"dc",
          3546 => x"93",
          3547 => x"ff",
          3548 => x"75",
          3549 => x"e6",
          3550 => x"84",
          3551 => x"74",
          3552 => x"a7",
          3553 => x"80",
          3554 => x"38",
          3555 => x"72",
          3556 => x"54",
          3557 => x"72",
          3558 => x"05",
          3559 => x"17",
          3560 => x"77",
          3561 => x"51",
          3562 => x"9f",
          3563 => x"72",
          3564 => x"79",
          3565 => x"81",
          3566 => x"72",
          3567 => x"38",
          3568 => x"05",
          3569 => x"ad",
          3570 => x"17",
          3571 => x"81",
          3572 => x"b0",
          3573 => x"38",
          3574 => x"81",
          3575 => x"06",
          3576 => x"9f",
          3577 => x"55",
          3578 => x"97",
          3579 => x"f9",
          3580 => x"81",
          3581 => x"8b",
          3582 => x"16",
          3583 => x"73",
          3584 => x"96",
          3585 => x"e0",
          3586 => x"17",
          3587 => x"33",
          3588 => x"f9",
          3589 => x"f2",
          3590 => x"16",
          3591 => x"7b",
          3592 => x"38",
          3593 => x"c6",
          3594 => x"96",
          3595 => x"fd",
          3596 => x"3d",
          3597 => x"05",
          3598 => x"52",
          3599 => x"e0",
          3600 => x"0d",
          3601 => x"0d",
          3602 => x"a0",
          3603 => x"88",
          3604 => x"51",
          3605 => x"82",
          3606 => x"53",
          3607 => x"80",
          3608 => x"a0",
          3609 => x"0d",
          3610 => x"0d",
          3611 => x"08",
          3612 => x"98",
          3613 => x"88",
          3614 => x"52",
          3615 => x"3f",
          3616 => x"98",
          3617 => x"0d",
          3618 => x"0d",
          3619 => x"93",
          3620 => x"56",
          3621 => x"80",
          3622 => x"2e",
          3623 => x"82",
          3624 => x"52",
          3625 => x"93",
          3626 => x"ff",
          3627 => x"80",
          3628 => x"38",
          3629 => x"b9",
          3630 => x"32",
          3631 => x"80",
          3632 => x"52",
          3633 => x"8b",
          3634 => x"2e",
          3635 => x"14",
          3636 => x"9f",
          3637 => x"38",
          3638 => x"73",
          3639 => x"38",
          3640 => x"72",
          3641 => x"14",
          3642 => x"f8",
          3643 => x"af",
          3644 => x"52",
          3645 => x"8a",
          3646 => x"3f",
          3647 => x"82",
          3648 => x"87",
          3649 => x"fe",
          3650 => x"93",
          3651 => x"82",
          3652 => x"77",
          3653 => x"53",
          3654 => x"72",
          3655 => x"0c",
          3656 => x"04",
          3657 => x"7a",
          3658 => x"80",
          3659 => x"58",
          3660 => x"33",
          3661 => x"a0",
          3662 => x"06",
          3663 => x"13",
          3664 => x"39",
          3665 => x"09",
          3666 => x"38",
          3667 => x"11",
          3668 => x"08",
          3669 => x"54",
          3670 => x"2e",
          3671 => x"80",
          3672 => x"08",
          3673 => x"0c",
          3674 => x"33",
          3675 => x"80",
          3676 => x"38",
          3677 => x"80",
          3678 => x"38",
          3679 => x"57",
          3680 => x"0c",
          3681 => x"33",
          3682 => x"39",
          3683 => x"74",
          3684 => x"38",
          3685 => x"80",
          3686 => x"89",
          3687 => x"38",
          3688 => x"d0",
          3689 => x"55",
          3690 => x"80",
          3691 => x"39",
          3692 => x"d9",
          3693 => x"80",
          3694 => x"27",
          3695 => x"80",
          3696 => x"89",
          3697 => x"70",
          3698 => x"55",
          3699 => x"70",
          3700 => x"55",
          3701 => x"27",
          3702 => x"14",
          3703 => x"06",
          3704 => x"74",
          3705 => x"73",
          3706 => x"38",
          3707 => x"14",
          3708 => x"05",
          3709 => x"08",
          3710 => x"54",
          3711 => x"39",
          3712 => x"84",
          3713 => x"55",
          3714 => x"81",
          3715 => x"93",
          3716 => x"3d",
          3717 => x"3d",
          3718 => x"5a",
          3719 => x"7a",
          3720 => x"08",
          3721 => x"53",
          3722 => x"09",
          3723 => x"38",
          3724 => x"0c",
          3725 => x"ad",
          3726 => x"06",
          3727 => x"76",
          3728 => x"0c",
          3729 => x"33",
          3730 => x"73",
          3731 => x"81",
          3732 => x"38",
          3733 => x"05",
          3734 => x"08",
          3735 => x"53",
          3736 => x"2e",
          3737 => x"57",
          3738 => x"2e",
          3739 => x"39",
          3740 => x"13",
          3741 => x"08",
          3742 => x"53",
          3743 => x"55",
          3744 => x"80",
          3745 => x"14",
          3746 => x"88",
          3747 => x"27",
          3748 => x"eb",
          3749 => x"53",
          3750 => x"89",
          3751 => x"38",
          3752 => x"55",
          3753 => x"8a",
          3754 => x"a0",
          3755 => x"c2",
          3756 => x"74",
          3757 => x"e0",
          3758 => x"ff",
          3759 => x"d0",
          3760 => x"ff",
          3761 => x"90",
          3762 => x"38",
          3763 => x"81",
          3764 => x"53",
          3765 => x"ca",
          3766 => x"27",
          3767 => x"77",
          3768 => x"08",
          3769 => x"0c",
          3770 => x"33",
          3771 => x"ff",
          3772 => x"80",
          3773 => x"74",
          3774 => x"79",
          3775 => x"74",
          3776 => x"0c",
          3777 => x"04",
          3778 => x"76",
          3779 => x"98",
          3780 => x"2b",
          3781 => x"72",
          3782 => x"82",
          3783 => x"51",
          3784 => x"80",
          3785 => x"e0",
          3786 => x"53",
          3787 => x"9c",
          3788 => x"dc",
          3789 => x"02",
          3790 => x"05",
          3791 => x"52",
          3792 => x"72",
          3793 => x"06",
          3794 => x"53",
          3795 => x"84",
          3796 => x"0d",
          3797 => x"0d",
          3798 => x"05",
          3799 => x"71",
          3800 => x"53",
          3801 => x"9f",
          3802 => x"f3",
          3803 => x"51",
          3804 => x"88",
          3805 => x"3f",
          3806 => x"05",
          3807 => x"34",
          3808 => x"06",
          3809 => x"76",
          3810 => x"3f",
          3811 => x"86",
          3812 => x"f6",
          3813 => x"02",
          3814 => x"05",
          3815 => x"05",
          3816 => x"82",
          3817 => x"70",
          3818 => x"8e",
          3819 => x"08",
          3820 => x"5a",
          3821 => x"80",
          3822 => x"74",
          3823 => x"3f",
          3824 => x"33",
          3825 => x"82",
          3826 => x"81",
          3827 => x"58",
          3828 => x"bc",
          3829 => x"84",
          3830 => x"82",
          3831 => x"70",
          3832 => x"8e",
          3833 => x"08",
          3834 => x"74",
          3835 => x"38",
          3836 => x"52",
          3837 => x"de",
          3838 => x"d0",
          3839 => x"55",
          3840 => x"d0",
          3841 => x"ff",
          3842 => x"75",
          3843 => x"80",
          3844 => x"d0",
          3845 => x"2e",
          3846 => x"8f",
          3847 => x"75",
          3848 => x"38",
          3849 => x"33",
          3850 => x"38",
          3851 => x"05",
          3852 => x"78",
          3853 => x"80",
          3854 => x"82",
          3855 => x"52",
          3856 => x"fd",
          3857 => x"8f",
          3858 => x"80",
          3859 => x"8c",
          3860 => x"dc",
          3861 => x"57",
          3862 => x"8f",
          3863 => x"80",
          3864 => x"82",
          3865 => x"80",
          3866 => x"8f",
          3867 => x"80",
          3868 => x"3d",
          3869 => x"80",
          3870 => x"82",
          3871 => x"80",
          3872 => x"75",
          3873 => x"3f",
          3874 => x"08",
          3875 => x"82",
          3876 => x"25",
          3877 => x"93",
          3878 => x"05",
          3879 => x"55",
          3880 => x"75",
          3881 => x"81",
          3882 => x"f4",
          3883 => x"ff",
          3884 => x"2e",
          3885 => x"ff",
          3886 => x"3d",
          3887 => x"3d",
          3888 => x"08",
          3889 => x"5a",
          3890 => x"58",
          3891 => x"82",
          3892 => x"51",
          3893 => x"3f",
          3894 => x"08",
          3895 => x"ff",
          3896 => x"cc",
          3897 => x"80",
          3898 => x"3d",
          3899 => x"80",
          3900 => x"82",
          3901 => x"80",
          3902 => x"75",
          3903 => x"3f",
          3904 => x"08",
          3905 => x"55",
          3906 => x"93",
          3907 => x"8e",
          3908 => x"84",
          3909 => x"70",
          3910 => x"80",
          3911 => x"09",
          3912 => x"72",
          3913 => x"51",
          3914 => x"77",
          3915 => x"73",
          3916 => x"82",
          3917 => x"8c",
          3918 => x"51",
          3919 => x"3f",
          3920 => x"08",
          3921 => x"38",
          3922 => x"51",
          3923 => x"78",
          3924 => x"81",
          3925 => x"75",
          3926 => x"d5",
          3927 => x"51",
          3928 => x"ab",
          3929 => x"82",
          3930 => x"74",
          3931 => x"77",
          3932 => x"0c",
          3933 => x"04",
          3934 => x"7c",
          3935 => x"71",
          3936 => x"59",
          3937 => x"a0",
          3938 => x"06",
          3939 => x"33",
          3940 => x"77",
          3941 => x"38",
          3942 => x"5b",
          3943 => x"56",
          3944 => x"a0",
          3945 => x"06",
          3946 => x"75",
          3947 => x"80",
          3948 => x"29",
          3949 => x"05",
          3950 => x"55",
          3951 => x"82",
          3952 => x"53",
          3953 => x"08",
          3954 => x"3f",
          3955 => x"08",
          3956 => x"84",
          3957 => x"74",
          3958 => x"38",
          3959 => x"88",
          3960 => x"fc",
          3961 => x"39",
          3962 => x"8c",
          3963 => x"53",
          3964 => x"f6",
          3965 => x"93",
          3966 => x"2e",
          3967 => x"53",
          3968 => x"51",
          3969 => x"82",
          3970 => x"81",
          3971 => x"74",
          3972 => x"54",
          3973 => x"14",
          3974 => x"06",
          3975 => x"74",
          3976 => x"38",
          3977 => x"82",
          3978 => x"8c",
          3979 => x"d3",
          3980 => x"3d",
          3981 => x"05",
          3982 => x"33",
          3983 => x"0b",
          3984 => x"82",
          3985 => x"5b",
          3986 => x"08",
          3987 => x"82",
          3988 => x"54",
          3989 => x"38",
          3990 => x"b4",
          3991 => x"84",
          3992 => x"cc",
          3993 => x"84",
          3994 => x"80",
          3995 => x"53",
          3996 => x"08",
          3997 => x"84",
          3998 => x"ed",
          3999 => x"84",
          4000 => x"8b",
          4001 => x"ac",
          4002 => x"3f",
          4003 => x"82",
          4004 => x"53",
          4005 => x"90",
          4006 => x"54",
          4007 => x"3f",
          4008 => x"08",
          4009 => x"84",
          4010 => x"09",
          4011 => x"c1",
          4012 => x"84",
          4013 => x"b9",
          4014 => x"84",
          4015 => x"0b",
          4016 => x"08",
          4017 => x"82",
          4018 => x"ff",
          4019 => x"55",
          4020 => x"34",
          4021 => x"81",
          4022 => x"75",
          4023 => x"3f",
          4024 => x"09",
          4025 => x"a7",
          4026 => x"81",
          4027 => x"c8",
          4028 => x"5d",
          4029 => x"82",
          4030 => x"98",
          4031 => x"2c",
          4032 => x"ff",
          4033 => x"78",
          4034 => x"82",
          4035 => x"70",
          4036 => x"98",
          4037 => x"a4",
          4038 => x"2b",
          4039 => x"71",
          4040 => x"70",
          4041 => x"fd",
          4042 => x"08",
          4043 => x"51",
          4044 => x"59",
          4045 => x"5d",
          4046 => x"73",
          4047 => x"e9",
          4048 => x"27",
          4049 => x"81",
          4050 => x"81",
          4051 => x"70",
          4052 => x"55",
          4053 => x"80",
          4054 => x"53",
          4055 => x"51",
          4056 => x"82",
          4057 => x"81",
          4058 => x"73",
          4059 => x"38",
          4060 => x"a4",
          4061 => x"b1",
          4062 => x"80",
          4063 => x"80",
          4064 => x"98",
          4065 => x"ff",
          4066 => x"55",
          4067 => x"97",
          4068 => x"74",
          4069 => x"f6",
          4070 => x"93",
          4071 => x"ff",
          4072 => x"cc",
          4073 => x"80",
          4074 => x"2e",
          4075 => x"81",
          4076 => x"82",
          4077 => x"74",
          4078 => x"98",
          4079 => x"a4",
          4080 => x"2b",
          4081 => x"70",
          4082 => x"82",
          4083 => x"e0",
          4084 => x"51",
          4085 => x"58",
          4086 => x"77",
          4087 => x"06",
          4088 => x"81",
          4089 => x"08",
          4090 => x"0b",
          4091 => x"34",
          4092 => x"93",
          4093 => x"39",
          4094 => x"a8",
          4095 => x"93",
          4096 => x"af",
          4097 => x"7d",
          4098 => x"73",
          4099 => x"e1",
          4100 => x"29",
          4101 => x"05",
          4102 => x"04",
          4103 => x"33",
          4104 => x"2e",
          4105 => x"82",
          4106 => x"55",
          4107 => x"ab",
          4108 => x"2b",
          4109 => x"51",
          4110 => x"24",
          4111 => x"1a",
          4112 => x"81",
          4113 => x"81",
          4114 => x"81",
          4115 => x"70",
          4116 => x"93",
          4117 => x"51",
          4118 => x"82",
          4119 => x"81",
          4120 => x"74",
          4121 => x"34",
          4122 => x"ae",
          4123 => x"34",
          4124 => x"33",
          4125 => x"27",
          4126 => x"14",
          4127 => x"93",
          4128 => x"93",
          4129 => x"81",
          4130 => x"81",
          4131 => x"70",
          4132 => x"93",
          4133 => x"51",
          4134 => x"77",
          4135 => x"74",
          4136 => x"52",
          4137 => x"3f",
          4138 => x"0a",
          4139 => x"0a",
          4140 => x"2c",
          4141 => x"33",
          4142 => x"73",
          4143 => x"38",
          4144 => x"33",
          4145 => x"70",
          4146 => x"93",
          4147 => x"51",
          4148 => x"77",
          4149 => x"38",
          4150 => x"92",
          4151 => x"80",
          4152 => x"80",
          4153 => x"98",
          4154 => x"ac",
          4155 => x"55",
          4156 => x"e4",
          4157 => x"39",
          4158 => x"33",
          4159 => x"06",
          4160 => x"80",
          4161 => x"38",
          4162 => x"33",
          4163 => x"73",
          4164 => x"34",
          4165 => x"73",
          4166 => x"34",
          4167 => x"ce",
          4168 => x"b0",
          4169 => x"2b",
          4170 => x"82",
          4171 => x"57",
          4172 => x"74",
          4173 => x"38",
          4174 => x"81",
          4175 => x"34",
          4176 => x"e7",
          4177 => x"81",
          4178 => x"81",
          4179 => x"70",
          4180 => x"93",
          4181 => x"51",
          4182 => x"24",
          4183 => x"51",
          4184 => x"82",
          4185 => x"70",
          4186 => x"98",
          4187 => x"ac",
          4188 => x"56",
          4189 => x"24",
          4190 => x"88",
          4191 => x"3f",
          4192 => x"0a",
          4193 => x"0a",
          4194 => x"2c",
          4195 => x"33",
          4196 => x"75",
          4197 => x"38",
          4198 => x"82",
          4199 => x"7a",
          4200 => x"74",
          4201 => x"e6",
          4202 => x"93",
          4203 => x"51",
          4204 => x"82",
          4205 => x"81",
          4206 => x"73",
          4207 => x"93",
          4208 => x"73",
          4209 => x"c9",
          4210 => x"73",
          4211 => x"f3",
          4212 => x"bd",
          4213 => x"34",
          4214 => x"82",
          4215 => x"54",
          4216 => x"fa",
          4217 => x"51",
          4218 => x"82",
          4219 => x"ff",
          4220 => x"82",
          4221 => x"73",
          4222 => x"54",
          4223 => x"93",
          4224 => x"93",
          4225 => x"55",
          4226 => x"f9",
          4227 => x"14",
          4228 => x"93",
          4229 => x"98",
          4230 => x"2c",
          4231 => x"06",
          4232 => x"74",
          4233 => x"38",
          4234 => x"81",
          4235 => x"34",
          4236 => x"e5",
          4237 => x"81",
          4238 => x"81",
          4239 => x"70",
          4240 => x"93",
          4241 => x"51",
          4242 => x"24",
          4243 => x"51",
          4244 => x"82",
          4245 => x"70",
          4246 => x"98",
          4247 => x"ac",
          4248 => x"56",
          4249 => x"24",
          4250 => x"88",
          4251 => x"3f",
          4252 => x"0a",
          4253 => x"0a",
          4254 => x"2c",
          4255 => x"33",
          4256 => x"75",
          4257 => x"38",
          4258 => x"82",
          4259 => x"70",
          4260 => x"82",
          4261 => x"59",
          4262 => x"77",
          4263 => x"38",
          4264 => x"73",
          4265 => x"34",
          4266 => x"33",
          4267 => x"be",
          4268 => x"b0",
          4269 => x"ff",
          4270 => x"ac",
          4271 => x"54",
          4272 => x"dc",
          4273 => x"39",
          4274 => x"82",
          4275 => x"55",
          4276 => x"a4",
          4277 => x"cb",
          4278 => x"93",
          4279 => x"93",
          4280 => x"93",
          4281 => x"ff",
          4282 => x"53",
          4283 => x"51",
          4284 => x"93",
          4285 => x"39",
          4286 => x"82",
          4287 => x"fc",
          4288 => x"54",
          4289 => x"a5",
          4290 => x"ca",
          4291 => x"93",
          4292 => x"93",
          4293 => x"93",
          4294 => x"ff",
          4295 => x"53",
          4296 => x"51",
          4297 => x"ff",
          4298 => x"de",
          4299 => x"55",
          4300 => x"f7",
          4301 => x"51",
          4302 => x"80",
          4303 => x"93",
          4304 => x"06",
          4305 => x"8e",
          4306 => x"74",
          4307 => x"38",
          4308 => x"9d",
          4309 => x"39",
          4310 => x"82",
          4311 => x"84",
          4312 => x"54",
          4313 => x"a9",
          4314 => x"ca",
          4315 => x"93",
          4316 => x"93",
          4317 => x"93",
          4318 => x"ff",
          4319 => x"53",
          4320 => x"51",
          4321 => x"81",
          4322 => x"81",
          4323 => x"a8",
          4324 => x"55",
          4325 => x"f6",
          4326 => x"51",
          4327 => x"82",
          4328 => x"82",
          4329 => x"82",
          4330 => x"81",
          4331 => x"05",
          4332 => x"79",
          4333 => x"3f",
          4334 => x"53",
          4335 => x"33",
          4336 => x"ef",
          4337 => x"a9",
          4338 => x"b0",
          4339 => x"ff",
          4340 => x"ac",
          4341 => x"54",
          4342 => x"f6",
          4343 => x"14",
          4344 => x"93",
          4345 => x"1a",
          4346 => x"54",
          4347 => x"f6",
          4348 => x"93",
          4349 => x"73",
          4350 => x"f5",
          4351 => x"e1",
          4352 => x"93",
          4353 => x"05",
          4354 => x"93",
          4355 => x"e1",
          4356 => x"82",
          4357 => x"80",
          4358 => x"ac",
          4359 => x"93",
          4360 => x"3d",
          4361 => x"3d",
          4362 => x"05",
          4363 => x"52",
          4364 => x"87",
          4365 => x"ec",
          4366 => x"71",
          4367 => x"0c",
          4368 => x"04",
          4369 => x"02",
          4370 => x"02",
          4371 => x"05",
          4372 => x"83",
          4373 => x"26",
          4374 => x"72",
          4375 => x"c0",
          4376 => x"53",
          4377 => x"74",
          4378 => x"38",
          4379 => x"73",
          4380 => x"c0",
          4381 => x"51",
          4382 => x"85",
          4383 => x"98",
          4384 => x"52",
          4385 => x"82",
          4386 => x"70",
          4387 => x"38",
          4388 => x"8c",
          4389 => x"ec",
          4390 => x"fc",
          4391 => x"52",
          4392 => x"87",
          4393 => x"08",
          4394 => x"2e",
          4395 => x"82",
          4396 => x"34",
          4397 => x"13",
          4398 => x"82",
          4399 => x"86",
          4400 => x"f3",
          4401 => x"62",
          4402 => x"05",
          4403 => x"57",
          4404 => x"83",
          4405 => x"fe",
          4406 => x"93",
          4407 => x"06",
          4408 => x"71",
          4409 => x"71",
          4410 => x"2b",
          4411 => x"80",
          4412 => x"92",
          4413 => x"c0",
          4414 => x"41",
          4415 => x"5a",
          4416 => x"87",
          4417 => x"0c",
          4418 => x"84",
          4419 => x"08",
          4420 => x"70",
          4421 => x"53",
          4422 => x"2e",
          4423 => x"08",
          4424 => x"70",
          4425 => x"34",
          4426 => x"80",
          4427 => x"53",
          4428 => x"2e",
          4429 => x"53",
          4430 => x"26",
          4431 => x"80",
          4432 => x"87",
          4433 => x"08",
          4434 => x"38",
          4435 => x"8c",
          4436 => x"80",
          4437 => x"78",
          4438 => x"99",
          4439 => x"0c",
          4440 => x"8c",
          4441 => x"08",
          4442 => x"51",
          4443 => x"38",
          4444 => x"8d",
          4445 => x"17",
          4446 => x"81",
          4447 => x"53",
          4448 => x"2e",
          4449 => x"fc",
          4450 => x"52",
          4451 => x"7d",
          4452 => x"ed",
          4453 => x"80",
          4454 => x"71",
          4455 => x"38",
          4456 => x"53",
          4457 => x"84",
          4458 => x"0d",
          4459 => x"0d",
          4460 => x"02",
          4461 => x"05",
          4462 => x"58",
          4463 => x"80",
          4464 => x"fc",
          4465 => x"93",
          4466 => x"06",
          4467 => x"71",
          4468 => x"81",
          4469 => x"38",
          4470 => x"2b",
          4471 => x"80",
          4472 => x"92",
          4473 => x"c0",
          4474 => x"40",
          4475 => x"5a",
          4476 => x"c0",
          4477 => x"76",
          4478 => x"76",
          4479 => x"75",
          4480 => x"2a",
          4481 => x"51",
          4482 => x"80",
          4483 => x"7a",
          4484 => x"5c",
          4485 => x"81",
          4486 => x"81",
          4487 => x"06",
          4488 => x"80",
          4489 => x"87",
          4490 => x"08",
          4491 => x"38",
          4492 => x"8c",
          4493 => x"80",
          4494 => x"77",
          4495 => x"99",
          4496 => x"0c",
          4497 => x"8c",
          4498 => x"08",
          4499 => x"51",
          4500 => x"38",
          4501 => x"8d",
          4502 => x"70",
          4503 => x"84",
          4504 => x"5b",
          4505 => x"2e",
          4506 => x"fc",
          4507 => x"52",
          4508 => x"7d",
          4509 => x"f8",
          4510 => x"80",
          4511 => x"71",
          4512 => x"38",
          4513 => x"53",
          4514 => x"84",
          4515 => x"0d",
          4516 => x"0d",
          4517 => x"05",
          4518 => x"02",
          4519 => x"05",
          4520 => x"54",
          4521 => x"fe",
          4522 => x"84",
          4523 => x"53",
          4524 => x"80",
          4525 => x"0b",
          4526 => x"8c",
          4527 => x"71",
          4528 => x"dc",
          4529 => x"24",
          4530 => x"84",
          4531 => x"92",
          4532 => x"54",
          4533 => x"8d",
          4534 => x"39",
          4535 => x"80",
          4536 => x"cb",
          4537 => x"70",
          4538 => x"81",
          4539 => x"52",
          4540 => x"8a",
          4541 => x"98",
          4542 => x"71",
          4543 => x"c0",
          4544 => x"52",
          4545 => x"81",
          4546 => x"c0",
          4547 => x"53",
          4548 => x"82",
          4549 => x"71",
          4550 => x"39",
          4551 => x"39",
          4552 => x"77",
          4553 => x"81",
          4554 => x"72",
          4555 => x"84",
          4556 => x"73",
          4557 => x"0c",
          4558 => x"04",
          4559 => x"74",
          4560 => x"71",
          4561 => x"2b",
          4562 => x"84",
          4563 => x"84",
          4564 => x"fd",
          4565 => x"83",
          4566 => x"12",
          4567 => x"2b",
          4568 => x"07",
          4569 => x"70",
          4570 => x"2b",
          4571 => x"07",
          4572 => x"0c",
          4573 => x"56",
          4574 => x"3d",
          4575 => x"3d",
          4576 => x"84",
          4577 => x"22",
          4578 => x"72",
          4579 => x"54",
          4580 => x"2a",
          4581 => x"34",
          4582 => x"04",
          4583 => x"73",
          4584 => x"70",
          4585 => x"05",
          4586 => x"88",
          4587 => x"72",
          4588 => x"54",
          4589 => x"2a",
          4590 => x"70",
          4591 => x"34",
          4592 => x"51",
          4593 => x"83",
          4594 => x"fe",
          4595 => x"75",
          4596 => x"51",
          4597 => x"92",
          4598 => x"81",
          4599 => x"73",
          4600 => x"55",
          4601 => x"51",
          4602 => x"3d",
          4603 => x"3d",
          4604 => x"76",
          4605 => x"72",
          4606 => x"05",
          4607 => x"11",
          4608 => x"38",
          4609 => x"04",
          4610 => x"78",
          4611 => x"56",
          4612 => x"81",
          4613 => x"74",
          4614 => x"56",
          4615 => x"31",
          4616 => x"52",
          4617 => x"80",
          4618 => x"71",
          4619 => x"38",
          4620 => x"84",
          4621 => x"0d",
          4622 => x"0d",
          4623 => x"51",
          4624 => x"73",
          4625 => x"81",
          4626 => x"33",
          4627 => x"38",
          4628 => x"93",
          4629 => x"3d",
          4630 => x"0b",
          4631 => x"0c",
          4632 => x"82",
          4633 => x"04",
          4634 => x"7b",
          4635 => x"83",
          4636 => x"5a",
          4637 => x"80",
          4638 => x"54",
          4639 => x"53",
          4640 => x"53",
          4641 => x"52",
          4642 => x"3f",
          4643 => x"08",
          4644 => x"81",
          4645 => x"82",
          4646 => x"83",
          4647 => x"16",
          4648 => x"18",
          4649 => x"18",
          4650 => x"58",
          4651 => x"9f",
          4652 => x"33",
          4653 => x"2e",
          4654 => x"93",
          4655 => x"76",
          4656 => x"52",
          4657 => x"51",
          4658 => x"83",
          4659 => x"79",
          4660 => x"0c",
          4661 => x"04",
          4662 => x"78",
          4663 => x"80",
          4664 => x"17",
          4665 => x"38",
          4666 => x"fc",
          4667 => x"84",
          4668 => x"93",
          4669 => x"38",
          4670 => x"53",
          4671 => x"81",
          4672 => x"f7",
          4673 => x"93",
          4674 => x"2e",
          4675 => x"55",
          4676 => x"b0",
          4677 => x"82",
          4678 => x"88",
          4679 => x"f8",
          4680 => x"70",
          4681 => x"c0",
          4682 => x"84",
          4683 => x"93",
          4684 => x"91",
          4685 => x"55",
          4686 => x"09",
          4687 => x"f0",
          4688 => x"33",
          4689 => x"2e",
          4690 => x"80",
          4691 => x"80",
          4692 => x"84",
          4693 => x"17",
          4694 => x"fd",
          4695 => x"d4",
          4696 => x"b2",
          4697 => x"96",
          4698 => x"85",
          4699 => x"75",
          4700 => x"3f",
          4701 => x"e4",
          4702 => x"98",
          4703 => x"9c",
          4704 => x"08",
          4705 => x"17",
          4706 => x"3f",
          4707 => x"52",
          4708 => x"51",
          4709 => x"a0",
          4710 => x"05",
          4711 => x"0c",
          4712 => x"75",
          4713 => x"33",
          4714 => x"3f",
          4715 => x"34",
          4716 => x"52",
          4717 => x"51",
          4718 => x"82",
          4719 => x"80",
          4720 => x"81",
          4721 => x"93",
          4722 => x"3d",
          4723 => x"3d",
          4724 => x"1a",
          4725 => x"fe",
          4726 => x"54",
          4727 => x"73",
          4728 => x"8a",
          4729 => x"71",
          4730 => x"08",
          4731 => x"75",
          4732 => x"0c",
          4733 => x"04",
          4734 => x"7a",
          4735 => x"56",
          4736 => x"77",
          4737 => x"38",
          4738 => x"08",
          4739 => x"38",
          4740 => x"54",
          4741 => x"2e",
          4742 => x"72",
          4743 => x"38",
          4744 => x"8d",
          4745 => x"39",
          4746 => x"81",
          4747 => x"b6",
          4748 => x"2a",
          4749 => x"2a",
          4750 => x"05",
          4751 => x"55",
          4752 => x"82",
          4753 => x"81",
          4754 => x"83",
          4755 => x"b4",
          4756 => x"17",
          4757 => x"a4",
          4758 => x"55",
          4759 => x"57",
          4760 => x"3f",
          4761 => x"08",
          4762 => x"74",
          4763 => x"14",
          4764 => x"70",
          4765 => x"07",
          4766 => x"71",
          4767 => x"52",
          4768 => x"72",
          4769 => x"75",
          4770 => x"58",
          4771 => x"76",
          4772 => x"15",
          4773 => x"73",
          4774 => x"3f",
          4775 => x"08",
          4776 => x"76",
          4777 => x"06",
          4778 => x"05",
          4779 => x"3f",
          4780 => x"08",
          4781 => x"06",
          4782 => x"76",
          4783 => x"15",
          4784 => x"73",
          4785 => x"3f",
          4786 => x"08",
          4787 => x"82",
          4788 => x"06",
          4789 => x"05",
          4790 => x"3f",
          4791 => x"08",
          4792 => x"58",
          4793 => x"58",
          4794 => x"84",
          4795 => x"0d",
          4796 => x"0d",
          4797 => x"5a",
          4798 => x"59",
          4799 => x"82",
          4800 => x"98",
          4801 => x"82",
          4802 => x"33",
          4803 => x"2e",
          4804 => x"72",
          4805 => x"38",
          4806 => x"8d",
          4807 => x"39",
          4808 => x"81",
          4809 => x"f7",
          4810 => x"2a",
          4811 => x"2a",
          4812 => x"05",
          4813 => x"55",
          4814 => x"82",
          4815 => x"59",
          4816 => x"08",
          4817 => x"74",
          4818 => x"16",
          4819 => x"16",
          4820 => x"59",
          4821 => x"53",
          4822 => x"8f",
          4823 => x"2b",
          4824 => x"74",
          4825 => x"71",
          4826 => x"72",
          4827 => x"0b",
          4828 => x"74",
          4829 => x"17",
          4830 => x"75",
          4831 => x"3f",
          4832 => x"08",
          4833 => x"84",
          4834 => x"38",
          4835 => x"06",
          4836 => x"78",
          4837 => x"54",
          4838 => x"77",
          4839 => x"33",
          4840 => x"71",
          4841 => x"51",
          4842 => x"34",
          4843 => x"76",
          4844 => x"17",
          4845 => x"75",
          4846 => x"3f",
          4847 => x"08",
          4848 => x"84",
          4849 => x"38",
          4850 => x"ff",
          4851 => x"10",
          4852 => x"76",
          4853 => x"51",
          4854 => x"be",
          4855 => x"2a",
          4856 => x"05",
          4857 => x"f9",
          4858 => x"93",
          4859 => x"82",
          4860 => x"ab",
          4861 => x"0a",
          4862 => x"2b",
          4863 => x"70",
          4864 => x"70",
          4865 => x"54",
          4866 => x"82",
          4867 => x"8f",
          4868 => x"07",
          4869 => x"f7",
          4870 => x"0b",
          4871 => x"78",
          4872 => x"0c",
          4873 => x"04",
          4874 => x"7a",
          4875 => x"08",
          4876 => x"59",
          4877 => x"a4",
          4878 => x"17",
          4879 => x"38",
          4880 => x"aa",
          4881 => x"73",
          4882 => x"fd",
          4883 => x"93",
          4884 => x"82",
          4885 => x"80",
          4886 => x"39",
          4887 => x"eb",
          4888 => x"80",
          4889 => x"93",
          4890 => x"80",
          4891 => x"52",
          4892 => x"84",
          4893 => x"84",
          4894 => x"93",
          4895 => x"2e",
          4896 => x"82",
          4897 => x"81",
          4898 => x"82",
          4899 => x"ff",
          4900 => x"80",
          4901 => x"75",
          4902 => x"3f",
          4903 => x"08",
          4904 => x"16",
          4905 => x"90",
          4906 => x"55",
          4907 => x"27",
          4908 => x"15",
          4909 => x"84",
          4910 => x"07",
          4911 => x"17",
          4912 => x"76",
          4913 => x"a6",
          4914 => x"73",
          4915 => x"0c",
          4916 => x"04",
          4917 => x"7c",
          4918 => x"59",
          4919 => x"95",
          4920 => x"08",
          4921 => x"2e",
          4922 => x"17",
          4923 => x"b2",
          4924 => x"ae",
          4925 => x"7a",
          4926 => x"3f",
          4927 => x"82",
          4928 => x"27",
          4929 => x"82",
          4930 => x"55",
          4931 => x"08",
          4932 => x"d2",
          4933 => x"08",
          4934 => x"08",
          4935 => x"38",
          4936 => x"17",
          4937 => x"54",
          4938 => x"82",
          4939 => x"7a",
          4940 => x"06",
          4941 => x"81",
          4942 => x"17",
          4943 => x"83",
          4944 => x"75",
          4945 => x"f9",
          4946 => x"59",
          4947 => x"08",
          4948 => x"81",
          4949 => x"82",
          4950 => x"59",
          4951 => x"08",
          4952 => x"70",
          4953 => x"25",
          4954 => x"82",
          4955 => x"54",
          4956 => x"55",
          4957 => x"38",
          4958 => x"08",
          4959 => x"38",
          4960 => x"54",
          4961 => x"90",
          4962 => x"18",
          4963 => x"38",
          4964 => x"39",
          4965 => x"38",
          4966 => x"16",
          4967 => x"08",
          4968 => x"38",
          4969 => x"78",
          4970 => x"38",
          4971 => x"51",
          4972 => x"82",
          4973 => x"80",
          4974 => x"80",
          4975 => x"84",
          4976 => x"09",
          4977 => x"38",
          4978 => x"08",
          4979 => x"84",
          4980 => x"30",
          4981 => x"80",
          4982 => x"07",
          4983 => x"55",
          4984 => x"38",
          4985 => x"09",
          4986 => x"ae",
          4987 => x"80",
          4988 => x"53",
          4989 => x"51",
          4990 => x"82",
          4991 => x"82",
          4992 => x"30",
          4993 => x"84",
          4994 => x"25",
          4995 => x"79",
          4996 => x"38",
          4997 => x"8f",
          4998 => x"79",
          4999 => x"f9",
          5000 => x"93",
          5001 => x"74",
          5002 => x"8c",
          5003 => x"17",
          5004 => x"90",
          5005 => x"54",
          5006 => x"86",
          5007 => x"90",
          5008 => x"17",
          5009 => x"54",
          5010 => x"34",
          5011 => x"56",
          5012 => x"90",
          5013 => x"80",
          5014 => x"82",
          5015 => x"55",
          5016 => x"56",
          5017 => x"82",
          5018 => x"8c",
          5019 => x"f8",
          5020 => x"70",
          5021 => x"f0",
          5022 => x"84",
          5023 => x"56",
          5024 => x"08",
          5025 => x"7b",
          5026 => x"f6",
          5027 => x"93",
          5028 => x"93",
          5029 => x"17",
          5030 => x"80",
          5031 => x"b4",
          5032 => x"57",
          5033 => x"77",
          5034 => x"81",
          5035 => x"15",
          5036 => x"78",
          5037 => x"81",
          5038 => x"53",
          5039 => x"15",
          5040 => x"e9",
          5041 => x"84",
          5042 => x"df",
          5043 => x"22",
          5044 => x"30",
          5045 => x"70",
          5046 => x"51",
          5047 => x"82",
          5048 => x"8a",
          5049 => x"f8",
          5050 => x"7c",
          5051 => x"56",
          5052 => x"80",
          5053 => x"f1",
          5054 => x"06",
          5055 => x"e9",
          5056 => x"18",
          5057 => x"08",
          5058 => x"38",
          5059 => x"82",
          5060 => x"38",
          5061 => x"54",
          5062 => x"74",
          5063 => x"82",
          5064 => x"22",
          5065 => x"79",
          5066 => x"38",
          5067 => x"98",
          5068 => x"cd",
          5069 => x"22",
          5070 => x"54",
          5071 => x"26",
          5072 => x"52",
          5073 => x"b0",
          5074 => x"84",
          5075 => x"93",
          5076 => x"2e",
          5077 => x"0b",
          5078 => x"08",
          5079 => x"98",
          5080 => x"93",
          5081 => x"85",
          5082 => x"bd",
          5083 => x"31",
          5084 => x"73",
          5085 => x"f4",
          5086 => x"93",
          5087 => x"18",
          5088 => x"18",
          5089 => x"08",
          5090 => x"72",
          5091 => x"38",
          5092 => x"58",
          5093 => x"89",
          5094 => x"18",
          5095 => x"ff",
          5096 => x"05",
          5097 => x"80",
          5098 => x"93",
          5099 => x"3d",
          5100 => x"3d",
          5101 => x"08",
          5102 => x"a0",
          5103 => x"54",
          5104 => x"77",
          5105 => x"80",
          5106 => x"0c",
          5107 => x"53",
          5108 => x"80",
          5109 => x"38",
          5110 => x"06",
          5111 => x"b5",
          5112 => x"98",
          5113 => x"14",
          5114 => x"92",
          5115 => x"2a",
          5116 => x"56",
          5117 => x"26",
          5118 => x"80",
          5119 => x"16",
          5120 => x"77",
          5121 => x"53",
          5122 => x"38",
          5123 => x"51",
          5124 => x"82",
          5125 => x"53",
          5126 => x"0b",
          5127 => x"08",
          5128 => x"38",
          5129 => x"93",
          5130 => x"2e",
          5131 => x"98",
          5132 => x"93",
          5133 => x"80",
          5134 => x"8a",
          5135 => x"15",
          5136 => x"80",
          5137 => x"14",
          5138 => x"51",
          5139 => x"82",
          5140 => x"53",
          5141 => x"93",
          5142 => x"2e",
          5143 => x"82",
          5144 => x"84",
          5145 => x"ba",
          5146 => x"82",
          5147 => x"ff",
          5148 => x"82",
          5149 => x"52",
          5150 => x"f3",
          5151 => x"84",
          5152 => x"72",
          5153 => x"72",
          5154 => x"f2",
          5155 => x"93",
          5156 => x"15",
          5157 => x"15",
          5158 => x"b4",
          5159 => x"0c",
          5160 => x"82",
          5161 => x"8a",
          5162 => x"f7",
          5163 => x"7d",
          5164 => x"5b",
          5165 => x"76",
          5166 => x"3f",
          5167 => x"08",
          5168 => x"84",
          5169 => x"38",
          5170 => x"08",
          5171 => x"08",
          5172 => x"f0",
          5173 => x"93",
          5174 => x"82",
          5175 => x"80",
          5176 => x"93",
          5177 => x"18",
          5178 => x"51",
          5179 => x"81",
          5180 => x"81",
          5181 => x"81",
          5182 => x"84",
          5183 => x"83",
          5184 => x"77",
          5185 => x"72",
          5186 => x"38",
          5187 => x"75",
          5188 => x"81",
          5189 => x"a5",
          5190 => x"84",
          5191 => x"52",
          5192 => x"8e",
          5193 => x"84",
          5194 => x"93",
          5195 => x"2e",
          5196 => x"73",
          5197 => x"81",
          5198 => x"87",
          5199 => x"93",
          5200 => x"3d",
          5201 => x"3d",
          5202 => x"11",
          5203 => x"ec",
          5204 => x"84",
          5205 => x"ff",
          5206 => x"33",
          5207 => x"71",
          5208 => x"81",
          5209 => x"94",
          5210 => x"d0",
          5211 => x"84",
          5212 => x"73",
          5213 => x"82",
          5214 => x"85",
          5215 => x"fc",
          5216 => x"79",
          5217 => x"ff",
          5218 => x"12",
          5219 => x"eb",
          5220 => x"70",
          5221 => x"72",
          5222 => x"81",
          5223 => x"73",
          5224 => x"94",
          5225 => x"d6",
          5226 => x"0d",
          5227 => x"0d",
          5228 => x"55",
          5229 => x"5a",
          5230 => x"08",
          5231 => x"8a",
          5232 => x"08",
          5233 => x"ee",
          5234 => x"93",
          5235 => x"82",
          5236 => x"80",
          5237 => x"15",
          5238 => x"55",
          5239 => x"38",
          5240 => x"e6",
          5241 => x"33",
          5242 => x"70",
          5243 => x"58",
          5244 => x"86",
          5245 => x"93",
          5246 => x"73",
          5247 => x"83",
          5248 => x"73",
          5249 => x"38",
          5250 => x"06",
          5251 => x"80",
          5252 => x"75",
          5253 => x"38",
          5254 => x"08",
          5255 => x"54",
          5256 => x"2e",
          5257 => x"83",
          5258 => x"73",
          5259 => x"38",
          5260 => x"51",
          5261 => x"82",
          5262 => x"58",
          5263 => x"08",
          5264 => x"15",
          5265 => x"38",
          5266 => x"0b",
          5267 => x"77",
          5268 => x"0c",
          5269 => x"04",
          5270 => x"77",
          5271 => x"54",
          5272 => x"51",
          5273 => x"82",
          5274 => x"55",
          5275 => x"08",
          5276 => x"14",
          5277 => x"51",
          5278 => x"82",
          5279 => x"55",
          5280 => x"08",
          5281 => x"53",
          5282 => x"08",
          5283 => x"08",
          5284 => x"3f",
          5285 => x"14",
          5286 => x"08",
          5287 => x"3f",
          5288 => x"17",
          5289 => x"93",
          5290 => x"3d",
          5291 => x"3d",
          5292 => x"08",
          5293 => x"54",
          5294 => x"53",
          5295 => x"82",
          5296 => x"8d",
          5297 => x"08",
          5298 => x"34",
          5299 => x"15",
          5300 => x"0d",
          5301 => x"0d",
          5302 => x"57",
          5303 => x"17",
          5304 => x"08",
          5305 => x"82",
          5306 => x"89",
          5307 => x"55",
          5308 => x"14",
          5309 => x"16",
          5310 => x"71",
          5311 => x"38",
          5312 => x"09",
          5313 => x"38",
          5314 => x"73",
          5315 => x"81",
          5316 => x"ae",
          5317 => x"05",
          5318 => x"15",
          5319 => x"70",
          5320 => x"34",
          5321 => x"8a",
          5322 => x"38",
          5323 => x"05",
          5324 => x"81",
          5325 => x"17",
          5326 => x"12",
          5327 => x"34",
          5328 => x"9c",
          5329 => x"e8",
          5330 => x"93",
          5331 => x"0c",
          5332 => x"e7",
          5333 => x"93",
          5334 => x"17",
          5335 => x"51",
          5336 => x"82",
          5337 => x"84",
          5338 => x"3d",
          5339 => x"3d",
          5340 => x"08",
          5341 => x"61",
          5342 => x"55",
          5343 => x"2e",
          5344 => x"55",
          5345 => x"2e",
          5346 => x"80",
          5347 => x"94",
          5348 => x"1c",
          5349 => x"81",
          5350 => x"61",
          5351 => x"56",
          5352 => x"2e",
          5353 => x"83",
          5354 => x"73",
          5355 => x"70",
          5356 => x"25",
          5357 => x"51",
          5358 => x"38",
          5359 => x"0c",
          5360 => x"51",
          5361 => x"26",
          5362 => x"80",
          5363 => x"34",
          5364 => x"51",
          5365 => x"82",
          5366 => x"55",
          5367 => x"91",
          5368 => x"1d",
          5369 => x"8b",
          5370 => x"79",
          5371 => x"3f",
          5372 => x"57",
          5373 => x"55",
          5374 => x"2e",
          5375 => x"80",
          5376 => x"18",
          5377 => x"1a",
          5378 => x"70",
          5379 => x"2a",
          5380 => x"07",
          5381 => x"5a",
          5382 => x"8c",
          5383 => x"54",
          5384 => x"81",
          5385 => x"39",
          5386 => x"70",
          5387 => x"2a",
          5388 => x"75",
          5389 => x"8c",
          5390 => x"2e",
          5391 => x"a0",
          5392 => x"38",
          5393 => x"0c",
          5394 => x"76",
          5395 => x"38",
          5396 => x"b8",
          5397 => x"70",
          5398 => x"5a",
          5399 => x"76",
          5400 => x"38",
          5401 => x"70",
          5402 => x"dc",
          5403 => x"72",
          5404 => x"80",
          5405 => x"51",
          5406 => x"73",
          5407 => x"38",
          5408 => x"18",
          5409 => x"1a",
          5410 => x"55",
          5411 => x"2e",
          5412 => x"83",
          5413 => x"73",
          5414 => x"70",
          5415 => x"25",
          5416 => x"51",
          5417 => x"38",
          5418 => x"75",
          5419 => x"81",
          5420 => x"81",
          5421 => x"27",
          5422 => x"73",
          5423 => x"38",
          5424 => x"70",
          5425 => x"32",
          5426 => x"80",
          5427 => x"2a",
          5428 => x"56",
          5429 => x"81",
          5430 => x"57",
          5431 => x"f5",
          5432 => x"2b",
          5433 => x"25",
          5434 => x"80",
          5435 => x"ff",
          5436 => x"57",
          5437 => x"e6",
          5438 => x"93",
          5439 => x"2e",
          5440 => x"18",
          5441 => x"1a",
          5442 => x"56",
          5443 => x"3f",
          5444 => x"08",
          5445 => x"e8",
          5446 => x"54",
          5447 => x"80",
          5448 => x"17",
          5449 => x"34",
          5450 => x"11",
          5451 => x"74",
          5452 => x"75",
          5453 => x"90",
          5454 => x"3f",
          5455 => x"08",
          5456 => x"9f",
          5457 => x"99",
          5458 => x"e0",
          5459 => x"ff",
          5460 => x"79",
          5461 => x"74",
          5462 => x"57",
          5463 => x"77",
          5464 => x"76",
          5465 => x"38",
          5466 => x"73",
          5467 => x"09",
          5468 => x"38",
          5469 => x"84",
          5470 => x"27",
          5471 => x"39",
          5472 => x"f2",
          5473 => x"80",
          5474 => x"54",
          5475 => x"34",
          5476 => x"58",
          5477 => x"f2",
          5478 => x"93",
          5479 => x"82",
          5480 => x"80",
          5481 => x"1b",
          5482 => x"51",
          5483 => x"82",
          5484 => x"56",
          5485 => x"08",
          5486 => x"9c",
          5487 => x"33",
          5488 => x"80",
          5489 => x"38",
          5490 => x"bf",
          5491 => x"86",
          5492 => x"15",
          5493 => x"2a",
          5494 => x"51",
          5495 => x"92",
          5496 => x"79",
          5497 => x"e4",
          5498 => x"93",
          5499 => x"2e",
          5500 => x"52",
          5501 => x"ba",
          5502 => x"39",
          5503 => x"33",
          5504 => x"80",
          5505 => x"74",
          5506 => x"81",
          5507 => x"38",
          5508 => x"70",
          5509 => x"82",
          5510 => x"54",
          5511 => x"96",
          5512 => x"06",
          5513 => x"2e",
          5514 => x"ff",
          5515 => x"1c",
          5516 => x"80",
          5517 => x"81",
          5518 => x"ba",
          5519 => x"b6",
          5520 => x"2a",
          5521 => x"51",
          5522 => x"38",
          5523 => x"70",
          5524 => x"81",
          5525 => x"55",
          5526 => x"e1",
          5527 => x"08",
          5528 => x"1d",
          5529 => x"7c",
          5530 => x"3f",
          5531 => x"08",
          5532 => x"fa",
          5533 => x"82",
          5534 => x"8f",
          5535 => x"f6",
          5536 => x"5b",
          5537 => x"70",
          5538 => x"59",
          5539 => x"73",
          5540 => x"c6",
          5541 => x"81",
          5542 => x"70",
          5543 => x"52",
          5544 => x"8d",
          5545 => x"38",
          5546 => x"09",
          5547 => x"a5",
          5548 => x"d0",
          5549 => x"ff",
          5550 => x"53",
          5551 => x"91",
          5552 => x"73",
          5553 => x"d0",
          5554 => x"71",
          5555 => x"f7",
          5556 => x"81",
          5557 => x"55",
          5558 => x"55",
          5559 => x"81",
          5560 => x"74",
          5561 => x"56",
          5562 => x"12",
          5563 => x"70",
          5564 => x"38",
          5565 => x"81",
          5566 => x"51",
          5567 => x"51",
          5568 => x"89",
          5569 => x"70",
          5570 => x"53",
          5571 => x"70",
          5572 => x"51",
          5573 => x"09",
          5574 => x"38",
          5575 => x"38",
          5576 => x"77",
          5577 => x"70",
          5578 => x"2a",
          5579 => x"07",
          5580 => x"51",
          5581 => x"8f",
          5582 => x"84",
          5583 => x"83",
          5584 => x"94",
          5585 => x"74",
          5586 => x"38",
          5587 => x"0c",
          5588 => x"86",
          5589 => x"c8",
          5590 => x"82",
          5591 => x"8c",
          5592 => x"fa",
          5593 => x"56",
          5594 => x"17",
          5595 => x"b0",
          5596 => x"52",
          5597 => x"e0",
          5598 => x"82",
          5599 => x"81",
          5600 => x"b2",
          5601 => x"b4",
          5602 => x"84",
          5603 => x"ff",
          5604 => x"55",
          5605 => x"d5",
          5606 => x"06",
          5607 => x"80",
          5608 => x"33",
          5609 => x"81",
          5610 => x"81",
          5611 => x"81",
          5612 => x"eb",
          5613 => x"70",
          5614 => x"07",
          5615 => x"73",
          5616 => x"81",
          5617 => x"81",
          5618 => x"83",
          5619 => x"a0",
          5620 => x"16",
          5621 => x"3f",
          5622 => x"08",
          5623 => x"84",
          5624 => x"9d",
          5625 => x"81",
          5626 => x"81",
          5627 => x"e0",
          5628 => x"93",
          5629 => x"82",
          5630 => x"80",
          5631 => x"82",
          5632 => x"93",
          5633 => x"3d",
          5634 => x"3d",
          5635 => x"84",
          5636 => x"05",
          5637 => x"80",
          5638 => x"51",
          5639 => x"82",
          5640 => x"58",
          5641 => x"0b",
          5642 => x"08",
          5643 => x"38",
          5644 => x"08",
          5645 => x"93",
          5646 => x"08",
          5647 => x"56",
          5648 => x"86",
          5649 => x"75",
          5650 => x"fe",
          5651 => x"54",
          5652 => x"2e",
          5653 => x"14",
          5654 => x"ca",
          5655 => x"84",
          5656 => x"06",
          5657 => x"54",
          5658 => x"38",
          5659 => x"86",
          5660 => x"82",
          5661 => x"06",
          5662 => x"56",
          5663 => x"38",
          5664 => x"80",
          5665 => x"81",
          5666 => x"52",
          5667 => x"51",
          5668 => x"82",
          5669 => x"81",
          5670 => x"81",
          5671 => x"83",
          5672 => x"87",
          5673 => x"2e",
          5674 => x"82",
          5675 => x"06",
          5676 => x"56",
          5677 => x"38",
          5678 => x"74",
          5679 => x"a3",
          5680 => x"84",
          5681 => x"06",
          5682 => x"2e",
          5683 => x"80",
          5684 => x"3d",
          5685 => x"83",
          5686 => x"15",
          5687 => x"53",
          5688 => x"8d",
          5689 => x"15",
          5690 => x"3f",
          5691 => x"08",
          5692 => x"70",
          5693 => x"0c",
          5694 => x"16",
          5695 => x"80",
          5696 => x"80",
          5697 => x"54",
          5698 => x"84",
          5699 => x"5b",
          5700 => x"80",
          5701 => x"7a",
          5702 => x"fc",
          5703 => x"93",
          5704 => x"ff",
          5705 => x"77",
          5706 => x"81",
          5707 => x"76",
          5708 => x"81",
          5709 => x"2e",
          5710 => x"8d",
          5711 => x"26",
          5712 => x"bf",
          5713 => x"f4",
          5714 => x"84",
          5715 => x"ff",
          5716 => x"84",
          5717 => x"81",
          5718 => x"38",
          5719 => x"51",
          5720 => x"82",
          5721 => x"83",
          5722 => x"58",
          5723 => x"80",
          5724 => x"db",
          5725 => x"93",
          5726 => x"77",
          5727 => x"80",
          5728 => x"82",
          5729 => x"c4",
          5730 => x"11",
          5731 => x"06",
          5732 => x"8d",
          5733 => x"26",
          5734 => x"74",
          5735 => x"78",
          5736 => x"c1",
          5737 => x"59",
          5738 => x"15",
          5739 => x"2e",
          5740 => x"13",
          5741 => x"72",
          5742 => x"38",
          5743 => x"eb",
          5744 => x"14",
          5745 => x"3f",
          5746 => x"08",
          5747 => x"84",
          5748 => x"23",
          5749 => x"57",
          5750 => x"83",
          5751 => x"c7",
          5752 => x"d8",
          5753 => x"84",
          5754 => x"ff",
          5755 => x"8d",
          5756 => x"14",
          5757 => x"3f",
          5758 => x"08",
          5759 => x"14",
          5760 => x"3f",
          5761 => x"08",
          5762 => x"06",
          5763 => x"72",
          5764 => x"97",
          5765 => x"22",
          5766 => x"84",
          5767 => x"5a",
          5768 => x"83",
          5769 => x"14",
          5770 => x"79",
          5771 => x"96",
          5772 => x"93",
          5773 => x"82",
          5774 => x"80",
          5775 => x"38",
          5776 => x"08",
          5777 => x"ff",
          5778 => x"38",
          5779 => x"83",
          5780 => x"83",
          5781 => x"74",
          5782 => x"85",
          5783 => x"89",
          5784 => x"76",
          5785 => x"c3",
          5786 => x"70",
          5787 => x"7b",
          5788 => x"73",
          5789 => x"17",
          5790 => x"ac",
          5791 => x"55",
          5792 => x"09",
          5793 => x"38",
          5794 => x"51",
          5795 => x"82",
          5796 => x"83",
          5797 => x"53",
          5798 => x"82",
          5799 => x"82",
          5800 => x"e0",
          5801 => x"ab",
          5802 => x"84",
          5803 => x"0c",
          5804 => x"53",
          5805 => x"56",
          5806 => x"81",
          5807 => x"13",
          5808 => x"74",
          5809 => x"82",
          5810 => x"74",
          5811 => x"81",
          5812 => x"06",
          5813 => x"83",
          5814 => x"2a",
          5815 => x"72",
          5816 => x"26",
          5817 => x"ff",
          5818 => x"0c",
          5819 => x"15",
          5820 => x"0b",
          5821 => x"76",
          5822 => x"81",
          5823 => x"38",
          5824 => x"51",
          5825 => x"82",
          5826 => x"83",
          5827 => x"53",
          5828 => x"09",
          5829 => x"f9",
          5830 => x"52",
          5831 => x"b8",
          5832 => x"84",
          5833 => x"38",
          5834 => x"08",
          5835 => x"84",
          5836 => x"d8",
          5837 => x"93",
          5838 => x"ff",
          5839 => x"72",
          5840 => x"2e",
          5841 => x"80",
          5842 => x"14",
          5843 => x"3f",
          5844 => x"08",
          5845 => x"a4",
          5846 => x"81",
          5847 => x"84",
          5848 => x"d7",
          5849 => x"93",
          5850 => x"8a",
          5851 => x"2e",
          5852 => x"9d",
          5853 => x"14",
          5854 => x"3f",
          5855 => x"08",
          5856 => x"84",
          5857 => x"d7",
          5858 => x"93",
          5859 => x"15",
          5860 => x"34",
          5861 => x"22",
          5862 => x"72",
          5863 => x"23",
          5864 => x"23",
          5865 => x"15",
          5866 => x"75",
          5867 => x"0c",
          5868 => x"04",
          5869 => x"77",
          5870 => x"73",
          5871 => x"38",
          5872 => x"72",
          5873 => x"38",
          5874 => x"71",
          5875 => x"38",
          5876 => x"84",
          5877 => x"52",
          5878 => x"09",
          5879 => x"38",
          5880 => x"51",
          5881 => x"82",
          5882 => x"81",
          5883 => x"88",
          5884 => x"08",
          5885 => x"39",
          5886 => x"73",
          5887 => x"74",
          5888 => x"0c",
          5889 => x"04",
          5890 => x"02",
          5891 => x"7a",
          5892 => x"fc",
          5893 => x"f4",
          5894 => x"54",
          5895 => x"93",
          5896 => x"bc",
          5897 => x"84",
          5898 => x"82",
          5899 => x"70",
          5900 => x"73",
          5901 => x"38",
          5902 => x"78",
          5903 => x"2e",
          5904 => x"74",
          5905 => x"0c",
          5906 => x"80",
          5907 => x"80",
          5908 => x"70",
          5909 => x"51",
          5910 => x"82",
          5911 => x"54",
          5912 => x"84",
          5913 => x"0d",
          5914 => x"0d",
          5915 => x"05",
          5916 => x"33",
          5917 => x"54",
          5918 => x"84",
          5919 => x"bf",
          5920 => x"98",
          5921 => x"53",
          5922 => x"05",
          5923 => x"fa",
          5924 => x"84",
          5925 => x"93",
          5926 => x"a4",
          5927 => x"68",
          5928 => x"70",
          5929 => x"c6",
          5930 => x"84",
          5931 => x"93",
          5932 => x"38",
          5933 => x"05",
          5934 => x"2b",
          5935 => x"80",
          5936 => x"86",
          5937 => x"06",
          5938 => x"2e",
          5939 => x"74",
          5940 => x"38",
          5941 => x"09",
          5942 => x"38",
          5943 => x"f8",
          5944 => x"84",
          5945 => x"39",
          5946 => x"33",
          5947 => x"73",
          5948 => x"77",
          5949 => x"81",
          5950 => x"73",
          5951 => x"38",
          5952 => x"bc",
          5953 => x"07",
          5954 => x"b4",
          5955 => x"2a",
          5956 => x"51",
          5957 => x"2e",
          5958 => x"62",
          5959 => x"e8",
          5960 => x"93",
          5961 => x"82",
          5962 => x"52",
          5963 => x"51",
          5964 => x"62",
          5965 => x"8b",
          5966 => x"53",
          5967 => x"51",
          5968 => x"80",
          5969 => x"05",
          5970 => x"3f",
          5971 => x"0b",
          5972 => x"75",
          5973 => x"f1",
          5974 => x"11",
          5975 => x"80",
          5976 => x"97",
          5977 => x"51",
          5978 => x"82",
          5979 => x"55",
          5980 => x"08",
          5981 => x"b7",
          5982 => x"c4",
          5983 => x"05",
          5984 => x"2a",
          5985 => x"51",
          5986 => x"80",
          5987 => x"84",
          5988 => x"39",
          5989 => x"70",
          5990 => x"54",
          5991 => x"a9",
          5992 => x"06",
          5993 => x"2e",
          5994 => x"55",
          5995 => x"73",
          5996 => x"d6",
          5997 => x"93",
          5998 => x"ff",
          5999 => x"0c",
          6000 => x"93",
          6001 => x"f8",
          6002 => x"2a",
          6003 => x"51",
          6004 => x"2e",
          6005 => x"80",
          6006 => x"7a",
          6007 => x"a0",
          6008 => x"a4",
          6009 => x"53",
          6010 => x"e6",
          6011 => x"93",
          6012 => x"93",
          6013 => x"1b",
          6014 => x"05",
          6015 => x"d3",
          6016 => x"84",
          6017 => x"84",
          6018 => x"0c",
          6019 => x"56",
          6020 => x"84",
          6021 => x"90",
          6022 => x"0b",
          6023 => x"80",
          6024 => x"0c",
          6025 => x"1a",
          6026 => x"2a",
          6027 => x"51",
          6028 => x"2e",
          6029 => x"82",
          6030 => x"80",
          6031 => x"38",
          6032 => x"08",
          6033 => x"8a",
          6034 => x"89",
          6035 => x"59",
          6036 => x"76",
          6037 => x"d7",
          6038 => x"93",
          6039 => x"82",
          6040 => x"81",
          6041 => x"82",
          6042 => x"84",
          6043 => x"09",
          6044 => x"38",
          6045 => x"78",
          6046 => x"30",
          6047 => x"80",
          6048 => x"77",
          6049 => x"38",
          6050 => x"06",
          6051 => x"c3",
          6052 => x"1a",
          6053 => x"38",
          6054 => x"06",
          6055 => x"2e",
          6056 => x"52",
          6057 => x"a6",
          6058 => x"84",
          6059 => x"82",
          6060 => x"75",
          6061 => x"93",
          6062 => x"9c",
          6063 => x"39",
          6064 => x"74",
          6065 => x"93",
          6066 => x"3d",
          6067 => x"3d",
          6068 => x"65",
          6069 => x"5d",
          6070 => x"0c",
          6071 => x"05",
          6072 => x"f9",
          6073 => x"93",
          6074 => x"82",
          6075 => x"8a",
          6076 => x"33",
          6077 => x"2e",
          6078 => x"56",
          6079 => x"90",
          6080 => x"06",
          6081 => x"74",
          6082 => x"b6",
          6083 => x"82",
          6084 => x"34",
          6085 => x"aa",
          6086 => x"91",
          6087 => x"56",
          6088 => x"8c",
          6089 => x"1a",
          6090 => x"74",
          6091 => x"38",
          6092 => x"80",
          6093 => x"38",
          6094 => x"70",
          6095 => x"56",
          6096 => x"b2",
          6097 => x"11",
          6098 => x"77",
          6099 => x"5b",
          6100 => x"38",
          6101 => x"88",
          6102 => x"8f",
          6103 => x"08",
          6104 => x"d5",
          6105 => x"93",
          6106 => x"81",
          6107 => x"9f",
          6108 => x"2e",
          6109 => x"74",
          6110 => x"98",
          6111 => x"7e",
          6112 => x"3f",
          6113 => x"08",
          6114 => x"83",
          6115 => x"84",
          6116 => x"89",
          6117 => x"77",
          6118 => x"d6",
          6119 => x"7f",
          6120 => x"58",
          6121 => x"75",
          6122 => x"75",
          6123 => x"77",
          6124 => x"7c",
          6125 => x"33",
          6126 => x"3f",
          6127 => x"08",
          6128 => x"7e",
          6129 => x"56",
          6130 => x"2e",
          6131 => x"16",
          6132 => x"55",
          6133 => x"94",
          6134 => x"53",
          6135 => x"b0",
          6136 => x"31",
          6137 => x"05",
          6138 => x"3f",
          6139 => x"56",
          6140 => x"9c",
          6141 => x"19",
          6142 => x"06",
          6143 => x"31",
          6144 => x"76",
          6145 => x"7b",
          6146 => x"08",
          6147 => x"d1",
          6148 => x"93",
          6149 => x"81",
          6150 => x"94",
          6151 => x"ff",
          6152 => x"05",
          6153 => x"cf",
          6154 => x"76",
          6155 => x"17",
          6156 => x"1e",
          6157 => x"18",
          6158 => x"5e",
          6159 => x"39",
          6160 => x"82",
          6161 => x"90",
          6162 => x"f2",
          6163 => x"63",
          6164 => x"40",
          6165 => x"7e",
          6166 => x"fc",
          6167 => x"51",
          6168 => x"82",
          6169 => x"55",
          6170 => x"08",
          6171 => x"18",
          6172 => x"80",
          6173 => x"74",
          6174 => x"39",
          6175 => x"70",
          6176 => x"81",
          6177 => x"56",
          6178 => x"80",
          6179 => x"38",
          6180 => x"0b",
          6181 => x"82",
          6182 => x"39",
          6183 => x"19",
          6184 => x"83",
          6185 => x"18",
          6186 => x"56",
          6187 => x"27",
          6188 => x"09",
          6189 => x"2e",
          6190 => x"94",
          6191 => x"83",
          6192 => x"56",
          6193 => x"38",
          6194 => x"22",
          6195 => x"89",
          6196 => x"55",
          6197 => x"75",
          6198 => x"18",
          6199 => x"9c",
          6200 => x"85",
          6201 => x"08",
          6202 => x"d7",
          6203 => x"93",
          6204 => x"82",
          6205 => x"80",
          6206 => x"38",
          6207 => x"ff",
          6208 => x"ff",
          6209 => x"38",
          6210 => x"0c",
          6211 => x"85",
          6212 => x"19",
          6213 => x"b0",
          6214 => x"19",
          6215 => x"81",
          6216 => x"74",
          6217 => x"3f",
          6218 => x"08",
          6219 => x"98",
          6220 => x"7e",
          6221 => x"3f",
          6222 => x"08",
          6223 => x"d2",
          6224 => x"84",
          6225 => x"89",
          6226 => x"78",
          6227 => x"d5",
          6228 => x"7f",
          6229 => x"58",
          6230 => x"75",
          6231 => x"75",
          6232 => x"78",
          6233 => x"7c",
          6234 => x"33",
          6235 => x"3f",
          6236 => x"08",
          6237 => x"7e",
          6238 => x"78",
          6239 => x"74",
          6240 => x"38",
          6241 => x"b0",
          6242 => x"31",
          6243 => x"05",
          6244 => x"51",
          6245 => x"7e",
          6246 => x"83",
          6247 => x"89",
          6248 => x"db",
          6249 => x"08",
          6250 => x"26",
          6251 => x"51",
          6252 => x"82",
          6253 => x"fd",
          6254 => x"77",
          6255 => x"55",
          6256 => x"0c",
          6257 => x"83",
          6258 => x"80",
          6259 => x"55",
          6260 => x"83",
          6261 => x"9c",
          6262 => x"7e",
          6263 => x"3f",
          6264 => x"08",
          6265 => x"75",
          6266 => x"94",
          6267 => x"ff",
          6268 => x"05",
          6269 => x"3f",
          6270 => x"0b",
          6271 => x"7b",
          6272 => x"08",
          6273 => x"76",
          6274 => x"08",
          6275 => x"1c",
          6276 => x"08",
          6277 => x"5c",
          6278 => x"83",
          6279 => x"74",
          6280 => x"fd",
          6281 => x"18",
          6282 => x"07",
          6283 => x"19",
          6284 => x"75",
          6285 => x"0c",
          6286 => x"04",
          6287 => x"7a",
          6288 => x"05",
          6289 => x"56",
          6290 => x"82",
          6291 => x"57",
          6292 => x"08",
          6293 => x"90",
          6294 => x"86",
          6295 => x"06",
          6296 => x"73",
          6297 => x"e9",
          6298 => x"08",
          6299 => x"cc",
          6300 => x"93",
          6301 => x"82",
          6302 => x"80",
          6303 => x"16",
          6304 => x"33",
          6305 => x"55",
          6306 => x"34",
          6307 => x"53",
          6308 => x"08",
          6309 => x"3f",
          6310 => x"52",
          6311 => x"c9",
          6312 => x"88",
          6313 => x"96",
          6314 => x"f0",
          6315 => x"92",
          6316 => x"ca",
          6317 => x"81",
          6318 => x"34",
          6319 => x"df",
          6320 => x"84",
          6321 => x"33",
          6322 => x"55",
          6323 => x"17",
          6324 => x"93",
          6325 => x"3d",
          6326 => x"3d",
          6327 => x"52",
          6328 => x"3f",
          6329 => x"08",
          6330 => x"84",
          6331 => x"86",
          6332 => x"52",
          6333 => x"bc",
          6334 => x"84",
          6335 => x"93",
          6336 => x"38",
          6337 => x"08",
          6338 => x"82",
          6339 => x"86",
          6340 => x"ff",
          6341 => x"3d",
          6342 => x"3f",
          6343 => x"0b",
          6344 => x"08",
          6345 => x"82",
          6346 => x"82",
          6347 => x"80",
          6348 => x"93",
          6349 => x"3d",
          6350 => x"3d",
          6351 => x"93",
          6352 => x"52",
          6353 => x"e9",
          6354 => x"93",
          6355 => x"82",
          6356 => x"80",
          6357 => x"58",
          6358 => x"3d",
          6359 => x"e0",
          6360 => x"93",
          6361 => x"82",
          6362 => x"bc",
          6363 => x"c7",
          6364 => x"98",
          6365 => x"73",
          6366 => x"38",
          6367 => x"12",
          6368 => x"39",
          6369 => x"33",
          6370 => x"70",
          6371 => x"55",
          6372 => x"2e",
          6373 => x"7f",
          6374 => x"54",
          6375 => x"82",
          6376 => x"94",
          6377 => x"39",
          6378 => x"08",
          6379 => x"81",
          6380 => x"85",
          6381 => x"93",
          6382 => x"3d",
          6383 => x"3d",
          6384 => x"5b",
          6385 => x"34",
          6386 => x"3d",
          6387 => x"52",
          6388 => x"e8",
          6389 => x"93",
          6390 => x"82",
          6391 => x"82",
          6392 => x"43",
          6393 => x"11",
          6394 => x"58",
          6395 => x"80",
          6396 => x"38",
          6397 => x"3d",
          6398 => x"d5",
          6399 => x"93",
          6400 => x"82",
          6401 => x"82",
          6402 => x"52",
          6403 => x"c8",
          6404 => x"84",
          6405 => x"93",
          6406 => x"c1",
          6407 => x"7b",
          6408 => x"3f",
          6409 => x"08",
          6410 => x"74",
          6411 => x"3f",
          6412 => x"08",
          6413 => x"84",
          6414 => x"38",
          6415 => x"51",
          6416 => x"82",
          6417 => x"57",
          6418 => x"08",
          6419 => x"52",
          6420 => x"f2",
          6421 => x"93",
          6422 => x"a6",
          6423 => x"74",
          6424 => x"3f",
          6425 => x"08",
          6426 => x"84",
          6427 => x"cc",
          6428 => x"2e",
          6429 => x"86",
          6430 => x"81",
          6431 => x"81",
          6432 => x"3d",
          6433 => x"52",
          6434 => x"c9",
          6435 => x"3d",
          6436 => x"11",
          6437 => x"5a",
          6438 => x"2e",
          6439 => x"b9",
          6440 => x"16",
          6441 => x"33",
          6442 => x"73",
          6443 => x"16",
          6444 => x"26",
          6445 => x"75",
          6446 => x"38",
          6447 => x"05",
          6448 => x"6f",
          6449 => x"ff",
          6450 => x"55",
          6451 => x"74",
          6452 => x"38",
          6453 => x"11",
          6454 => x"74",
          6455 => x"39",
          6456 => x"09",
          6457 => x"38",
          6458 => x"11",
          6459 => x"74",
          6460 => x"82",
          6461 => x"70",
          6462 => x"ff",
          6463 => x"08",
          6464 => x"5c",
          6465 => x"73",
          6466 => x"38",
          6467 => x"1a",
          6468 => x"55",
          6469 => x"38",
          6470 => x"73",
          6471 => x"38",
          6472 => x"76",
          6473 => x"74",
          6474 => x"33",
          6475 => x"05",
          6476 => x"15",
          6477 => x"ba",
          6478 => x"05",
          6479 => x"ff",
          6480 => x"06",
          6481 => x"57",
          6482 => x"18",
          6483 => x"54",
          6484 => x"70",
          6485 => x"34",
          6486 => x"ee",
          6487 => x"34",
          6488 => x"84",
          6489 => x"0d",
          6490 => x"0d",
          6491 => x"3d",
          6492 => x"71",
          6493 => x"ec",
          6494 => x"93",
          6495 => x"82",
          6496 => x"82",
          6497 => x"15",
          6498 => x"82",
          6499 => x"15",
          6500 => x"76",
          6501 => x"90",
          6502 => x"81",
          6503 => x"06",
          6504 => x"72",
          6505 => x"56",
          6506 => x"54",
          6507 => x"17",
          6508 => x"78",
          6509 => x"38",
          6510 => x"22",
          6511 => x"59",
          6512 => x"78",
          6513 => x"76",
          6514 => x"51",
          6515 => x"3f",
          6516 => x"08",
          6517 => x"54",
          6518 => x"53",
          6519 => x"3f",
          6520 => x"08",
          6521 => x"38",
          6522 => x"75",
          6523 => x"18",
          6524 => x"31",
          6525 => x"57",
          6526 => x"b1",
          6527 => x"08",
          6528 => x"38",
          6529 => x"51",
          6530 => x"82",
          6531 => x"54",
          6532 => x"08",
          6533 => x"9a",
          6534 => x"84",
          6535 => x"81",
          6536 => x"93",
          6537 => x"16",
          6538 => x"16",
          6539 => x"2e",
          6540 => x"76",
          6541 => x"dc",
          6542 => x"31",
          6543 => x"18",
          6544 => x"90",
          6545 => x"81",
          6546 => x"06",
          6547 => x"56",
          6548 => x"9a",
          6549 => x"74",
          6550 => x"3f",
          6551 => x"08",
          6552 => x"84",
          6553 => x"82",
          6554 => x"56",
          6555 => x"52",
          6556 => x"84",
          6557 => x"84",
          6558 => x"ff",
          6559 => x"81",
          6560 => x"38",
          6561 => x"98",
          6562 => x"a6",
          6563 => x"16",
          6564 => x"39",
          6565 => x"16",
          6566 => x"75",
          6567 => x"53",
          6568 => x"aa",
          6569 => x"79",
          6570 => x"3f",
          6571 => x"08",
          6572 => x"0b",
          6573 => x"82",
          6574 => x"39",
          6575 => x"16",
          6576 => x"bb",
          6577 => x"2a",
          6578 => x"08",
          6579 => x"15",
          6580 => x"15",
          6581 => x"90",
          6582 => x"16",
          6583 => x"33",
          6584 => x"53",
          6585 => x"34",
          6586 => x"06",
          6587 => x"2e",
          6588 => x"9c",
          6589 => x"85",
          6590 => x"16",
          6591 => x"72",
          6592 => x"0c",
          6593 => x"04",
          6594 => x"79",
          6595 => x"75",
          6596 => x"8a",
          6597 => x"89",
          6598 => x"52",
          6599 => x"05",
          6600 => x"3f",
          6601 => x"08",
          6602 => x"84",
          6603 => x"38",
          6604 => x"7a",
          6605 => x"d8",
          6606 => x"93",
          6607 => x"82",
          6608 => x"80",
          6609 => x"16",
          6610 => x"2b",
          6611 => x"74",
          6612 => x"86",
          6613 => x"84",
          6614 => x"06",
          6615 => x"73",
          6616 => x"38",
          6617 => x"52",
          6618 => x"da",
          6619 => x"84",
          6620 => x"0c",
          6621 => x"14",
          6622 => x"23",
          6623 => x"51",
          6624 => x"82",
          6625 => x"55",
          6626 => x"09",
          6627 => x"38",
          6628 => x"39",
          6629 => x"84",
          6630 => x"0c",
          6631 => x"82",
          6632 => x"89",
          6633 => x"fc",
          6634 => x"87",
          6635 => x"53",
          6636 => x"e7",
          6637 => x"93",
          6638 => x"38",
          6639 => x"08",
          6640 => x"3d",
          6641 => x"3d",
          6642 => x"89",
          6643 => x"54",
          6644 => x"54",
          6645 => x"82",
          6646 => x"53",
          6647 => x"08",
          6648 => x"74",
          6649 => x"93",
          6650 => x"73",
          6651 => x"3f",
          6652 => x"08",
          6653 => x"39",
          6654 => x"08",
          6655 => x"d3",
          6656 => x"93",
          6657 => x"82",
          6658 => x"84",
          6659 => x"06",
          6660 => x"53",
          6661 => x"93",
          6662 => x"38",
          6663 => x"51",
          6664 => x"72",
          6665 => x"cf",
          6666 => x"93",
          6667 => x"32",
          6668 => x"72",
          6669 => x"70",
          6670 => x"08",
          6671 => x"54",
          6672 => x"93",
          6673 => x"3d",
          6674 => x"3d",
          6675 => x"80",
          6676 => x"70",
          6677 => x"52",
          6678 => x"3f",
          6679 => x"08",
          6680 => x"84",
          6681 => x"64",
          6682 => x"d6",
          6683 => x"93",
          6684 => x"82",
          6685 => x"a0",
          6686 => x"cb",
          6687 => x"98",
          6688 => x"73",
          6689 => x"38",
          6690 => x"39",
          6691 => x"88",
          6692 => x"75",
          6693 => x"3f",
          6694 => x"84",
          6695 => x"0d",
          6696 => x"0d",
          6697 => x"5c",
          6698 => x"3d",
          6699 => x"93",
          6700 => x"d6",
          6701 => x"84",
          6702 => x"93",
          6703 => x"80",
          6704 => x"0c",
          6705 => x"11",
          6706 => x"90",
          6707 => x"56",
          6708 => x"74",
          6709 => x"75",
          6710 => x"e4",
          6711 => x"81",
          6712 => x"5b",
          6713 => x"82",
          6714 => x"75",
          6715 => x"73",
          6716 => x"81",
          6717 => x"82",
          6718 => x"76",
          6719 => x"f0",
          6720 => x"f4",
          6721 => x"84",
          6722 => x"d1",
          6723 => x"84",
          6724 => x"ce",
          6725 => x"84",
          6726 => x"82",
          6727 => x"07",
          6728 => x"05",
          6729 => x"53",
          6730 => x"98",
          6731 => x"26",
          6732 => x"f9",
          6733 => x"08",
          6734 => x"08",
          6735 => x"98",
          6736 => x"81",
          6737 => x"58",
          6738 => x"3f",
          6739 => x"08",
          6740 => x"84",
          6741 => x"38",
          6742 => x"77",
          6743 => x"5d",
          6744 => x"74",
          6745 => x"81",
          6746 => x"b4",
          6747 => x"bb",
          6748 => x"93",
          6749 => x"ff",
          6750 => x"30",
          6751 => x"1b",
          6752 => x"5b",
          6753 => x"39",
          6754 => x"ff",
          6755 => x"82",
          6756 => x"f0",
          6757 => x"30",
          6758 => x"1b",
          6759 => x"5b",
          6760 => x"83",
          6761 => x"58",
          6762 => x"92",
          6763 => x"0c",
          6764 => x"12",
          6765 => x"33",
          6766 => x"54",
          6767 => x"34",
          6768 => x"84",
          6769 => x"0d",
          6770 => x"0d",
          6771 => x"fc",
          6772 => x"52",
          6773 => x"3f",
          6774 => x"08",
          6775 => x"84",
          6776 => x"38",
          6777 => x"56",
          6778 => x"38",
          6779 => x"70",
          6780 => x"81",
          6781 => x"55",
          6782 => x"80",
          6783 => x"38",
          6784 => x"54",
          6785 => x"08",
          6786 => x"38",
          6787 => x"82",
          6788 => x"53",
          6789 => x"52",
          6790 => x"8c",
          6791 => x"84",
          6792 => x"19",
          6793 => x"c9",
          6794 => x"08",
          6795 => x"ff",
          6796 => x"82",
          6797 => x"ff",
          6798 => x"06",
          6799 => x"56",
          6800 => x"08",
          6801 => x"81",
          6802 => x"82",
          6803 => x"75",
          6804 => x"54",
          6805 => x"08",
          6806 => x"27",
          6807 => x"17",
          6808 => x"93",
          6809 => x"76",
          6810 => x"3f",
          6811 => x"08",
          6812 => x"08",
          6813 => x"90",
          6814 => x"c0",
          6815 => x"90",
          6816 => x"80",
          6817 => x"75",
          6818 => x"75",
          6819 => x"93",
          6820 => x"3d",
          6821 => x"3d",
          6822 => x"a0",
          6823 => x"05",
          6824 => x"51",
          6825 => x"82",
          6826 => x"55",
          6827 => x"08",
          6828 => x"78",
          6829 => x"08",
          6830 => x"70",
          6831 => x"ae",
          6832 => x"84",
          6833 => x"93",
          6834 => x"db",
          6835 => x"fb",
          6836 => x"85",
          6837 => x"06",
          6838 => x"86",
          6839 => x"c7",
          6840 => x"2b",
          6841 => x"24",
          6842 => x"02",
          6843 => x"33",
          6844 => x"58",
          6845 => x"76",
          6846 => x"6b",
          6847 => x"cc",
          6848 => x"93",
          6849 => x"84",
          6850 => x"06",
          6851 => x"73",
          6852 => x"d4",
          6853 => x"82",
          6854 => x"94",
          6855 => x"81",
          6856 => x"5a",
          6857 => x"08",
          6858 => x"8a",
          6859 => x"54",
          6860 => x"82",
          6861 => x"55",
          6862 => x"08",
          6863 => x"82",
          6864 => x"52",
          6865 => x"e5",
          6866 => x"84",
          6867 => x"93",
          6868 => x"38",
          6869 => x"cf",
          6870 => x"84",
          6871 => x"88",
          6872 => x"84",
          6873 => x"38",
          6874 => x"c2",
          6875 => x"84",
          6876 => x"84",
          6877 => x"82",
          6878 => x"07",
          6879 => x"55",
          6880 => x"2e",
          6881 => x"80",
          6882 => x"80",
          6883 => x"77",
          6884 => x"3f",
          6885 => x"08",
          6886 => x"38",
          6887 => x"ba",
          6888 => x"93",
          6889 => x"74",
          6890 => x"0c",
          6891 => x"04",
          6892 => x"82",
          6893 => x"c0",
          6894 => x"3d",
          6895 => x"3f",
          6896 => x"08",
          6897 => x"84",
          6898 => x"38",
          6899 => x"52",
          6900 => x"52",
          6901 => x"3f",
          6902 => x"08",
          6903 => x"84",
          6904 => x"88",
          6905 => x"39",
          6906 => x"08",
          6907 => x"81",
          6908 => x"38",
          6909 => x"05",
          6910 => x"2a",
          6911 => x"55",
          6912 => x"81",
          6913 => x"5a",
          6914 => x"3d",
          6915 => x"c1",
          6916 => x"93",
          6917 => x"55",
          6918 => x"84",
          6919 => x"87",
          6920 => x"84",
          6921 => x"09",
          6922 => x"38",
          6923 => x"93",
          6924 => x"2e",
          6925 => x"86",
          6926 => x"81",
          6927 => x"81",
          6928 => x"93",
          6929 => x"78",
          6930 => x"3f",
          6931 => x"08",
          6932 => x"84",
          6933 => x"38",
          6934 => x"52",
          6935 => x"ff",
          6936 => x"78",
          6937 => x"b4",
          6938 => x"54",
          6939 => x"15",
          6940 => x"b2",
          6941 => x"ca",
          6942 => x"b6",
          6943 => x"53",
          6944 => x"53",
          6945 => x"3f",
          6946 => x"b4",
          6947 => x"d4",
          6948 => x"b6",
          6949 => x"54",
          6950 => x"d5",
          6951 => x"53",
          6952 => x"11",
          6953 => x"d7",
          6954 => x"81",
          6955 => x"34",
          6956 => x"a4",
          6957 => x"84",
          6958 => x"93",
          6959 => x"38",
          6960 => x"0a",
          6961 => x"05",
          6962 => x"d0",
          6963 => x"64",
          6964 => x"c9",
          6965 => x"54",
          6966 => x"15",
          6967 => x"81",
          6968 => x"34",
          6969 => x"b8",
          6970 => x"93",
          6971 => x"8b",
          6972 => x"75",
          6973 => x"ff",
          6974 => x"73",
          6975 => x"0c",
          6976 => x"04",
          6977 => x"a9",
          6978 => x"51",
          6979 => x"82",
          6980 => x"ff",
          6981 => x"a9",
          6982 => x"ee",
          6983 => x"84",
          6984 => x"93",
          6985 => x"d3",
          6986 => x"a9",
          6987 => x"9d",
          6988 => x"58",
          6989 => x"82",
          6990 => x"55",
          6991 => x"08",
          6992 => x"02",
          6993 => x"33",
          6994 => x"54",
          6995 => x"82",
          6996 => x"53",
          6997 => x"52",
          6998 => x"88",
          6999 => x"b4",
          7000 => x"53",
          7001 => x"3d",
          7002 => x"ff",
          7003 => x"aa",
          7004 => x"73",
          7005 => x"3f",
          7006 => x"08",
          7007 => x"84",
          7008 => x"63",
          7009 => x"81",
          7010 => x"65",
          7011 => x"2e",
          7012 => x"55",
          7013 => x"82",
          7014 => x"84",
          7015 => x"06",
          7016 => x"73",
          7017 => x"3f",
          7018 => x"08",
          7019 => x"84",
          7020 => x"38",
          7021 => x"53",
          7022 => x"95",
          7023 => x"16",
          7024 => x"87",
          7025 => x"05",
          7026 => x"34",
          7027 => x"70",
          7028 => x"81",
          7029 => x"55",
          7030 => x"74",
          7031 => x"73",
          7032 => x"78",
          7033 => x"83",
          7034 => x"16",
          7035 => x"2a",
          7036 => x"51",
          7037 => x"80",
          7038 => x"38",
          7039 => x"80",
          7040 => x"52",
          7041 => x"be",
          7042 => x"84",
          7043 => x"51",
          7044 => x"3f",
          7045 => x"93",
          7046 => x"2e",
          7047 => x"82",
          7048 => x"52",
          7049 => x"b5",
          7050 => x"93",
          7051 => x"80",
          7052 => x"58",
          7053 => x"84",
          7054 => x"38",
          7055 => x"54",
          7056 => x"09",
          7057 => x"38",
          7058 => x"52",
          7059 => x"af",
          7060 => x"81",
          7061 => x"34",
          7062 => x"93",
          7063 => x"38",
          7064 => x"ca",
          7065 => x"84",
          7066 => x"93",
          7067 => x"38",
          7068 => x"b5",
          7069 => x"93",
          7070 => x"74",
          7071 => x"0c",
          7072 => x"04",
          7073 => x"02",
          7074 => x"33",
          7075 => x"80",
          7076 => x"57",
          7077 => x"95",
          7078 => x"52",
          7079 => x"d2",
          7080 => x"93",
          7081 => x"82",
          7082 => x"80",
          7083 => x"5a",
          7084 => x"3d",
          7085 => x"c9",
          7086 => x"93",
          7087 => x"82",
          7088 => x"b8",
          7089 => x"cf",
          7090 => x"a0",
          7091 => x"55",
          7092 => x"75",
          7093 => x"71",
          7094 => x"33",
          7095 => x"74",
          7096 => x"57",
          7097 => x"8b",
          7098 => x"54",
          7099 => x"15",
          7100 => x"ff",
          7101 => x"82",
          7102 => x"55",
          7103 => x"84",
          7104 => x"0d",
          7105 => x"0d",
          7106 => x"53",
          7107 => x"05",
          7108 => x"51",
          7109 => x"82",
          7110 => x"55",
          7111 => x"08",
          7112 => x"76",
          7113 => x"93",
          7114 => x"51",
          7115 => x"82",
          7116 => x"55",
          7117 => x"08",
          7118 => x"80",
          7119 => x"81",
          7120 => x"86",
          7121 => x"38",
          7122 => x"86",
          7123 => x"90",
          7124 => x"54",
          7125 => x"ff",
          7126 => x"76",
          7127 => x"83",
          7128 => x"51",
          7129 => x"3f",
          7130 => x"08",
          7131 => x"93",
          7132 => x"3d",
          7133 => x"3d",
          7134 => x"5c",
          7135 => x"98",
          7136 => x"52",
          7137 => x"d1",
          7138 => x"93",
          7139 => x"93",
          7140 => x"70",
          7141 => x"08",
          7142 => x"51",
          7143 => x"80",
          7144 => x"38",
          7145 => x"06",
          7146 => x"80",
          7147 => x"38",
          7148 => x"5f",
          7149 => x"3d",
          7150 => x"ff",
          7151 => x"82",
          7152 => x"57",
          7153 => x"08",
          7154 => x"74",
          7155 => x"c3",
          7156 => x"93",
          7157 => x"82",
          7158 => x"bf",
          7159 => x"84",
          7160 => x"84",
          7161 => x"59",
          7162 => x"81",
          7163 => x"56",
          7164 => x"33",
          7165 => x"16",
          7166 => x"27",
          7167 => x"56",
          7168 => x"80",
          7169 => x"80",
          7170 => x"ff",
          7171 => x"70",
          7172 => x"56",
          7173 => x"e8",
          7174 => x"76",
          7175 => x"81",
          7176 => x"80",
          7177 => x"57",
          7178 => x"78",
          7179 => x"51",
          7180 => x"2e",
          7181 => x"73",
          7182 => x"38",
          7183 => x"08",
          7184 => x"b1",
          7185 => x"93",
          7186 => x"82",
          7187 => x"a7",
          7188 => x"33",
          7189 => x"c3",
          7190 => x"2e",
          7191 => x"e4",
          7192 => x"2e",
          7193 => x"56",
          7194 => x"05",
          7195 => x"e3",
          7196 => x"84",
          7197 => x"76",
          7198 => x"0c",
          7199 => x"04",
          7200 => x"82",
          7201 => x"ff",
          7202 => x"9d",
          7203 => x"fa",
          7204 => x"84",
          7205 => x"84",
          7206 => x"82",
          7207 => x"83",
          7208 => x"53",
          7209 => x"3d",
          7210 => x"ff",
          7211 => x"73",
          7212 => x"70",
          7213 => x"52",
          7214 => x"9f",
          7215 => x"bc",
          7216 => x"74",
          7217 => x"6d",
          7218 => x"70",
          7219 => x"af",
          7220 => x"93",
          7221 => x"2e",
          7222 => x"70",
          7223 => x"57",
          7224 => x"fd",
          7225 => x"84",
          7226 => x"8d",
          7227 => x"2b",
          7228 => x"81",
          7229 => x"86",
          7230 => x"84",
          7231 => x"9f",
          7232 => x"ff",
          7233 => x"54",
          7234 => x"8a",
          7235 => x"70",
          7236 => x"06",
          7237 => x"ff",
          7238 => x"38",
          7239 => x"15",
          7240 => x"80",
          7241 => x"74",
          7242 => x"f0",
          7243 => x"89",
          7244 => x"84",
          7245 => x"81",
          7246 => x"88",
          7247 => x"26",
          7248 => x"39",
          7249 => x"86",
          7250 => x"81",
          7251 => x"ff",
          7252 => x"38",
          7253 => x"54",
          7254 => x"81",
          7255 => x"81",
          7256 => x"78",
          7257 => x"5a",
          7258 => x"6d",
          7259 => x"81",
          7260 => x"57",
          7261 => x"9f",
          7262 => x"38",
          7263 => x"54",
          7264 => x"81",
          7265 => x"b1",
          7266 => x"2e",
          7267 => x"a7",
          7268 => x"15",
          7269 => x"54",
          7270 => x"09",
          7271 => x"38",
          7272 => x"76",
          7273 => x"41",
          7274 => x"52",
          7275 => x"52",
          7276 => x"b3",
          7277 => x"84",
          7278 => x"93",
          7279 => x"f7",
          7280 => x"74",
          7281 => x"e5",
          7282 => x"84",
          7283 => x"93",
          7284 => x"38",
          7285 => x"38",
          7286 => x"74",
          7287 => x"39",
          7288 => x"08",
          7289 => x"81",
          7290 => x"38",
          7291 => x"74",
          7292 => x"38",
          7293 => x"51",
          7294 => x"3f",
          7295 => x"08",
          7296 => x"84",
          7297 => x"a0",
          7298 => x"84",
          7299 => x"51",
          7300 => x"3f",
          7301 => x"0b",
          7302 => x"8b",
          7303 => x"67",
          7304 => x"a7",
          7305 => x"81",
          7306 => x"34",
          7307 => x"ad",
          7308 => x"93",
          7309 => x"73",
          7310 => x"93",
          7311 => x"3d",
          7312 => x"3d",
          7313 => x"02",
          7314 => x"cb",
          7315 => x"3d",
          7316 => x"72",
          7317 => x"5a",
          7318 => x"82",
          7319 => x"58",
          7320 => x"08",
          7321 => x"91",
          7322 => x"77",
          7323 => x"7c",
          7324 => x"38",
          7325 => x"59",
          7326 => x"90",
          7327 => x"81",
          7328 => x"06",
          7329 => x"73",
          7330 => x"54",
          7331 => x"82",
          7332 => x"39",
          7333 => x"8b",
          7334 => x"11",
          7335 => x"2b",
          7336 => x"54",
          7337 => x"fe",
          7338 => x"ff",
          7339 => x"70",
          7340 => x"07",
          7341 => x"93",
          7342 => x"8c",
          7343 => x"40",
          7344 => x"55",
          7345 => x"88",
          7346 => x"08",
          7347 => x"38",
          7348 => x"77",
          7349 => x"56",
          7350 => x"51",
          7351 => x"3f",
          7352 => x"55",
          7353 => x"08",
          7354 => x"38",
          7355 => x"93",
          7356 => x"2e",
          7357 => x"82",
          7358 => x"ff",
          7359 => x"38",
          7360 => x"08",
          7361 => x"16",
          7362 => x"2e",
          7363 => x"87",
          7364 => x"74",
          7365 => x"74",
          7366 => x"81",
          7367 => x"38",
          7368 => x"ff",
          7369 => x"2e",
          7370 => x"7b",
          7371 => x"80",
          7372 => x"81",
          7373 => x"81",
          7374 => x"06",
          7375 => x"56",
          7376 => x"52",
          7377 => x"af",
          7378 => x"93",
          7379 => x"82",
          7380 => x"80",
          7381 => x"81",
          7382 => x"56",
          7383 => x"d3",
          7384 => x"ff",
          7385 => x"7c",
          7386 => x"55",
          7387 => x"b3",
          7388 => x"1b",
          7389 => x"1b",
          7390 => x"33",
          7391 => x"54",
          7392 => x"34",
          7393 => x"fe",
          7394 => x"08",
          7395 => x"74",
          7396 => x"75",
          7397 => x"16",
          7398 => x"33",
          7399 => x"73",
          7400 => x"77",
          7401 => x"93",
          7402 => x"3d",
          7403 => x"3d",
          7404 => x"02",
          7405 => x"eb",
          7406 => x"3d",
          7407 => x"59",
          7408 => x"8b",
          7409 => x"82",
          7410 => x"24",
          7411 => x"82",
          7412 => x"84",
          7413 => x"b4",
          7414 => x"51",
          7415 => x"2e",
          7416 => x"75",
          7417 => x"84",
          7418 => x"06",
          7419 => x"7e",
          7420 => x"d0",
          7421 => x"84",
          7422 => x"06",
          7423 => x"56",
          7424 => x"74",
          7425 => x"76",
          7426 => x"81",
          7427 => x"8a",
          7428 => x"b2",
          7429 => x"fc",
          7430 => x"52",
          7431 => x"a4",
          7432 => x"93",
          7433 => x"38",
          7434 => x"80",
          7435 => x"74",
          7436 => x"26",
          7437 => x"15",
          7438 => x"74",
          7439 => x"38",
          7440 => x"80",
          7441 => x"84",
          7442 => x"92",
          7443 => x"80",
          7444 => x"38",
          7445 => x"06",
          7446 => x"2e",
          7447 => x"56",
          7448 => x"78",
          7449 => x"89",
          7450 => x"2b",
          7451 => x"43",
          7452 => x"38",
          7453 => x"30",
          7454 => x"77",
          7455 => x"91",
          7456 => x"c2",
          7457 => x"f8",
          7458 => x"52",
          7459 => x"a4",
          7460 => x"56",
          7461 => x"08",
          7462 => x"77",
          7463 => x"77",
          7464 => x"84",
          7465 => x"45",
          7466 => x"bf",
          7467 => x"8e",
          7468 => x"26",
          7469 => x"74",
          7470 => x"48",
          7471 => x"75",
          7472 => x"38",
          7473 => x"81",
          7474 => x"fa",
          7475 => x"2a",
          7476 => x"56",
          7477 => x"2e",
          7478 => x"87",
          7479 => x"82",
          7480 => x"38",
          7481 => x"55",
          7482 => x"83",
          7483 => x"81",
          7484 => x"56",
          7485 => x"80",
          7486 => x"38",
          7487 => x"83",
          7488 => x"06",
          7489 => x"78",
          7490 => x"91",
          7491 => x"0b",
          7492 => x"22",
          7493 => x"80",
          7494 => x"74",
          7495 => x"38",
          7496 => x"56",
          7497 => x"17",
          7498 => x"57",
          7499 => x"2e",
          7500 => x"75",
          7501 => x"79",
          7502 => x"fe",
          7503 => x"82",
          7504 => x"84",
          7505 => x"05",
          7506 => x"5e",
          7507 => x"80",
          7508 => x"84",
          7509 => x"8a",
          7510 => x"fd",
          7511 => x"75",
          7512 => x"38",
          7513 => x"78",
          7514 => x"8c",
          7515 => x"0b",
          7516 => x"22",
          7517 => x"80",
          7518 => x"74",
          7519 => x"38",
          7520 => x"56",
          7521 => x"17",
          7522 => x"57",
          7523 => x"2e",
          7524 => x"75",
          7525 => x"79",
          7526 => x"fe",
          7527 => x"82",
          7528 => x"10",
          7529 => x"82",
          7530 => x"9f",
          7531 => x"38",
          7532 => x"93",
          7533 => x"82",
          7534 => x"05",
          7535 => x"2a",
          7536 => x"56",
          7537 => x"17",
          7538 => x"81",
          7539 => x"60",
          7540 => x"65",
          7541 => x"12",
          7542 => x"30",
          7543 => x"74",
          7544 => x"59",
          7545 => x"7d",
          7546 => x"81",
          7547 => x"76",
          7548 => x"41",
          7549 => x"76",
          7550 => x"90",
          7551 => x"62",
          7552 => x"51",
          7553 => x"26",
          7554 => x"75",
          7555 => x"31",
          7556 => x"65",
          7557 => x"fe",
          7558 => x"82",
          7559 => x"58",
          7560 => x"09",
          7561 => x"38",
          7562 => x"08",
          7563 => x"26",
          7564 => x"78",
          7565 => x"79",
          7566 => x"78",
          7567 => x"86",
          7568 => x"82",
          7569 => x"06",
          7570 => x"83",
          7571 => x"82",
          7572 => x"27",
          7573 => x"8f",
          7574 => x"55",
          7575 => x"26",
          7576 => x"59",
          7577 => x"62",
          7578 => x"74",
          7579 => x"38",
          7580 => x"88",
          7581 => x"84",
          7582 => x"26",
          7583 => x"86",
          7584 => x"1a",
          7585 => x"79",
          7586 => x"38",
          7587 => x"80",
          7588 => x"2e",
          7589 => x"83",
          7590 => x"9f",
          7591 => x"8b",
          7592 => x"06",
          7593 => x"74",
          7594 => x"84",
          7595 => x"52",
          7596 => x"a2",
          7597 => x"53",
          7598 => x"52",
          7599 => x"a2",
          7600 => x"80",
          7601 => x"51",
          7602 => x"3f",
          7603 => x"34",
          7604 => x"ff",
          7605 => x"1b",
          7606 => x"a2",
          7607 => x"90",
          7608 => x"83",
          7609 => x"70",
          7610 => x"80",
          7611 => x"55",
          7612 => x"ff",
          7613 => x"66",
          7614 => x"ff",
          7615 => x"38",
          7616 => x"ff",
          7617 => x"1b",
          7618 => x"f2",
          7619 => x"74",
          7620 => x"51",
          7621 => x"3f",
          7622 => x"1c",
          7623 => x"98",
          7624 => x"a0",
          7625 => x"ff",
          7626 => x"51",
          7627 => x"3f",
          7628 => x"1b",
          7629 => x"e4",
          7630 => x"2e",
          7631 => x"80",
          7632 => x"88",
          7633 => x"80",
          7634 => x"ff",
          7635 => x"7c",
          7636 => x"51",
          7637 => x"3f",
          7638 => x"1b",
          7639 => x"bc",
          7640 => x"b0",
          7641 => x"a0",
          7642 => x"52",
          7643 => x"ff",
          7644 => x"ff",
          7645 => x"c0",
          7646 => x"0b",
          7647 => x"34",
          7648 => x"ff",
          7649 => x"c7",
          7650 => x"39",
          7651 => x"0a",
          7652 => x"51",
          7653 => x"3f",
          7654 => x"ff",
          7655 => x"1b",
          7656 => x"da",
          7657 => x"0b",
          7658 => x"a9",
          7659 => x"34",
          7660 => x"ff",
          7661 => x"1b",
          7662 => x"8f",
          7663 => x"d5",
          7664 => x"1b",
          7665 => x"ff",
          7666 => x"81",
          7667 => x"7a",
          7668 => x"ff",
          7669 => x"81",
          7670 => x"84",
          7671 => x"38",
          7672 => x"09",
          7673 => x"ee",
          7674 => x"60",
          7675 => x"7a",
          7676 => x"ff",
          7677 => x"84",
          7678 => x"52",
          7679 => x"9f",
          7680 => x"8b",
          7681 => x"52",
          7682 => x"9f",
          7683 => x"8a",
          7684 => x"52",
          7685 => x"51",
          7686 => x"3f",
          7687 => x"83",
          7688 => x"ff",
          7689 => x"82",
          7690 => x"1b",
          7691 => x"ec",
          7692 => x"d5",
          7693 => x"ff",
          7694 => x"75",
          7695 => x"05",
          7696 => x"7e",
          7697 => x"e5",
          7698 => x"60",
          7699 => x"52",
          7700 => x"9a",
          7701 => x"53",
          7702 => x"51",
          7703 => x"3f",
          7704 => x"58",
          7705 => x"09",
          7706 => x"38",
          7707 => x"51",
          7708 => x"3f",
          7709 => x"1b",
          7710 => x"a0",
          7711 => x"52",
          7712 => x"91",
          7713 => x"ff",
          7714 => x"81",
          7715 => x"f8",
          7716 => x"7a",
          7717 => x"84",
          7718 => x"61",
          7719 => x"26",
          7720 => x"57",
          7721 => x"53",
          7722 => x"51",
          7723 => x"3f",
          7724 => x"08",
          7725 => x"84",
          7726 => x"93",
          7727 => x"7a",
          7728 => x"aa",
          7729 => x"75",
          7730 => x"56",
          7731 => x"81",
          7732 => x"80",
          7733 => x"38",
          7734 => x"83",
          7735 => x"63",
          7736 => x"74",
          7737 => x"38",
          7738 => x"54",
          7739 => x"52",
          7740 => x"99",
          7741 => x"93",
          7742 => x"c1",
          7743 => x"75",
          7744 => x"56",
          7745 => x"8c",
          7746 => x"2e",
          7747 => x"56",
          7748 => x"ff",
          7749 => x"84",
          7750 => x"2e",
          7751 => x"56",
          7752 => x"58",
          7753 => x"38",
          7754 => x"77",
          7755 => x"ff",
          7756 => x"82",
          7757 => x"78",
          7758 => x"c2",
          7759 => x"1b",
          7760 => x"34",
          7761 => x"16",
          7762 => x"82",
          7763 => x"83",
          7764 => x"84",
          7765 => x"67",
          7766 => x"fd",
          7767 => x"51",
          7768 => x"3f",
          7769 => x"16",
          7770 => x"84",
          7771 => x"bf",
          7772 => x"86",
          7773 => x"93",
          7774 => x"16",
          7775 => x"83",
          7776 => x"ff",
          7777 => x"66",
          7778 => x"1b",
          7779 => x"8c",
          7780 => x"77",
          7781 => x"7e",
          7782 => x"91",
          7783 => x"82",
          7784 => x"a2",
          7785 => x"80",
          7786 => x"ff",
          7787 => x"81",
          7788 => x"84",
          7789 => x"89",
          7790 => x"8a",
          7791 => x"86",
          7792 => x"84",
          7793 => x"82",
          7794 => x"99",
          7795 => x"f5",
          7796 => x"60",
          7797 => x"79",
          7798 => x"5a",
          7799 => x"78",
          7800 => x"8d",
          7801 => x"55",
          7802 => x"fc",
          7803 => x"51",
          7804 => x"7a",
          7805 => x"81",
          7806 => x"8c",
          7807 => x"74",
          7808 => x"38",
          7809 => x"81",
          7810 => x"81",
          7811 => x"8a",
          7812 => x"06",
          7813 => x"76",
          7814 => x"76",
          7815 => x"55",
          7816 => x"84",
          7817 => x"0d",
          7818 => x"0d",
          7819 => x"05",
          7820 => x"59",
          7821 => x"2e",
          7822 => x"87",
          7823 => x"76",
          7824 => x"84",
          7825 => x"80",
          7826 => x"38",
          7827 => x"77",
          7828 => x"56",
          7829 => x"34",
          7830 => x"bb",
          7831 => x"38",
          7832 => x"05",
          7833 => x"8c",
          7834 => x"08",
          7835 => x"3f",
          7836 => x"70",
          7837 => x"07",
          7838 => x"30",
          7839 => x"56",
          7840 => x"0c",
          7841 => x"18",
          7842 => x"0d",
          7843 => x"0d",
          7844 => x"08",
          7845 => x"75",
          7846 => x"89",
          7847 => x"54",
          7848 => x"16",
          7849 => x"51",
          7850 => x"82",
          7851 => x"91",
          7852 => x"08",
          7853 => x"81",
          7854 => x"88",
          7855 => x"83",
          7856 => x"74",
          7857 => x"0c",
          7858 => x"04",
          7859 => x"75",
          7860 => x"53",
          7861 => x"51",
          7862 => x"3f",
          7863 => x"85",
          7864 => x"ea",
          7865 => x"80",
          7866 => x"6a",
          7867 => x"70",
          7868 => x"d8",
          7869 => x"72",
          7870 => x"3f",
          7871 => x"8d",
          7872 => x"0d",
          7873 => x"0d",
          7874 => x"70",
          7875 => x"74",
          7876 => x"e1",
          7877 => x"77",
          7878 => x"85",
          7879 => x"80",
          7880 => x"33",
          7881 => x"2e",
          7882 => x"86",
          7883 => x"55",
          7884 => x"57",
          7885 => x"82",
          7886 => x"70",
          7887 => x"fe",
          7888 => x"82",
          7889 => x"82",
          7890 => x"54",
          7891 => x"08",
          7892 => x"da",
          7893 => x"93",
          7894 => x"38",
          7895 => x"54",
          7896 => x"ff",
          7897 => x"17",
          7898 => x"06",
          7899 => x"77",
          7900 => x"ff",
          7901 => x"93",
          7902 => x"3d",
          7903 => x"3d",
          7904 => x"71",
          7905 => x"8e",
          7906 => x"29",
          7907 => x"05",
          7908 => x"04",
          7909 => x"51",
          7910 => x"82",
          7911 => x"80",
          7912 => x"82",
          7913 => x"f2",
          7914 => x"80",
          7915 => x"39",
          7916 => x"51",
          7917 => x"82",
          7918 => x"80",
          7919 => x"83",
          7920 => x"d6",
          7921 => x"c4",
          7922 => x"39",
          7923 => x"51",
          7924 => x"82",
          7925 => x"80",
          7926 => x"84",
          7927 => x"39",
          7928 => x"51",
          7929 => x"84",
          7930 => x"39",
          7931 => x"51",
          7932 => x"84",
          7933 => x"39",
          7934 => x"51",
          7935 => x"85",
          7936 => x"39",
          7937 => x"51",
          7938 => x"85",
          7939 => x"39",
          7940 => x"51",
          7941 => x"86",
          7942 => x"f2",
          7943 => x"3d",
          7944 => x"3d",
          7945 => x"56",
          7946 => x"e7",
          7947 => x"74",
          7948 => x"e8",
          7949 => x"39",
          7950 => x"74",
          7951 => x"9e",
          7952 => x"84",
          7953 => x"51",
          7954 => x"3f",
          7955 => x"08",
          7956 => x"75",
          7957 => x"94",
          7958 => x"d3",
          7959 => x"0d",
          7960 => x"0d",
          7961 => x"05",
          7962 => x"33",
          7963 => x"68",
          7964 => x"7a",
          7965 => x"51",
          7966 => x"78",
          7967 => x"ff",
          7968 => x"81",
          7969 => x"07",
          7970 => x"06",
          7971 => x"56",
          7972 => x"38",
          7973 => x"52",
          7974 => x"52",
          7975 => x"c9",
          7976 => x"84",
          7977 => x"93",
          7978 => x"38",
          7979 => x"08",
          7980 => x"88",
          7981 => x"84",
          7982 => x"3d",
          7983 => x"84",
          7984 => x"52",
          7985 => x"86",
          7986 => x"84",
          7987 => x"93",
          7988 => x"38",
          7989 => x"80",
          7990 => x"74",
          7991 => x"59",
          7992 => x"96",
          7993 => x"51",
          7994 => x"76",
          7995 => x"07",
          7996 => x"30",
          7997 => x"72",
          7998 => x"51",
          7999 => x"2e",
          8000 => x"86",
          8001 => x"c0",
          8002 => x"52",
          8003 => x"92",
          8004 => x"75",
          8005 => x"0c",
          8006 => x"04",
          8007 => x"7b",
          8008 => x"b3",
          8009 => x"58",
          8010 => x"53",
          8011 => x"51",
          8012 => x"82",
          8013 => x"a4",
          8014 => x"2e",
          8015 => x"81",
          8016 => x"98",
          8017 => x"7f",
          8018 => x"84",
          8019 => x"7d",
          8020 => x"82",
          8021 => x"57",
          8022 => x"04",
          8023 => x"84",
          8024 => x"0d",
          8025 => x"0d",
          8026 => x"02",
          8027 => x"cf",
          8028 => x"73",
          8029 => x"5f",
          8030 => x"5e",
          8031 => x"82",
          8032 => x"fe",
          8033 => x"82",
          8034 => x"fe",
          8035 => x"80",
          8036 => x"27",
          8037 => x"7b",
          8038 => x"38",
          8039 => x"a7",
          8040 => x"39",
          8041 => x"72",
          8042 => x"38",
          8043 => x"82",
          8044 => x"fe",
          8045 => x"89",
          8046 => x"d8",
          8047 => x"8b",
          8048 => x"55",
          8049 => x"74",
          8050 => x"7a",
          8051 => x"72",
          8052 => x"86",
          8053 => x"f4",
          8054 => x"39",
          8055 => x"51",
          8056 => x"3f",
          8057 => x"a1",
          8058 => x"53",
          8059 => x"8e",
          8060 => x"52",
          8061 => x"51",
          8062 => x"3f",
          8063 => x"86",
          8064 => x"ee",
          8065 => x"15",
          8066 => x"fe",
          8067 => x"ff",
          8068 => x"86",
          8069 => x"ee",
          8070 => x"55",
          8071 => x"bc",
          8072 => x"70",
          8073 => x"80",
          8074 => x"27",
          8075 => x"56",
          8076 => x"74",
          8077 => x"81",
          8078 => x"06",
          8079 => x"06",
          8080 => x"80",
          8081 => x"73",
          8082 => x"85",
          8083 => x"83",
          8084 => x"fe",
          8085 => x"81",
          8086 => x"39",
          8087 => x"51",
          8088 => x"3f",
          8089 => x"1c",
          8090 => x"de",
          8091 => x"93",
          8092 => x"2b",
          8093 => x"51",
          8094 => x"2e",
          8095 => x"ab",
          8096 => x"fd",
          8097 => x"84",
          8098 => x"70",
          8099 => x"a0",
          8100 => x"72",
          8101 => x"30",
          8102 => x"73",
          8103 => x"51",
          8104 => x"57",
          8105 => x"73",
          8106 => x"76",
          8107 => x"81",
          8108 => x"80",
          8109 => x"7c",
          8110 => x"78",
          8111 => x"38",
          8112 => x"82",
          8113 => x"8f",
          8114 => x"fc",
          8115 => x"9b",
          8116 => x"86",
          8117 => x"86",
          8118 => x"fe",
          8119 => x"82",
          8120 => x"51",
          8121 => x"3f",
          8122 => x"54",
          8123 => x"53",
          8124 => x"33",
          8125 => x"9c",
          8126 => x"b3",
          8127 => x"2e",
          8128 => x"e2",
          8129 => x"3d",
          8130 => x"3d",
          8131 => x"96",
          8132 => x"fe",
          8133 => x"81",
          8134 => x"f9",
          8135 => x"b8",
          8136 => x"f1",
          8137 => x"fe",
          8138 => x"72",
          8139 => x"81",
          8140 => x"71",
          8141 => x"38",
          8142 => x"d8",
          8143 => x"87",
          8144 => x"da",
          8145 => x"51",
          8146 => x"3f",
          8147 => x"70",
          8148 => x"52",
          8149 => x"95",
          8150 => x"fe",
          8151 => x"82",
          8152 => x"fe",
          8153 => x"80",
          8154 => x"a9",
          8155 => x"2a",
          8156 => x"51",
          8157 => x"2e",
          8158 => x"51",
          8159 => x"3f",
          8160 => x"51",
          8161 => x"3f",
          8162 => x"d8",
          8163 => x"84",
          8164 => x"06",
          8165 => x"80",
          8166 => x"81",
          8167 => x"f5",
          8168 => x"8c",
          8169 => x"ed",
          8170 => x"fe",
          8171 => x"72",
          8172 => x"81",
          8173 => x"71",
          8174 => x"38",
          8175 => x"d7",
          8176 => x"88",
          8177 => x"d9",
          8178 => x"51",
          8179 => x"3f",
          8180 => x"70",
          8181 => x"52",
          8182 => x"95",
          8183 => x"fe",
          8184 => x"82",
          8185 => x"fe",
          8186 => x"80",
          8187 => x"a5",
          8188 => x"2a",
          8189 => x"51",
          8190 => x"2e",
          8191 => x"51",
          8192 => x"3f",
          8193 => x"51",
          8194 => x"3f",
          8195 => x"d7",
          8196 => x"88",
          8197 => x"06",
          8198 => x"80",
          8199 => x"81",
          8200 => x"f1",
          8201 => x"dc",
          8202 => x"e9",
          8203 => x"fe",
          8204 => x"fe",
          8205 => x"84",
          8206 => x"fb",
          8207 => x"02",
          8208 => x"05",
          8209 => x"56",
          8210 => x"75",
          8211 => x"a1",
          8212 => x"f0",
          8213 => x"a7",
          8214 => x"82",
          8215 => x"82",
          8216 => x"ff",
          8217 => x"82",
          8218 => x"30",
          8219 => x"84",
          8220 => x"25",
          8221 => x"51",
          8222 => x"82",
          8223 => x"82",
          8224 => x"54",
          8225 => x"09",
          8226 => x"38",
          8227 => x"53",
          8228 => x"51",
          8229 => x"82",
          8230 => x"80",
          8231 => x"82",
          8232 => x"51",
          8233 => x"3f",
          8234 => x"aa",
          8235 => x"aa",
          8236 => x"82",
          8237 => x"82",
          8238 => x"54",
          8239 => x"09",
          8240 => x"38",
          8241 => x"51",
          8242 => x"3f",
          8243 => x"93",
          8244 => x"3d",
          8245 => x"3d",
          8246 => x"71",
          8247 => x"0c",
          8248 => x"52",
          8249 => x"86",
          8250 => x"93",
          8251 => x"ff",
          8252 => x"7d",
          8253 => x"06",
          8254 => x"89",
          8255 => x"3d",
          8256 => x"fe",
          8257 => x"7c",
          8258 => x"82",
          8259 => x"ff",
          8260 => x"82",
          8261 => x"7d",
          8262 => x"82",
          8263 => x"91",
          8264 => x"70",
          8265 => x"89",
          8266 => x"e8",
          8267 => x"3d",
          8268 => x"80",
          8269 => x"51",
          8270 => x"b4",
          8271 => x"05",
          8272 => x"3f",
          8273 => x"08",
          8274 => x"90",
          8275 => x"78",
          8276 => x"89",
          8277 => x"80",
          8278 => x"d9",
          8279 => x"2e",
          8280 => x"78",
          8281 => x"38",
          8282 => x"81",
          8283 => x"82",
          8284 => x"78",
          8285 => x"ae",
          8286 => x"39",
          8287 => x"82",
          8288 => x"94",
          8289 => x"38",
          8290 => x"78",
          8291 => x"8c",
          8292 => x"24",
          8293 => x"b0",
          8294 => x"38",
          8295 => x"84",
          8296 => x"fc",
          8297 => x"2e",
          8298 => x"78",
          8299 => x"86",
          8300 => x"ec",
          8301 => x"d5",
          8302 => x"38",
          8303 => x"24",
          8304 => x"80",
          8305 => x"f6",
          8306 => x"d0",
          8307 => x"78",
          8308 => x"8a",
          8309 => x"80",
          8310 => x"c2",
          8311 => x"39",
          8312 => x"2e",
          8313 => x"78",
          8314 => x"8c",
          8315 => x"b0",
          8316 => x"82",
          8317 => x"38",
          8318 => x"24",
          8319 => x"80",
          8320 => x"96",
          8321 => x"f9",
          8322 => x"38",
          8323 => x"78",
          8324 => x"8d",
          8325 => x"81",
          8326 => x"fd",
          8327 => x"39",
          8328 => x"80",
          8329 => x"84",
          8330 => x"ed",
          8331 => x"93",
          8332 => x"38",
          8333 => x"51",
          8334 => x"b4",
          8335 => x"11",
          8336 => x"05",
          8337 => x"dc",
          8338 => x"84",
          8339 => x"88",
          8340 => x"25",
          8341 => x"43",
          8342 => x"05",
          8343 => x"80",
          8344 => x"51",
          8345 => x"3f",
          8346 => x"08",
          8347 => x"59",
          8348 => x"82",
          8349 => x"fe",
          8350 => x"81",
          8351 => x"39",
          8352 => x"51",
          8353 => x"b4",
          8354 => x"11",
          8355 => x"05",
          8356 => x"90",
          8357 => x"84",
          8358 => x"fd",
          8359 => x"53",
          8360 => x"80",
          8361 => x"51",
          8362 => x"3f",
          8363 => x"08",
          8364 => x"a4",
          8365 => x"39",
          8366 => x"80",
          8367 => x"84",
          8368 => x"ec",
          8369 => x"93",
          8370 => x"2e",
          8371 => x"89",
          8372 => x"38",
          8373 => x"fc",
          8374 => x"84",
          8375 => x"ec",
          8376 => x"93",
          8377 => x"38",
          8378 => x"08",
          8379 => x"82",
          8380 => x"79",
          8381 => x"cd",
          8382 => x"cb",
          8383 => x"79",
          8384 => x"b4",
          8385 => x"c8",
          8386 => x"b1",
          8387 => x"93",
          8388 => x"93",
          8389 => x"fc",
          8390 => x"af",
          8391 => x"fc",
          8392 => x"3d",
          8393 => x"51",
          8394 => x"3f",
          8395 => x"08",
          8396 => x"84",
          8397 => x"fe",
          8398 => x"81",
          8399 => x"84",
          8400 => x"51",
          8401 => x"80",
          8402 => x"3d",
          8403 => x"51",
          8404 => x"3f",
          8405 => x"08",
          8406 => x"84",
          8407 => x"fe",
          8408 => x"82",
          8409 => x"b5",
          8410 => x"05",
          8411 => x"cd",
          8412 => x"93",
          8413 => x"3d",
          8414 => x"52",
          8415 => x"a8",
          8416 => x"80",
          8417 => x"cc",
          8418 => x"80",
          8419 => x"84",
          8420 => x"06",
          8421 => x"79",
          8422 => x"f2",
          8423 => x"93",
          8424 => x"2e",
          8425 => x"82",
          8426 => x"51",
          8427 => x"fa",
          8428 => x"3d",
          8429 => x"53",
          8430 => x"51",
          8431 => x"3f",
          8432 => x"08",
          8433 => x"de",
          8434 => x"fe",
          8435 => x"ff",
          8436 => x"fe",
          8437 => x"82",
          8438 => x"80",
          8439 => x"38",
          8440 => x"f8",
          8441 => x"84",
          8442 => x"ea",
          8443 => x"93",
          8444 => x"38",
          8445 => x"08",
          8446 => x"b0",
          8447 => x"cb",
          8448 => x"5c",
          8449 => x"27",
          8450 => x"61",
          8451 => x"70",
          8452 => x"0c",
          8453 => x"f5",
          8454 => x"39",
          8455 => x"80",
          8456 => x"84",
          8457 => x"e9",
          8458 => x"93",
          8459 => x"2e",
          8460 => x"b4",
          8461 => x"11",
          8462 => x"05",
          8463 => x"e4",
          8464 => x"84",
          8465 => x"f9",
          8466 => x"3d",
          8467 => x"53",
          8468 => x"51",
          8469 => x"3f",
          8470 => x"08",
          8471 => x"c6",
          8472 => x"c0",
          8473 => x"e3",
          8474 => x"79",
          8475 => x"8c",
          8476 => x"79",
          8477 => x"5b",
          8478 => x"61",
          8479 => x"eb",
          8480 => x"ff",
          8481 => x"ff",
          8482 => x"fe",
          8483 => x"82",
          8484 => x"80",
          8485 => x"38",
          8486 => x"fc",
          8487 => x"84",
          8488 => x"e8",
          8489 => x"93",
          8490 => x"2e",
          8491 => x"b4",
          8492 => x"11",
          8493 => x"05",
          8494 => x"e8",
          8495 => x"84",
          8496 => x"f8",
          8497 => x"8a",
          8498 => x"e0",
          8499 => x"5a",
          8500 => x"a8",
          8501 => x"33",
          8502 => x"5a",
          8503 => x"2e",
          8504 => x"55",
          8505 => x"33",
          8506 => x"82",
          8507 => x"fe",
          8508 => x"81",
          8509 => x"05",
          8510 => x"39",
          8511 => x"51",
          8512 => x"b4",
          8513 => x"11",
          8514 => x"05",
          8515 => x"94",
          8516 => x"84",
          8517 => x"38",
          8518 => x"33",
          8519 => x"2e",
          8520 => x"8e",
          8521 => x"80",
          8522 => x"8e",
          8523 => x"78",
          8524 => x"38",
          8525 => x"08",
          8526 => x"82",
          8527 => x"59",
          8528 => x"88",
          8529 => x"90",
          8530 => x"39",
          8531 => x"33",
          8532 => x"2e",
          8533 => x"8e",
          8534 => x"9a",
          8535 => x"c6",
          8536 => x"80",
          8537 => x"82",
          8538 => x"44",
          8539 => x"8e",
          8540 => x"80",
          8541 => x"3d",
          8542 => x"53",
          8543 => x"51",
          8544 => x"3f",
          8545 => x"08",
          8546 => x"82",
          8547 => x"59",
          8548 => x"89",
          8549 => x"84",
          8550 => x"cc",
          8551 => x"c9",
          8552 => x"80",
          8553 => x"82",
          8554 => x"43",
          8555 => x"8e",
          8556 => x"78",
          8557 => x"38",
          8558 => x"08",
          8559 => x"82",
          8560 => x"59",
          8561 => x"88",
          8562 => x"9c",
          8563 => x"39",
          8564 => x"33",
          8565 => x"2e",
          8566 => x"8e",
          8567 => x"88",
          8568 => x"b0",
          8569 => x"43",
          8570 => x"f8",
          8571 => x"84",
          8572 => x"e6",
          8573 => x"93",
          8574 => x"2e",
          8575 => x"62",
          8576 => x"88",
          8577 => x"81",
          8578 => x"32",
          8579 => x"72",
          8580 => x"70",
          8581 => x"51",
          8582 => x"80",
          8583 => x"7a",
          8584 => x"38",
          8585 => x"8a",
          8586 => x"de",
          8587 => x"55",
          8588 => x"53",
          8589 => x"51",
          8590 => x"82",
          8591 => x"fe",
          8592 => x"f5",
          8593 => x"3d",
          8594 => x"53",
          8595 => x"51",
          8596 => x"3f",
          8597 => x"08",
          8598 => x"ca",
          8599 => x"fe",
          8600 => x"ff",
          8601 => x"fe",
          8602 => x"82",
          8603 => x"80",
          8604 => x"63",
          8605 => x"cb",
          8606 => x"34",
          8607 => x"44",
          8608 => x"fc",
          8609 => x"84",
          8610 => x"e5",
          8611 => x"93",
          8612 => x"38",
          8613 => x"63",
          8614 => x"52",
          8615 => x"51",
          8616 => x"3f",
          8617 => x"79",
          8618 => x"dd",
          8619 => x"79",
          8620 => x"ae",
          8621 => x"38",
          8622 => x"a0",
          8623 => x"fe",
          8624 => x"ff",
          8625 => x"fe",
          8626 => x"82",
          8627 => x"80",
          8628 => x"63",
          8629 => x"cb",
          8630 => x"34",
          8631 => x"44",
          8632 => x"82",
          8633 => x"fe",
          8634 => x"ff",
          8635 => x"3d",
          8636 => x"53",
          8637 => x"51",
          8638 => x"3f",
          8639 => x"08",
          8640 => x"a2",
          8641 => x"fe",
          8642 => x"ff",
          8643 => x"fe",
          8644 => x"82",
          8645 => x"80",
          8646 => x"60",
          8647 => x"05",
          8648 => x"82",
          8649 => x"78",
          8650 => x"fe",
          8651 => x"ff",
          8652 => x"fe",
          8653 => x"82",
          8654 => x"df",
          8655 => x"39",
          8656 => x"54",
          8657 => x"a8",
          8658 => x"e3",
          8659 => x"52",
          8660 => x"e2",
          8661 => x"45",
          8662 => x"78",
          8663 => x"c6",
          8664 => x"26",
          8665 => x"82",
          8666 => x"39",
          8667 => x"f0",
          8668 => x"84",
          8669 => x"e5",
          8670 => x"93",
          8671 => x"2e",
          8672 => x"59",
          8673 => x"22",
          8674 => x"05",
          8675 => x"41",
          8676 => x"82",
          8677 => x"fe",
          8678 => x"ff",
          8679 => x"3d",
          8680 => x"53",
          8681 => x"51",
          8682 => x"3f",
          8683 => x"08",
          8684 => x"f2",
          8685 => x"fe",
          8686 => x"ff",
          8687 => x"fe",
          8688 => x"82",
          8689 => x"80",
          8690 => x"60",
          8691 => x"59",
          8692 => x"41",
          8693 => x"f0",
          8694 => x"84",
          8695 => x"e4",
          8696 => x"93",
          8697 => x"38",
          8698 => x"60",
          8699 => x"52",
          8700 => x"51",
          8701 => x"3f",
          8702 => x"79",
          8703 => x"89",
          8704 => x"79",
          8705 => x"ae",
          8706 => x"38",
          8707 => x"9c",
          8708 => x"fe",
          8709 => x"ff",
          8710 => x"fe",
          8711 => x"82",
          8712 => x"80",
          8713 => x"60",
          8714 => x"59",
          8715 => x"41",
          8716 => x"82",
          8717 => x"fe",
          8718 => x"ff",
          8719 => x"8b",
          8720 => x"da",
          8721 => x"51",
          8722 => x"3f",
          8723 => x"82",
          8724 => x"fe",
          8725 => x"a2",
          8726 => x"aa",
          8727 => x"39",
          8728 => x"51",
          8729 => x"3f",
          8730 => x"0b",
          8731 => x"84",
          8732 => x"81",
          8733 => x"94",
          8734 => x"aa",
          8735 => x"84",
          8736 => x"c7",
          8737 => x"83",
          8738 => x"94",
          8739 => x"80",
          8740 => x"c0",
          8741 => x"f1",
          8742 => x"3d",
          8743 => x"53",
          8744 => x"51",
          8745 => x"3f",
          8746 => x"08",
          8747 => x"f6",
          8748 => x"82",
          8749 => x"fe",
          8750 => x"63",
          8751 => x"b4",
          8752 => x"11",
          8753 => x"05",
          8754 => x"d8",
          8755 => x"84",
          8756 => x"f0",
          8757 => x"52",
          8758 => x"51",
          8759 => x"3f",
          8760 => x"2d",
          8761 => x"08",
          8762 => x"ba",
          8763 => x"84",
          8764 => x"8c",
          8765 => x"de",
          8766 => x"aa",
          8767 => x"ec",
          8768 => x"c7",
          8769 => x"b6",
          8770 => x"39",
          8771 => x"51",
          8772 => x"3f",
          8773 => x"a5",
          8774 => x"89",
          8775 => x"39",
          8776 => x"33",
          8777 => x"2e",
          8778 => x"7d",
          8779 => x"78",
          8780 => x"d3",
          8781 => x"ff",
          8782 => x"fe",
          8783 => x"82",
          8784 => x"5b",
          8785 => x"82",
          8786 => x"7b",
          8787 => x"38",
          8788 => x"8c",
          8789 => x"39",
          8790 => x"b0",
          8791 => x"39",
          8792 => x"56",
          8793 => x"8d",
          8794 => x"53",
          8795 => x"52",
          8796 => x"b0",
          8797 => x"dd",
          8798 => x"39",
          8799 => x"52",
          8800 => x"b0",
          8801 => x"dd",
          8802 => x"39",
          8803 => x"8d",
          8804 => x"53",
          8805 => x"52",
          8806 => x"b0",
          8807 => x"dd",
          8808 => x"39",
          8809 => x"53",
          8810 => x"52",
          8811 => x"b0",
          8812 => x"dd",
          8813 => x"8e",
          8814 => x"93",
          8815 => x"56",
          8816 => x"54",
          8817 => x"53",
          8818 => x"52",
          8819 => x"b0",
          8820 => x"c8",
          8821 => x"84",
          8822 => x"84",
          8823 => x"30",
          8824 => x"80",
          8825 => x"5b",
          8826 => x"7b",
          8827 => x"38",
          8828 => x"7a",
          8829 => x"80",
          8830 => x"81",
          8831 => x"ff",
          8832 => x"7b",
          8833 => x"7d",
          8834 => x"81",
          8835 => x"78",
          8836 => x"ff",
          8837 => x"06",
          8838 => x"82",
          8839 => x"fe",
          8840 => x"ee",
          8841 => x"3d",
          8842 => x"82",
          8843 => x"87",
          8844 => x"70",
          8845 => x"87",
          8846 => x"72",
          8847 => x"9e",
          8848 => x"84",
          8849 => x"75",
          8850 => x"87",
          8851 => x"73",
          8852 => x"8a",
          8853 => x"93",
          8854 => x"75",
          8855 => x"94",
          8856 => x"54",
          8857 => x"80",
          8858 => x"fe",
          8859 => x"82",
          8860 => x"90",
          8861 => x"55",
          8862 => x"80",
          8863 => x"fe",
          8864 => x"72",
          8865 => x"08",
          8866 => x"8c",
          8867 => x"87",
          8868 => x"0c",
          8869 => x"0b",
          8870 => x"94",
          8871 => x"0b",
          8872 => x"0c",
          8873 => x"82",
          8874 => x"fe",
          8875 => x"fe",
          8876 => x"82",
          8877 => x"fe",
          8878 => x"82",
          8879 => x"fe",
          8880 => x"81",
          8881 => x"fe",
          8882 => x"81",
          8883 => x"3f",
          8884 => x"80",
          8885 => x"00",
          8886 => x"00",
          8887 => x"00",
          8888 => x"00",
          8889 => x"00",
          8890 => x"00",
          8891 => x"00",
          8892 => x"00",
          8893 => x"00",
          8894 => x"00",
          8895 => x"00",
          8896 => x"00",
          8897 => x"00",
          8898 => x"00",
          8899 => x"00",
          8900 => x"00",
          8901 => x"00",
          8902 => x"00",
          8903 => x"00",
          8904 => x"00",
          8905 => x"00",
          8906 => x"00",
          8907 => x"00",
          8908 => x"00",
          8909 => x"00",
          8910 => x"00",
          8911 => x"00",
          8912 => x"00",
          8913 => x"00",
          8914 => x"00",
          8915 => x"00",
          8916 => x"00",
          8917 => x"00",
          8918 => x"00",
          8919 => x"00",
          8920 => x"00",
          8921 => x"00",
          8922 => x"25",
          8923 => x"64",
          8924 => x"20",
          8925 => x"25",
          8926 => x"64",
          8927 => x"25",
          8928 => x"53",
          8929 => x"43",
          8930 => x"69",
          8931 => x"61",
          8932 => x"6e",
          8933 => x"20",
          8934 => x"6f",
          8935 => x"6f",
          8936 => x"6f",
          8937 => x"67",
          8938 => x"3a",
          8939 => x"76",
          8940 => x"73",
          8941 => x"70",
          8942 => x"65",
          8943 => x"64",
          8944 => x"20",
          8945 => x"57",
          8946 => x"44",
          8947 => x"20",
          8948 => x"30",
          8949 => x"25",
          8950 => x"29",
          8951 => x"20",
          8952 => x"53",
          8953 => x"4d",
          8954 => x"20",
          8955 => x"30",
          8956 => x"25",
          8957 => x"29",
          8958 => x"20",
          8959 => x"49",
          8960 => x"20",
          8961 => x"4d",
          8962 => x"30",
          8963 => x"25",
          8964 => x"29",
          8965 => x"20",
          8966 => x"42",
          8967 => x"20",
          8968 => x"20",
          8969 => x"30",
          8970 => x"25",
          8971 => x"29",
          8972 => x"20",
          8973 => x"52",
          8974 => x"20",
          8975 => x"20",
          8976 => x"30",
          8977 => x"25",
          8978 => x"29",
          8979 => x"20",
          8980 => x"53",
          8981 => x"41",
          8982 => x"20",
          8983 => x"65",
          8984 => x"65",
          8985 => x"25",
          8986 => x"29",
          8987 => x"20",
          8988 => x"54",
          8989 => x"52",
          8990 => x"20",
          8991 => x"69",
          8992 => x"73",
          8993 => x"25",
          8994 => x"29",
          8995 => x"20",
          8996 => x"49",
          8997 => x"20",
          8998 => x"4c",
          8999 => x"68",
          9000 => x"65",
          9001 => x"25",
          9002 => x"29",
          9003 => x"20",
          9004 => x"57",
          9005 => x"42",
          9006 => x"20",
          9007 => x"0a",
          9008 => x"20",
          9009 => x"57",
          9010 => x"32",
          9011 => x"20",
          9012 => x"49",
          9013 => x"4c",
          9014 => x"20",
          9015 => x"50",
          9016 => x"00",
          9017 => x"20",
          9018 => x"53",
          9019 => x"00",
          9020 => x"41",
          9021 => x"65",
          9022 => x"73",
          9023 => x"20",
          9024 => x"43",
          9025 => x"52",
          9026 => x"74",
          9027 => x"63",
          9028 => x"20",
          9029 => x"72",
          9030 => x"20",
          9031 => x"30",
          9032 => x"00",
          9033 => x"20",
          9034 => x"43",
          9035 => x"4d",
          9036 => x"72",
          9037 => x"74",
          9038 => x"20",
          9039 => x"72",
          9040 => x"20",
          9041 => x"30",
          9042 => x"00",
          9043 => x"20",
          9044 => x"53",
          9045 => x"6b",
          9046 => x"61",
          9047 => x"41",
          9048 => x"65",
          9049 => x"20",
          9050 => x"20",
          9051 => x"30",
          9052 => x"00",
          9053 => x"4d",
          9054 => x"3a",
          9055 => x"20",
          9056 => x"5a",
          9057 => x"49",
          9058 => x"20",
          9059 => x"20",
          9060 => x"20",
          9061 => x"20",
          9062 => x"20",
          9063 => x"30",
          9064 => x"00",
          9065 => x"20",
          9066 => x"53",
          9067 => x"65",
          9068 => x"6c",
          9069 => x"20",
          9070 => x"71",
          9071 => x"20",
          9072 => x"20",
          9073 => x"64",
          9074 => x"34",
          9075 => x"7a",
          9076 => x"20",
          9077 => x"53",
          9078 => x"4d",
          9079 => x"6f",
          9080 => x"46",
          9081 => x"20",
          9082 => x"20",
          9083 => x"20",
          9084 => x"64",
          9085 => x"34",
          9086 => x"7a",
          9087 => x"20",
          9088 => x"57",
          9089 => x"62",
          9090 => x"20",
          9091 => x"41",
          9092 => x"6c",
          9093 => x"20",
          9094 => x"71",
          9095 => x"64",
          9096 => x"34",
          9097 => x"7a",
          9098 => x"53",
          9099 => x"6c",
          9100 => x"4d",
          9101 => x"75",
          9102 => x"46",
          9103 => x"00",
          9104 => x"45",
          9105 => x"45",
          9106 => x"69",
          9107 => x"55",
          9108 => x"6f",
          9109 => x"68",
          9110 => x"6f",
          9111 => x"74",
          9112 => x"68",
          9113 => x"6f",
          9114 => x"68",
          9115 => x"00",
          9116 => x"21",
          9117 => x"25",
          9118 => x"20",
          9119 => x"0a",
          9120 => x"46",
          9121 => x"65",
          9122 => x"6f",
          9123 => x"73",
          9124 => x"74",
          9125 => x"68",
          9126 => x"6f",
          9127 => x"66",
          9128 => x"20",
          9129 => x"45",
          9130 => x"0a",
          9131 => x"43",
          9132 => x"6f",
          9133 => x"70",
          9134 => x"63",
          9135 => x"74",
          9136 => x"69",
          9137 => x"72",
          9138 => x"69",
          9139 => x"20",
          9140 => x"61",
          9141 => x"6e",
          9142 => x"00",
          9143 => x"00",
          9144 => x"01",
          9145 => x"00",
          9146 => x"00",
          9147 => x"01",
          9148 => x"00",
          9149 => x"00",
          9150 => x"04",
          9151 => x"00",
          9152 => x"00",
          9153 => x"04",
          9154 => x"00",
          9155 => x"00",
          9156 => x"04",
          9157 => x"00",
          9158 => x"00",
          9159 => x"04",
          9160 => x"00",
          9161 => x"00",
          9162 => x"04",
          9163 => x"00",
          9164 => x"00",
          9165 => x"03",
          9166 => x"00",
          9167 => x"00",
          9168 => x"03",
          9169 => x"00",
          9170 => x"00",
          9171 => x"03",
          9172 => x"00",
          9173 => x"00",
          9174 => x"03",
          9175 => x"00",
          9176 => x"1b",
          9177 => x"1b",
          9178 => x"1b",
          9179 => x"1b",
          9180 => x"1b",
          9181 => x"1b",
          9182 => x"1b",
          9183 => x"1b",
          9184 => x"1b",
          9185 => x"0d",
          9186 => x"08",
          9187 => x"53",
          9188 => x"22",
          9189 => x"3a",
          9190 => x"3e",
          9191 => x"7c",
          9192 => x"46",
          9193 => x"46",
          9194 => x"32",
          9195 => x"eb",
          9196 => x"53",
          9197 => x"35",
          9198 => x"4e",
          9199 => x"41",
          9200 => x"20",
          9201 => x"41",
          9202 => x"20",
          9203 => x"4e",
          9204 => x"41",
          9205 => x"20",
          9206 => x"41",
          9207 => x"20",
          9208 => x"00",
          9209 => x"00",
          9210 => x"00",
          9211 => x"00",
          9212 => x"80",
          9213 => x"8e",
          9214 => x"45",
          9215 => x"49",
          9216 => x"90",
          9217 => x"99",
          9218 => x"59",
          9219 => x"9c",
          9220 => x"41",
          9221 => x"a5",
          9222 => x"a8",
          9223 => x"ac",
          9224 => x"b0",
          9225 => x"b4",
          9226 => x"b8",
          9227 => x"bc",
          9228 => x"c0",
          9229 => x"c4",
          9230 => x"c8",
          9231 => x"cc",
          9232 => x"d0",
          9233 => x"d4",
          9234 => x"d8",
          9235 => x"dc",
          9236 => x"e0",
          9237 => x"e4",
          9238 => x"e8",
          9239 => x"ec",
          9240 => x"f0",
          9241 => x"f4",
          9242 => x"f8",
          9243 => x"fc",
          9244 => x"2b",
          9245 => x"3d",
          9246 => x"5c",
          9247 => x"3c",
          9248 => x"7f",
          9249 => x"00",
          9250 => x"00",
          9251 => x"01",
          9252 => x"00",
          9253 => x"00",
          9254 => x"00",
          9255 => x"00",
          9256 => x"00",
          9257 => x"64",
          9258 => x"74",
          9259 => x"64",
          9260 => x"74",
          9261 => x"66",
          9262 => x"74",
          9263 => x"66",
          9264 => x"64",
          9265 => x"66",
          9266 => x"63",
          9267 => x"6d",
          9268 => x"61",
          9269 => x"6d",
          9270 => x"79",
          9271 => x"6d",
          9272 => x"66",
          9273 => x"6d",
          9274 => x"70",
          9275 => x"6d",
          9276 => x"6d",
          9277 => x"6d",
          9278 => x"68",
          9279 => x"68",
          9280 => x"68",
          9281 => x"68",
          9282 => x"63",
          9283 => x"00",
          9284 => x"6a",
          9285 => x"72",
          9286 => x"61",
          9287 => x"72",
          9288 => x"74",
          9289 => x"69",
          9290 => x"00",
          9291 => x"74",
          9292 => x"00",
          9293 => x"74",
          9294 => x"69",
          9295 => x"6d",
          9296 => x"69",
          9297 => x"6b",
          9298 => x"00",
          9299 => x"44",
          9300 => x"20",
          9301 => x"6f",
          9302 => x"49",
          9303 => x"72",
          9304 => x"20",
          9305 => x"6f",
          9306 => x"00",
          9307 => x"44",
          9308 => x"20",
          9309 => x"20",
          9310 => x"64",
          9311 => x"00",
          9312 => x"4e",
          9313 => x"69",
          9314 => x"66",
          9315 => x"64",
          9316 => x"4e",
          9317 => x"61",
          9318 => x"66",
          9319 => x"64",
          9320 => x"49",
          9321 => x"6c",
          9322 => x"66",
          9323 => x"6e",
          9324 => x"2e",
          9325 => x"41",
          9326 => x"73",
          9327 => x"65",
          9328 => x"64",
          9329 => x"46",
          9330 => x"20",
          9331 => x"65",
          9332 => x"20",
          9333 => x"73",
          9334 => x"0a",
          9335 => x"46",
          9336 => x"20",
          9337 => x"64",
          9338 => x"69",
          9339 => x"6c",
          9340 => x"0a",
          9341 => x"53",
          9342 => x"73",
          9343 => x"69",
          9344 => x"70",
          9345 => x"65",
          9346 => x"64",
          9347 => x"44",
          9348 => x"65",
          9349 => x"6d",
          9350 => x"20",
          9351 => x"69",
          9352 => x"6c",
          9353 => x"0a",
          9354 => x"44",
          9355 => x"20",
          9356 => x"20",
          9357 => x"62",
          9358 => x"2e",
          9359 => x"4e",
          9360 => x"6f",
          9361 => x"74",
          9362 => x"65",
          9363 => x"6c",
          9364 => x"73",
          9365 => x"20",
          9366 => x"6e",
          9367 => x"6e",
          9368 => x"73",
          9369 => x"00",
          9370 => x"46",
          9371 => x"61",
          9372 => x"62",
          9373 => x"65",
          9374 => x"00",
          9375 => x"54",
          9376 => x"6f",
          9377 => x"20",
          9378 => x"72",
          9379 => x"6f",
          9380 => x"61",
          9381 => x"6c",
          9382 => x"2e",
          9383 => x"46",
          9384 => x"20",
          9385 => x"6c",
          9386 => x"65",
          9387 => x"00",
          9388 => x"49",
          9389 => x"66",
          9390 => x"69",
          9391 => x"20",
          9392 => x"6f",
          9393 => x"0a",
          9394 => x"54",
          9395 => x"6d",
          9396 => x"20",
          9397 => x"6e",
          9398 => x"6c",
          9399 => x"0a",
          9400 => x"50",
          9401 => x"6d",
          9402 => x"72",
          9403 => x"6e",
          9404 => x"72",
          9405 => x"2e",
          9406 => x"53",
          9407 => x"65",
          9408 => x"0a",
          9409 => x"55",
          9410 => x"6f",
          9411 => x"65",
          9412 => x"72",
          9413 => x"0a",
          9414 => x"20",
          9415 => x"65",
          9416 => x"73",
          9417 => x"20",
          9418 => x"20",
          9419 => x"65",
          9420 => x"65",
          9421 => x"00",
          9422 => x"72",
          9423 => x"00",
          9424 => x"25",
          9425 => x"00",
          9426 => x"3a",
          9427 => x"25",
          9428 => x"00",
          9429 => x"20",
          9430 => x"20",
          9431 => x"00",
          9432 => x"25",
          9433 => x"00",
          9434 => x"20",
          9435 => x"20",
          9436 => x"7c",
          9437 => x"5a",
          9438 => x"41",
          9439 => x"0a",
          9440 => x"25",
          9441 => x"00",
          9442 => x"32",
          9443 => x"34",
          9444 => x"32",
          9445 => x"76",
          9446 => x"31",
          9447 => x"20",
          9448 => x"2c",
          9449 => x"76",
          9450 => x"32",
          9451 => x"25",
          9452 => x"73",
          9453 => x"0a",
          9454 => x"5a",
          9455 => x"41",
          9456 => x"74",
          9457 => x"75",
          9458 => x"48",
          9459 => x"6c",
          9460 => x"00",
          9461 => x"54",
          9462 => x"72",
          9463 => x"74",
          9464 => x"75",
          9465 => x"00",
          9466 => x"50",
          9467 => x"69",
          9468 => x"72",
          9469 => x"74",
          9470 => x"49",
          9471 => x"4c",
          9472 => x"20",
          9473 => x"65",
          9474 => x"70",
          9475 => x"49",
          9476 => x"4c",
          9477 => x"20",
          9478 => x"65",
          9479 => x"70",
          9480 => x"55",
          9481 => x"30",
          9482 => x"20",
          9483 => x"65",
          9484 => x"70",
          9485 => x"55",
          9486 => x"30",
          9487 => x"20",
          9488 => x"65",
          9489 => x"70",
          9490 => x"55",
          9491 => x"31",
          9492 => x"20",
          9493 => x"65",
          9494 => x"70",
          9495 => x"55",
          9496 => x"31",
          9497 => x"20",
          9498 => x"65",
          9499 => x"70",
          9500 => x"53",
          9501 => x"69",
          9502 => x"75",
          9503 => x"69",
          9504 => x"2e",
          9505 => x"00",
          9506 => x"45",
          9507 => x"6c",
          9508 => x"20",
          9509 => x"65",
          9510 => x"2e",
          9511 => x"61",
          9512 => x"65",
          9513 => x"2e",
          9514 => x"00",
          9515 => x"30",
          9516 => x"46",
          9517 => x"65",
          9518 => x"6f",
          9519 => x"69",
          9520 => x"6c",
          9521 => x"20",
          9522 => x"63",
          9523 => x"20",
          9524 => x"70",
          9525 => x"73",
          9526 => x"6e",
          9527 => x"6d",
          9528 => x"61",
          9529 => x"2e",
          9530 => x"2a",
          9531 => x"42",
          9532 => x"64",
          9533 => x"20",
          9534 => x"0a",
          9535 => x"49",
          9536 => x"69",
          9537 => x"73",
          9538 => x"0a",
          9539 => x"46",
          9540 => x"65",
          9541 => x"6f",
          9542 => x"69",
          9543 => x"6c",
          9544 => x"2e",
          9545 => x"72",
          9546 => x"64",
          9547 => x"25",
          9548 => x"43",
          9549 => x"72",
          9550 => x"2e",
          9551 => x"00",
          9552 => x"43",
          9553 => x"69",
          9554 => x"2e",
          9555 => x"43",
          9556 => x"61",
          9557 => x"67",
          9558 => x"00",
          9559 => x"25",
          9560 => x"78",
          9561 => x"38",
          9562 => x"3e",
          9563 => x"6c",
          9564 => x"30",
          9565 => x"0a",
          9566 => x"44",
          9567 => x"20",
          9568 => x"6f",
          9569 => x"00",
          9570 => x"0a",
          9571 => x"70",
          9572 => x"65",
          9573 => x"25",
          9574 => x"20",
          9575 => x"58",
          9576 => x"3f",
          9577 => x"00",
          9578 => x"25",
          9579 => x"20",
          9580 => x"58",
          9581 => x"25",
          9582 => x"20",
          9583 => x"58",
          9584 => x"44",
          9585 => x"62",
          9586 => x"67",
          9587 => x"74",
          9588 => x"75",
          9589 => x"0a",
          9590 => x"45",
          9591 => x"6c",
          9592 => x"20",
          9593 => x"65",
          9594 => x"70",
          9595 => x"00",
          9596 => x"44",
          9597 => x"62",
          9598 => x"20",
          9599 => x"74",
          9600 => x"66",
          9601 => x"45",
          9602 => x"6c",
          9603 => x"20",
          9604 => x"74",
          9605 => x"66",
          9606 => x"45",
          9607 => x"75",
          9608 => x"67",
          9609 => x"64",
          9610 => x"20",
          9611 => x"78",
          9612 => x"2e",
          9613 => x"43",
          9614 => x"69",
          9615 => x"63",
          9616 => x"20",
          9617 => x"30",
          9618 => x"2e",
          9619 => x"00",
          9620 => x"43",
          9621 => x"20",
          9622 => x"75",
          9623 => x"64",
          9624 => x"64",
          9625 => x"25",
          9626 => x"0a",
          9627 => x"52",
          9628 => x"61",
          9629 => x"6e",
          9630 => x"70",
          9631 => x"63",
          9632 => x"6f",
          9633 => x"2e",
          9634 => x"43",
          9635 => x"20",
          9636 => x"6f",
          9637 => x"6e",
          9638 => x"2e",
          9639 => x"5a",
          9640 => x"62",
          9641 => x"25",
          9642 => x"25",
          9643 => x"73",
          9644 => x"00",
          9645 => x"25",
          9646 => x"25",
          9647 => x"73",
          9648 => x"25",
          9649 => x"25",
          9650 => x"42",
          9651 => x"63",
          9652 => x"61",
          9653 => x"0a",
          9654 => x"52",
          9655 => x"69",
          9656 => x"2e",
          9657 => x"45",
          9658 => x"6c",
          9659 => x"20",
          9660 => x"65",
          9661 => x"70",
          9662 => x"2e",
          9663 => x"00",
          9664 => x"00",
          9665 => x"00",
          9666 => x"00",
          9667 => x"00",
          9668 => x"00",
          9669 => x"00",
          9670 => x"00",
          9671 => x"00",
          9672 => x"01",
          9673 => x"01",
          9674 => x"00",
          9675 => x"00",
          9676 => x"00",
          9677 => x"00",
          9678 => x"05",
          9679 => x"05",
          9680 => x"05",
          9681 => x"00",
          9682 => x"01",
          9683 => x"01",
          9684 => x"01",
          9685 => x"01",
          9686 => x"00",
          9687 => x"00",
          9688 => x"00",
          9689 => x"00",
          9690 => x"00",
          9691 => x"00",
          9692 => x"00",
          9693 => x"00",
          9694 => x"00",
          9695 => x"00",
          9696 => x"00",
          9697 => x"00",
          9698 => x"00",
          9699 => x"00",
          9700 => x"00",
          9701 => x"00",
          9702 => x"00",
          9703 => x"00",
          9704 => x"00",
          9705 => x"00",
          9706 => x"00",
          9707 => x"00",
          9708 => x"00",
          9709 => x"00",
          9710 => x"00",
          9711 => x"00",
          9712 => x"00",
          9713 => x"00",
          9714 => x"00",
          9715 => x"00",
          9716 => x"00",
          9717 => x"00",
          9718 => x"01",
          9719 => x"00",
          9720 => x"01",
          9721 => x"00",
          9722 => x"02",
          9723 => x"01",
          9724 => x"00",
          9725 => x"00",
          9726 => x"01",
          9727 => x"00",
          9728 => x"00",
          9729 => x"00",
          9730 => x"01",
          9731 => x"00",
          9732 => x"00",
          9733 => x"00",
          9734 => x"01",
          9735 => x"00",
          9736 => x"00",
          9737 => x"00",
          9738 => x"01",
          9739 => x"00",
          9740 => x"00",
          9741 => x"00",
          9742 => x"01",
          9743 => x"00",
          9744 => x"00",
          9745 => x"00",
          9746 => x"01",
          9747 => x"00",
          9748 => x"00",
          9749 => x"00",
          9750 => x"01",
          9751 => x"00",
          9752 => x"00",
          9753 => x"00",
          9754 => x"01",
          9755 => x"00",
          9756 => x"00",
          9757 => x"00",
          9758 => x"01",
          9759 => x"00",
          9760 => x"00",
          9761 => x"00",
          9762 => x"01",
          9763 => x"00",
          9764 => x"00",
          9765 => x"00",
          9766 => x"01",
          9767 => x"00",
          9768 => x"00",
          9769 => x"00",
          9770 => x"01",
          9771 => x"00",
          9772 => x"00",
          9773 => x"00",
          9774 => x"01",
          9775 => x"00",
          9776 => x"00",
          9777 => x"00",
          9778 => x"01",
          9779 => x"00",
          9780 => x"00",
          9781 => x"00",
          9782 => x"01",
          9783 => x"00",
          9784 => x"00",
          9785 => x"00",
          9786 => x"01",
          9787 => x"00",
          9788 => x"00",
          9789 => x"00",
          9790 => x"01",
          9791 => x"00",
          9792 => x"00",
          9793 => x"00",
          9794 => x"01",
          9795 => x"00",
          9796 => x"00",
          9797 => x"00",
          9798 => x"01",
          9799 => x"00",
          9800 => x"00",
          9801 => x"00",
          9802 => x"01",
          9803 => x"00",
          9804 => x"00",
          9805 => x"00",
          9806 => x"01",
          9807 => x"00",
          9808 => x"00",
          9809 => x"00",
          9810 => x"01",
          9811 => x"00",
          9812 => x"00",
          9813 => x"00",
          9814 => x"01",
          9815 => x"00",
          9816 => x"00",
          9817 => x"00",
          9818 => x"01",
          9819 => x"00",
          9820 => x"00",
          9821 => x"00",
          9822 => x"01",
          9823 => x"00",
          9824 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);

    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
