-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Philip Smart 02/2019 for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity BootROM is
port (
        clk                  : in  std_logic;
        areset               : in  std_logic := '0';
        memAWriteEnable      : in  std_logic;
        memAAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memBWriteEnable      : in  std_logic;
        memBAddr             : in  std_logic_vector(ADDR_32BIT_BRAM_RANGE);
        memBWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE);
        memBRead             : out std_logic_vector(WORD_32BIT_RANGE)
);
end BootROM;

architecture arch of BootROM is

type ram_type is array(natural range 0 to (2**(SOC_MAX_ADDR_BRAM_BIT-2))-1) of std_logic_vector(WORD_32BIT_RANGE);

shared variable ram : ram_type :=
(
             0 => x"0b0b0b88",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"88088c08",
             9 => x"90080b0b",
            10 => x"0b888008",
            11 => x"2d900c8c",
            12 => x"0c880c04",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a50400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"09810572",
            51 => x"0a100a72",
            52 => x"0a100a31",
            53 => x"050a8106",
            54 => x"51515351",
            55 => x"04000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c4040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a7",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"04067383",
           106 => x"06098105",
           107 => x"8205832b",
           108 => x"0b2b0772",
           109 => x"fc060c51",
           110 => x"51040000",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9f",
           162 => x"d0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88ac0400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"88088c08",
           169 => x"90087575",
           170 => x"0b0b0b89",
           171 => x"cf2d5050",
           172 => x"88085690",
           173 => x"0c8c0c88",
           174 => x"0c510400",
           175 => x"00000000",
           176 => x"88088c08",
           177 => x"90087575",
           178 => x"0b0b0b8b",
           179 => x"812d5050",
           180 => x"88085690",
           181 => x"0c8c0c88",
           182 => x"0c510400",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"04000000",
           209 => x"00000000",
           210 => x"00000000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"04000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"00000404",
           257 => x"04000000",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10101053",
           266 => x"51040000",
           267 => x"7381ff06",
           268 => x"73830609",
           269 => x"81058305",
           270 => x"1010102b",
           271 => x"0772fc06",
           272 => x"0c515104",
           273 => x"72728072",
           274 => x"8106ff05",
           275 => x"09720605",
           276 => x"71105272",
           277 => x"0a100a53",
           278 => x"72ed3851",
           279 => x"51535104",
           280 => x"9ff470a0",
           281 => x"a4278e38",
           282 => x"80717084",
           283 => x"05530c0b",
           284 => x"0b0b88e2",
           285 => x"0488fe51",
           286 => x"9e9d0400",
           287 => x"80040088",
           288 => x"fe040000",
           289 => x"00940802",
           290 => x"940cfd3d",
           291 => x"0d805394",
           292 => x"088c0508",
           293 => x"52940888",
           294 => x"05085182",
           295 => x"de3f8808",
           296 => x"70880c54",
           297 => x"853d0d94",
           298 => x"0c049408",
           299 => x"02940cfd",
           300 => x"3d0d8153",
           301 => x"94088c05",
           302 => x"08529408",
           303 => x"88050851",
           304 => x"82b93f88",
           305 => x"0870880c",
           306 => x"54853d0d",
           307 => x"940c0494",
           308 => x"0802940c",
           309 => x"f93d0d80",
           310 => x"0b9408fc",
           311 => x"050c9408",
           312 => x"88050880",
           313 => x"25ab3894",
           314 => x"08880508",
           315 => x"30940888",
           316 => x"050c800b",
           317 => x"9408f405",
           318 => x"0c9408fc",
           319 => x"05088838",
           320 => x"810b9408",
           321 => x"f4050c94",
           322 => x"08f40508",
           323 => x"9408fc05",
           324 => x"0c94088c",
           325 => x"05088025",
           326 => x"ab389408",
           327 => x"8c050830",
           328 => x"94088c05",
           329 => x"0c800b94",
           330 => x"08f0050c",
           331 => x"9408fc05",
           332 => x"08883881",
           333 => x"0b9408f0",
           334 => x"050c9408",
           335 => x"f0050894",
           336 => x"08fc050c",
           337 => x"80539408",
           338 => x"8c050852",
           339 => x"94088805",
           340 => x"085181a7",
           341 => x"3f880870",
           342 => x"9408f805",
           343 => x"0c549408",
           344 => x"fc050880",
           345 => x"2e8c3894",
           346 => x"08f80508",
           347 => x"309408f8",
           348 => x"050c9408",
           349 => x"f8050870",
           350 => x"880c5489",
           351 => x"3d0d940c",
           352 => x"04940802",
           353 => x"940cfb3d",
           354 => x"0d800b94",
           355 => x"08fc050c",
           356 => x"94088805",
           357 => x"08802593",
           358 => x"38940888",
           359 => x"05083094",
           360 => x"0888050c",
           361 => x"810b9408",
           362 => x"fc050c94",
           363 => x"088c0508",
           364 => x"80258c38",
           365 => x"94088c05",
           366 => x"08309408",
           367 => x"8c050c81",
           368 => x"5394088c",
           369 => x"05085294",
           370 => x"08880508",
           371 => x"51ad3f88",
           372 => x"08709408",
           373 => x"f8050c54",
           374 => x"9408fc05",
           375 => x"08802e8c",
           376 => x"389408f8",
           377 => x"05083094",
           378 => x"08f8050c",
           379 => x"9408f805",
           380 => x"0870880c",
           381 => x"54873d0d",
           382 => x"940c0494",
           383 => x"0802940c",
           384 => x"fd3d0d81",
           385 => x"0b9408fc",
           386 => x"050c800b",
           387 => x"9408f805",
           388 => x"0c94088c",
           389 => x"05089408",
           390 => x"88050827",
           391 => x"ac389408",
           392 => x"fc050880",
           393 => x"2ea33880",
           394 => x"0b94088c",
           395 => x"05082499",
           396 => x"3894088c",
           397 => x"05081094",
           398 => x"088c050c",
           399 => x"9408fc05",
           400 => x"08109408",
           401 => x"fc050cc9",
           402 => x"399408fc",
           403 => x"0508802e",
           404 => x"80c93894",
           405 => x"088c0508",
           406 => x"94088805",
           407 => x"0826a138",
           408 => x"94088805",
           409 => x"0894088c",
           410 => x"05083194",
           411 => x"0888050c",
           412 => x"9408f805",
           413 => x"089408fc",
           414 => x"05080794",
           415 => x"08f8050c",
           416 => x"9408fc05",
           417 => x"08812a94",
           418 => x"08fc050c",
           419 => x"94088c05",
           420 => x"08812a94",
           421 => x"088c050c",
           422 => x"ffaf3994",
           423 => x"08900508",
           424 => x"802e8f38",
           425 => x"94088805",
           426 => x"08709408",
           427 => x"f4050c51",
           428 => x"8d399408",
           429 => x"f8050870",
           430 => x"9408f405",
           431 => x"0c519408",
           432 => x"f4050888",
           433 => x"0c853d0d",
           434 => x"940c04ff",
           435 => x"3d0d8188",
           436 => x"0b87c092",
           437 => x"8c0c810b",
           438 => x"87c0928c",
           439 => x"0c850b87",
           440 => x"c0988c0c",
           441 => x"87c0928c",
           442 => x"08708206",
           443 => x"51517080",
           444 => x"2e8a3887",
           445 => x"c0988c08",
           446 => x"5170e938",
           447 => x"87c0928c",
           448 => x"08fc8080",
           449 => x"06527193",
           450 => x"3887c098",
           451 => x"8c085170",
           452 => x"802e8838",
           453 => x"710b0b0b",
           454 => x"9ff0340b",
           455 => x"0b0b9ff0",
           456 => x"33880c83",
           457 => x"3d0d04fa",
           458 => x"3d0d787b",
           459 => x"7d565856",
           460 => x"800b0b0b",
           461 => x"0b9ff033",
           462 => x"81065255",
           463 => x"82527075",
           464 => x"2e098106",
           465 => x"819e3885",
           466 => x"0b87c098",
           467 => x"8c0c7987",
           468 => x"c092800c",
           469 => x"840b87c0",
           470 => x"928c0c87",
           471 => x"c0928c08",
           472 => x"70852a70",
           473 => x"81065152",
           474 => x"5370802e",
           475 => x"a73887c0",
           476 => x"92840870",
           477 => x"81ff0676",
           478 => x"79275253",
           479 => x"5173802e",
           480 => x"90387080",
           481 => x"2e8b3871",
           482 => x"76708105",
           483 => x"5834ff14",
           484 => x"54811555",
           485 => x"72a20651",
           486 => x"70802e8b",
           487 => x"3887c098",
           488 => x"8c085170",
           489 => x"ffb53887",
           490 => x"c0988c08",
           491 => x"51709538",
           492 => x"810b87c0",
           493 => x"928c0c87",
           494 => x"c0928c08",
           495 => x"70820651",
           496 => x"5170f438",
           497 => x"8073fc80",
           498 => x"80065252",
           499 => x"70722e09",
           500 => x"81068f38",
           501 => x"87c0988c",
           502 => x"08517072",
           503 => x"2e098106",
           504 => x"83388152",
           505 => x"71880c88",
           506 => x"3d0d04fe",
           507 => x"3d0d7481",
           508 => x"11337133",
           509 => x"71882b07",
           510 => x"880c5351",
           511 => x"843d0d04",
           512 => x"fd3d0d75",
           513 => x"83113382",
           514 => x"12337190",
           515 => x"2b71882b",
           516 => x"07811433",
           517 => x"70720788",
           518 => x"2b753371",
           519 => x"07880c52",
           520 => x"53545654",
           521 => x"52853d0d",
           522 => x"04f93d0d",
           523 => x"790b0b0b",
           524 => x"9ff40857",
           525 => x"57817727",
           526 => x"80ed3876",
           527 => x"88170827",
           528 => x"80e53875",
           529 => x"33557482",
           530 => x"2e893874",
           531 => x"832eae38",
           532 => x"80d53974",
           533 => x"54761083",
           534 => x"fe065376",
           535 => x"882a8c17",
           536 => x"08055288",
           537 => x"3d705255",
           538 => x"fdbd3f88",
           539 => x"08b93874",
           540 => x"51fef83f",
           541 => x"880883ff",
           542 => x"ff0655ad",
           543 => x"39845476",
           544 => x"822b83fc",
           545 => x"06537687",
           546 => x"2a8c1708",
           547 => x"0552883d",
           548 => x"705255fd",
           549 => x"923f8808",
           550 => x"8e387451",
           551 => x"fee23f88",
           552 => x"08f00a06",
           553 => x"55833981",
           554 => x"5574880c",
           555 => x"893d0d04",
           556 => x"fb3d0d0b",
           557 => x"0b0b9ff4",
           558 => x"08fe1988",
           559 => x"1208fe05",
           560 => x"55565480",
           561 => x"56747327",
           562 => x"8d388214",
           563 => x"33757129",
           564 => x"94160805",
           565 => x"57537588",
           566 => x"0c873d0d",
           567 => x"04fd3d0d",
           568 => x"7554800b",
           569 => x"0b0b0b9f",
           570 => x"f4087033",
           571 => x"51535371",
           572 => x"832e0981",
           573 => x"068c3894",
           574 => x"1451fdef",
           575 => x"3f880890",
           576 => x"2b539a14",
           577 => x"51fde43f",
           578 => x"880883ff",
           579 => x"ff067307",
           580 => x"880c853d",
           581 => x"0d04fc3d",
           582 => x"0d760b0b",
           583 => x"0b9ff408",
           584 => x"55558075",
           585 => x"23881508",
           586 => x"5372812e",
           587 => x"88388814",
           588 => x"08732685",
           589 => x"388152b0",
           590 => x"39729038",
           591 => x"73335271",
           592 => x"832e0981",
           593 => x"06853890",
           594 => x"14085372",
           595 => x"8c160c72",
           596 => x"802e8b38",
           597 => x"7251fed8",
           598 => x"3f880852",
           599 => x"85399014",
           600 => x"08527190",
           601 => x"160c8052",
           602 => x"71880c86",
           603 => x"3d0d04fa",
           604 => x"3d0d780b",
           605 => x"0b0b9ff4",
           606 => x"08712281",
           607 => x"057083ff",
           608 => x"ff065754",
           609 => x"57557380",
           610 => x"2e883890",
           611 => x"15085372",
           612 => x"86388352",
           613 => x"80dc3973",
           614 => x"8f065271",
           615 => x"80cf3881",
           616 => x"1390160c",
           617 => x"8c150853",
           618 => x"728f3883",
           619 => x"0b841722",
           620 => x"57527376",
           621 => x"27bc38b5",
           622 => x"39821633",
           623 => x"ff057484",
           624 => x"2a065271",
           625 => x"a8387251",
           626 => x"fcdf3f81",
           627 => x"52718808",
           628 => x"27a03883",
           629 => x"52880888",
           630 => x"17082796",
           631 => x"3888088c",
           632 => x"160c8808",
           633 => x"51fdc93f",
           634 => x"88089016",
           635 => x"0c737523",
           636 => x"80527188",
           637 => x"0c883d0d",
           638 => x"04f23d0d",
           639 => x"60626458",
           640 => x"5e5c7533",
           641 => x"5574a02e",
           642 => x"09810688",
           643 => x"38811670",
           644 => x"4456ef39",
           645 => x"62703356",
           646 => x"5674af2e",
           647 => x"09810684",
           648 => x"38811643",
           649 => x"800b881d",
           650 => x"0c627033",
           651 => x"5155749f",
           652 => x"268f387b",
           653 => x"51fddf3f",
           654 => x"88085680",
           655 => x"7d3482d3",
           656 => x"39933d84",
           657 => x"1d087058",
           658 => x"5a5f8a55",
           659 => x"a0767081",
           660 => x"055834ff",
           661 => x"155574ff",
           662 => x"2e098106",
           663 => x"ef388070",
           664 => x"595b887f",
           665 => x"085f5a7a",
           666 => x"811c7081",
           667 => x"ff066013",
           668 => x"703370af",
           669 => x"327030a0",
           670 => x"73277180",
           671 => x"25075151",
           672 => x"525b535d",
           673 => x"57557480",
           674 => x"c73876ae",
           675 => x"2e098106",
           676 => x"83388155",
           677 => x"777a2775",
           678 => x"07557480",
           679 => x"2e9f3879",
           680 => x"88327030",
           681 => x"78ae3270",
           682 => x"30707307",
           683 => x"9f2a5351",
           684 => x"57515675",
           685 => x"9b388858",
           686 => x"8b5affab",
           687 => x"39778119",
           688 => x"7081ff06",
           689 => x"721c535a",
           690 => x"57557675",
           691 => x"34ff9839",
           692 => x"7a1e7f0c",
           693 => x"805576a0",
           694 => x"26833881",
           695 => x"55748b1a",
           696 => x"347b51fc",
           697 => x"b13f8808",
           698 => x"80ef38a0",
           699 => x"547b2270",
           700 => x"852b83e0",
           701 => x"06545590",
           702 => x"1c08527c",
           703 => x"51f8a83f",
           704 => x"88085788",
           705 => x"0880fb38",
           706 => x"7c335574",
           707 => x"802e80ee",
           708 => x"388b1d33",
           709 => x"70832a70",
           710 => x"81065156",
           711 => x"5674b238",
           712 => x"8b7d841e",
           713 => x"08880859",
           714 => x"5b5b58ff",
           715 => x"185877ff",
           716 => x"2e9a3879",
           717 => x"7081055b",
           718 => x"33797081",
           719 => x"055b3371",
           720 => x"71315256",
           721 => x"5675802e",
           722 => x"e2388639",
           723 => x"75802e92",
           724 => x"387b51fc",
           725 => x"9a3fff8e",
           726 => x"39880856",
           727 => x"8808b438",
           728 => x"83397656",
           729 => x"841c088b",
           730 => x"11335155",
           731 => x"74a5388b",
           732 => x"1d337084",
           733 => x"2a708106",
           734 => x"51565674",
           735 => x"89388356",
           736 => x"92398156",
           737 => x"8e397c51",
           738 => x"fad33f88",
           739 => x"08881d0c",
           740 => x"fdaf3975",
           741 => x"880c903d",
           742 => x"0d04f93d",
           743 => x"0d797b59",
           744 => x"57825483",
           745 => x"fe537752",
           746 => x"7651f6fb",
           747 => x"3f835688",
           748 => x"0880e738",
           749 => x"7651f8b3",
           750 => x"3f880883",
           751 => x"ffff0655",
           752 => x"82567482",
           753 => x"d4d52e09",
           754 => x"810680ce",
           755 => x"387554b6",
           756 => x"53775276",
           757 => x"51f6d03f",
           758 => x"88085688",
           759 => x"08943876",
           760 => x"51f8883f",
           761 => x"880883ff",
           762 => x"ff065574",
           763 => x"8182c62e",
           764 => x"a9388254",
           765 => x"80d25377",
           766 => x"527651f6",
           767 => x"aa3f8808",
           768 => x"56880894",
           769 => x"387651f7",
           770 => x"e23f8808",
           771 => x"83ffff06",
           772 => x"55748182",
           773 => x"c62e8338",
           774 => x"81567588",
           775 => x"0c893d0d",
           776 => x"04ed3d0d",
           777 => x"6559800b",
           778 => x"0b0b0b9f",
           779 => x"f40cf59b",
           780 => x"3f880881",
           781 => x"06558256",
           782 => x"7482f238",
           783 => x"7475538d",
           784 => x"3d705357",
           785 => x"5afed33f",
           786 => x"880881ff",
           787 => x"06577681",
           788 => x"2e098106",
           789 => x"b3389054",
           790 => x"83be5374",
           791 => x"527551f5",
           792 => x"c63f8808",
           793 => x"ab388d3d",
           794 => x"33557480",
           795 => x"2eac3895",
           796 => x"3de40551",
           797 => x"f78a3f88",
           798 => x"08880853",
           799 => x"76525afe",
           800 => x"993f8808",
           801 => x"81ff0657",
           802 => x"76832e09",
           803 => x"81068638",
           804 => x"81568299",
           805 => x"3976802e",
           806 => x"86388656",
           807 => x"828f39a4",
           808 => x"548d5379",
           809 => x"527551f4",
           810 => x"fe3f8156",
           811 => x"880881fd",
           812 => x"38953de5",
           813 => x"0551f6b3",
           814 => x"3f880883",
           815 => x"ffff0658",
           816 => x"778c3895",
           817 => x"3df30551",
           818 => x"f6b63f88",
           819 => x"085802af",
           820 => x"05337871",
           821 => x"29028805",
           822 => x"ad057054",
           823 => x"52595bf6",
           824 => x"8a3f8808",
           825 => x"83ffff06",
           826 => x"7a058c1a",
           827 => x"0c8c3d33",
           828 => x"821a3495",
           829 => x"3de00551",
           830 => x"f5f13f88",
           831 => x"08841a23",
           832 => x"953de205",
           833 => x"51f5e43f",
           834 => x"880883ff",
           835 => x"ff065675",
           836 => x"8c38953d",
           837 => x"ef0551f5",
           838 => x"e73f8808",
           839 => x"567a51f5",
           840 => x"ca3f8808",
           841 => x"83ffff06",
           842 => x"76713179",
           843 => x"31841b22",
           844 => x"70842a82",
           845 => x"1d335672",
           846 => x"71315559",
           847 => x"5c5155ee",
           848 => x"c43f8808",
           849 => x"82057088",
           850 => x"1b0c8808",
           851 => x"e08a0556",
           852 => x"567483df",
           853 => x"fe268338",
           854 => x"825783ff",
           855 => x"f6762785",
           856 => x"38835789",
           857 => x"39865676",
           858 => x"802e80c1",
           859 => x"38767934",
           860 => x"76832e09",
           861 => x"81069038",
           862 => x"953dfb05",
           863 => x"51f5813f",
           864 => x"8808901a",
           865 => x"0c88398c",
           866 => x"19081890",
           867 => x"1a0c7983",
           868 => x"ffff068c",
           869 => x"1a081971",
           870 => x"842a0594",
           871 => x"1b0c5580",
           872 => x"0b811a34",
           873 => x"780b0b0b",
           874 => x"9ff40c80",
           875 => x"5675880c",
           876 => x"953d0d04",
           877 => x"ea3d0d0b",
           878 => x"0b0b9ff4",
           879 => x"08558554",
           880 => x"74802e80",
           881 => x"df38800b",
           882 => x"81163498",
           883 => x"3de01145",
           884 => x"6954893d",
           885 => x"705457ec",
           886 => x"0551f89d",
           887 => x"3f880854",
           888 => x"880880c0",
           889 => x"38883d33",
           890 => x"5473802e",
           891 => x"933802a7",
           892 => x"05337084",
           893 => x"2a708106",
           894 => x"51555773",
           895 => x"802e8538",
           896 => x"8354a139",
           897 => x"7551f5d5",
           898 => x"3f8808a0",
           899 => x"160c983d",
           900 => x"dc0551f3",
           901 => x"eb3f8808",
           902 => x"9c160c73",
           903 => x"98160c81",
           904 => x"0b811634",
           905 => x"73880c98",
           906 => x"3d0d04f6",
           907 => x"3d0d7d7f",
           908 => x"7e0b0b0b",
           909 => x"9ff40859",
           910 => x"5b5c5880",
           911 => x"7b0c8557",
           912 => x"75802e81",
           913 => x"d1388116",
           914 => x"33810655",
           915 => x"84577480",
           916 => x"2e81c338",
           917 => x"91397481",
           918 => x"17348639",
           919 => x"800b8117",
           920 => x"34815781",
           921 => x"b1399c16",
           922 => x"08981708",
           923 => x"31557478",
           924 => x"27833874",
           925 => x"5877802e",
           926 => x"819a3898",
           927 => x"16087083",
           928 => x"ff065657",
           929 => x"7480c738",
           930 => x"821633ff",
           931 => x"0577892a",
           932 => x"067081ff",
           933 => x"065b5579",
           934 => x"9e387687",
           935 => x"38a01608",
           936 => x"558b39a4",
           937 => x"160851f3",
           938 => x"803f8808",
           939 => x"55817527",
           940 => x"ffaa3874",
           941 => x"a4170ca4",
           942 => x"160851f3",
           943 => x"f33f8808",
           944 => x"55880880",
           945 => x"2eff8f38",
           946 => x"88081aa8",
           947 => x"170c9816",
           948 => x"0883ff06",
           949 => x"84807131",
           950 => x"51557775",
           951 => x"27833877",
           952 => x"55745498",
           953 => x"160883ff",
           954 => x"0653a816",
           955 => x"08527851",
           956 => x"f0b53f88",
           957 => x"08fee538",
           958 => x"98160815",
           959 => x"98170c77",
           960 => x"75317b08",
           961 => x"167c0c58",
           962 => x"78802efe",
           963 => x"e8387419",
           964 => x"59fee239",
           965 => x"80577688",
           966 => x"0c8c3d0d",
           967 => x"04fb3d0d",
           968 => x"87c0948c",
           969 => x"08548784",
           970 => x"80527351",
           971 => x"ead73f88",
           972 => x"08902b87",
           973 => x"c0948c08",
           974 => x"56548784",
           975 => x"80527451",
           976 => x"eac33f73",
           977 => x"88080787",
           978 => x"c0948c0c",
           979 => x"87c0949c",
           980 => x"08548784",
           981 => x"80527351",
           982 => x"eaab3f88",
           983 => x"08902b87",
           984 => x"c0949c08",
           985 => x"56548784",
           986 => x"80527451",
           987 => x"ea973f73",
           988 => x"88080787",
           989 => x"c0949c0c",
           990 => x"8c80830b",
           991 => x"87c09484",
           992 => x"0c8c8083",
           993 => x"0b87c094",
           994 => x"940c9ff8",
           995 => x"51f9923f",
           996 => x"8808b838",
           997 => x"9fe051fc",
           998 => x"9b3f8808",
           999 => x"ae38a080",
          1000 => x"0b880887",
          1001 => x"c098880c",
          1002 => x"55873dfc",
          1003 => x"05538480",
          1004 => x"527451fc",
          1005 => x"f63f8808",
          1006 => x"8d387554",
          1007 => x"73802e86",
          1008 => x"38731555",
          1009 => x"e439a080",
          1010 => x"54730480",
          1011 => x"54fb3900",
          1012 => x"00ffffff",
          1013 => x"ff00ffff",
          1014 => x"ffff00ff",
          1015 => x"ffffff00",
          1016 => x"424f4f54",
          1017 => x"54494e59",
          1018 => x"2e524f4d",
          1019 => x"00000000",
          1020 => x"01000000",
          2048 => x"0b0b87ff",
          2049 => x"f80d0b0b",
          2050 => x"0b93b904",
          2051 => x"00000000",
          2052 => x"00000000",
          2053 => x"00000000",
          2054 => x"00000000",
          2055 => x"00000000",
          2056 => x"88088c08",
          2057 => x"90088880",
          2058 => x"082d900c",
          2059 => x"8c0c880c",
          2060 => x"04000000",
          2061 => x"00000000",
          2062 => x"00000000",
          2063 => x"00000000",
          2064 => x"71fd0608",
          2065 => x"72830609",
          2066 => x"81058205",
          2067 => x"832b2a83",
          2068 => x"ffff0652",
          2069 => x"04000000",
          2070 => x"00000000",
          2071 => x"00000000",
          2072 => x"71fd0608",
          2073 => x"83ffff73",
          2074 => x"83060981",
          2075 => x"05820583",
          2076 => x"2b2b0906",
          2077 => x"7383ffff",
          2078 => x"0b0b0b0b",
          2079 => x"83a50400",
          2080 => x"72098105",
          2081 => x"72057373",
          2082 => x"09060906",
          2083 => x"73097306",
          2084 => x"070a8106",
          2085 => x"53510400",
          2086 => x"00000000",
          2087 => x"00000000",
          2088 => x"72722473",
          2089 => x"732e0753",
          2090 => x"51040000",
          2091 => x"00000000",
          2092 => x"00000000",
          2093 => x"00000000",
          2094 => x"00000000",
          2095 => x"00000000",
          2096 => x"71737109",
          2097 => x"71068106",
          2098 => x"09810572",
          2099 => x"0a100a72",
          2100 => x"0a100a31",
          2101 => x"050a8106",
          2102 => x"51515351",
          2103 => x"04000000",
          2104 => x"72722673",
          2105 => x"732e0753",
          2106 => x"51040000",
          2107 => x"00000000",
          2108 => x"00000000",
          2109 => x"00000000",
          2110 => x"00000000",
          2111 => x"00000000",
          2112 => x"00000000",
          2113 => x"00000000",
          2114 => x"00000000",
          2115 => x"00000000",
          2116 => x"00000000",
          2117 => x"00000000",
          2118 => x"00000000",
          2119 => x"00000000",
          2120 => x"0b0b0b93",
          2121 => x"9d040000",
          2122 => x"00000000",
          2123 => x"00000000",
          2124 => x"00000000",
          2125 => x"00000000",
          2126 => x"00000000",
          2127 => x"00000000",
          2128 => x"720a722b",
          2129 => x"0a535104",
          2130 => x"00000000",
          2131 => x"00000000",
          2132 => x"00000000",
          2133 => x"00000000",
          2134 => x"00000000",
          2135 => x"00000000",
          2136 => x"72729f06",
          2137 => x"0981050b",
          2138 => x"0b0b9380",
          2139 => x"05040000",
          2140 => x"00000000",
          2141 => x"00000000",
          2142 => x"00000000",
          2143 => x"00000000",
          2144 => x"72722aff",
          2145 => x"739f062a",
          2146 => x"0974090a",
          2147 => x"8106ff05",
          2148 => x"06075351",
          2149 => x"04000000",
          2150 => x"00000000",
          2151 => x"00000000",
          2152 => x"71715351",
          2153 => x"04067383",
          2154 => x"06098105",
          2155 => x"8205832b",
          2156 => x"0b2b0772",
          2157 => x"fc060c51",
          2158 => x"51040000",
          2159 => x"00000000",
          2160 => x"72098105",
          2161 => x"72050970",
          2162 => x"81050906",
          2163 => x"0a810653",
          2164 => x"51040000",
          2165 => x"00000000",
          2166 => x"00000000",
          2167 => x"00000000",
          2168 => x"72098105",
          2169 => x"72050970",
          2170 => x"81050906",
          2171 => x"0a098106",
          2172 => x"53510400",
          2173 => x"00000000",
          2174 => x"00000000",
          2175 => x"00000000",
          2176 => x"71098105",
          2177 => x"52040000",
          2178 => x"00000000",
          2179 => x"00000000",
          2180 => x"00000000",
          2181 => x"00000000",
          2182 => x"00000000",
          2183 => x"00000000",
          2184 => x"72720981",
          2185 => x"05055351",
          2186 => x"04000000",
          2187 => x"00000000",
          2188 => x"00000000",
          2189 => x"00000000",
          2190 => x"00000000",
          2191 => x"00000000",
          2192 => x"72097206",
          2193 => x"73730906",
          2194 => x"07535104",
          2195 => x"00000000",
          2196 => x"00000000",
          2197 => x"00000000",
          2198 => x"00000000",
          2199 => x"00000000",
          2200 => x"71fc0608",
          2201 => x"72830609",
          2202 => x"81058305",
          2203 => x"1010102a",
          2204 => x"81ff0652",
          2205 => x"04000000",
          2206 => x"00000000",
          2207 => x"00000000",
          2208 => x"71fc0608",
          2209 => x"0b0b82ae",
          2210 => x"e4738306",
          2211 => x"10100508",
          2212 => x"060b0b0b",
          2213 => x"93850400",
          2214 => x"00000000",
          2215 => x"00000000",
          2216 => x"88088c08",
          2217 => x"90087575",
          2218 => x"0b0b80c3",
          2219 => x"f42d5050",
          2220 => x"88085690",
          2221 => x"0c8c0c88",
          2222 => x"0c510400",
          2223 => x"00000000",
          2224 => x"88088c08",
          2225 => x"90087575",
          2226 => x"0b0b80c5",
          2227 => x"e02d5050",
          2228 => x"88085690",
          2229 => x"0c8c0c88",
          2230 => x"0c510400",
          2231 => x"00000000",
          2232 => x"72097081",
          2233 => x"0509060a",
          2234 => x"8106ff05",
          2235 => x"70547106",
          2236 => x"73097274",
          2237 => x"05ff0506",
          2238 => x"07515151",
          2239 => x"04000000",
          2240 => x"72097081",
          2241 => x"0509060a",
          2242 => x"098106ff",
          2243 => x"05705471",
          2244 => x"06730972",
          2245 => x"7405ff05",
          2246 => x"06075151",
          2247 => x"51040000",
          2248 => x"05ff0504",
          2249 => x"00000000",
          2250 => x"00000000",
          2251 => x"00000000",
          2252 => x"00000000",
          2253 => x"00000000",
          2254 => x"00000000",
          2255 => x"00000000",
          2256 => x"04000000",
          2257 => x"00000000",
          2258 => x"00000000",
          2259 => x"00000000",
          2260 => x"00000000",
          2261 => x"00000000",
          2262 => x"00000000",
          2263 => x"00000000",
          2264 => x"71810552",
          2265 => x"04000000",
          2266 => x"00000000",
          2267 => x"00000000",
          2268 => x"00000000",
          2269 => x"00000000",
          2270 => x"00000000",
          2271 => x"00000000",
          2272 => x"04000000",
          2273 => x"00000000",
          2274 => x"00000000",
          2275 => x"00000000",
          2276 => x"00000000",
          2277 => x"00000000",
          2278 => x"00000000",
          2279 => x"00000000",
          2280 => x"02840572",
          2281 => x"10100552",
          2282 => x"04000000",
          2283 => x"00000000",
          2284 => x"00000000",
          2285 => x"00000000",
          2286 => x"00000000",
          2287 => x"00000000",
          2288 => x"00000000",
          2289 => x"00000000",
          2290 => x"00000000",
          2291 => x"00000000",
          2292 => x"00000000",
          2293 => x"00000000",
          2294 => x"00000000",
          2295 => x"00000000",
          2296 => x"717105ff",
          2297 => x"05715351",
          2298 => x"020d04ff",
          2299 => x"ffffffff",
          2300 => x"ffffffff",
          2301 => x"ffffffff",
          2302 => x"ffffffff",
          2303 => x"ffffffff",
          2304 => x"00000600",
          2305 => x"ffffffff",
          2306 => x"ffffffff",
          2307 => x"ffffffff",
          2308 => x"ffffffff",
          2309 => x"ffffffff",
          2310 => x"ffffffff",
          2311 => x"ffffffff",
          2312 => x"0b0b0b8c",
          2313 => x"81040b0b",
          2314 => x"0b8c8504",
          2315 => x"0b0b0b8c",
          2316 => x"95040b0b",
          2317 => x"0b8ca404",
          2318 => x"0b0b0b8c",
          2319 => x"b3040b0b",
          2320 => x"0b8cc204",
          2321 => x"0b0b0b8c",
          2322 => x"d1040b0b",
          2323 => x"0b8ce004",
          2324 => x"0b0b0b8c",
          2325 => x"f0040b0b",
          2326 => x"0b8d8004",
          2327 => x"0b0b0b8d",
          2328 => x"8f040b0b",
          2329 => x"0b8d9e04",
          2330 => x"0b0b0b8d",
          2331 => x"ad040b0b",
          2332 => x"0b8dbd04",
          2333 => x"0b0b0b8d",
          2334 => x"cd040b0b",
          2335 => x"0b8ddd04",
          2336 => x"0b0b0b8d",
          2337 => x"ed040b0b",
          2338 => x"0b8dfd04",
          2339 => x"0b0b0b8e",
          2340 => x"8d040b0b",
          2341 => x"0b8e9d04",
          2342 => x"0b0b0b8e",
          2343 => x"ad040b0b",
          2344 => x"0b8ebd04",
          2345 => x"0b0b0b8e",
          2346 => x"cd040b0b",
          2347 => x"0b8edd04",
          2348 => x"0b0b0b8e",
          2349 => x"ed040b0b",
          2350 => x"0b8efd04",
          2351 => x"0b0b0b8f",
          2352 => x"8d040b0b",
          2353 => x"0b8f9d04",
          2354 => x"0b0b0b8f",
          2355 => x"ad040b0b",
          2356 => x"0b8fbd04",
          2357 => x"0b0b0b8f",
          2358 => x"cd040b0b",
          2359 => x"0b8fdd04",
          2360 => x"0b0b0b8f",
          2361 => x"ed040b0b",
          2362 => x"0b8ffd04",
          2363 => x"0b0b0b90",
          2364 => x"8d040b0b",
          2365 => x"0b909d04",
          2366 => x"0b0b0b90",
          2367 => x"ad040b0b",
          2368 => x"0b90bd04",
          2369 => x"0b0b0b90",
          2370 => x"cd040b0b",
          2371 => x"0b90dd04",
          2372 => x"0b0b0b90",
          2373 => x"ed040b0b",
          2374 => x"0b90fd04",
          2375 => x"0b0b0b91",
          2376 => x"8d040b0b",
          2377 => x"0b919d04",
          2378 => x"0b0b0b91",
          2379 => x"ad040b0b",
          2380 => x"0b91bd04",
          2381 => x"0b0b0b91",
          2382 => x"cd040b0b",
          2383 => x"0b91dd04",
          2384 => x"0b0b0b91",
          2385 => x"ed040b0b",
          2386 => x"0b91fd04",
          2387 => x"0b0b0b92",
          2388 => x"8d040b0b",
          2389 => x"0b929d04",
          2390 => x"0b0b0b92",
          2391 => x"ad040b0b",
          2392 => x"0b92bd04",
          2393 => x"0b0b0b92",
          2394 => x"cd04ffff",
          2395 => x"ffffffff",
          2396 => x"ffffffff",
          2397 => x"ffffffff",
          2398 => x"ffffffff",
          2399 => x"ffffffff",
          2400 => x"ffffffff",
          2401 => x"ffffffff",
          2402 => x"ffffffff",
          2403 => x"ffffffff",
          2404 => x"ffffffff",
          2405 => x"ffffffff",
          2406 => x"ffffffff",
          2407 => x"ffffffff",
          2408 => x"ffffffff",
          2409 => x"ffffffff",
          2410 => x"ffffffff",
          2411 => x"ffffffff",
          2412 => x"ffffffff",
          2413 => x"ffffffff",
          2414 => x"ffffffff",
          2415 => x"ffffffff",
          2416 => x"ffffffff",
          2417 => x"ffffffff",
          2418 => x"ffffffff",
          2419 => x"ffffffff",
          2420 => x"ffffffff",
          2421 => x"ffffffff",
          2422 => x"ffffffff",
          2423 => x"ffffffff",
          2424 => x"ffffffff",
          2425 => x"ffffffff",
          2426 => x"ffffffff",
          2427 => x"ffffffff",
          2428 => x"ffffffff",
          2429 => x"ffffffff",
          2430 => x"ffffffff",
          2431 => x"ffffffff",
          2432 => x"04008c81",
          2433 => x"0482d8d4",
          2434 => x"0c80f9b3",
          2435 => x"2d82d8d4",
          2436 => x"08848090",
          2437 => x"0482d8d4",
          2438 => x"0cb3b22d",
          2439 => x"82d8d408",
          2440 => x"84809004",
          2441 => x"82d8d40c",
          2442 => x"afe32d82",
          2443 => x"d8d40884",
          2444 => x"80900482",
          2445 => x"d8d40caf",
          2446 => x"ad2d82d8",
          2447 => x"d4088480",
          2448 => x"900482d8",
          2449 => x"d40c94ad",
          2450 => x"2d82d8d4",
          2451 => x"08848090",
          2452 => x"0482d8d4",
          2453 => x"0cb1c22d",
          2454 => x"82d8d408",
          2455 => x"84809004",
          2456 => x"82d8d40c",
          2457 => x"80cfcc2d",
          2458 => x"82d8d408",
          2459 => x"84809004",
          2460 => x"82d8d40c",
          2461 => x"80c9fb2d",
          2462 => x"82d8d408",
          2463 => x"84809004",
          2464 => x"82d8d40c",
          2465 => x"93d82d82",
          2466 => x"d8d40884",
          2467 => x"80900482",
          2468 => x"d8d40c96",
          2469 => x"c02d82d8",
          2470 => x"d4088480",
          2471 => x"900482d8",
          2472 => x"d40c97cd",
          2473 => x"2d82d8d4",
          2474 => x"08848090",
          2475 => x"0482d8d4",
          2476 => x"0c80fcdd",
          2477 => x"2d82d8d4",
          2478 => x"08848090",
          2479 => x"0482d8d4",
          2480 => x"0c80fdbb",
          2481 => x"2d82d8d4",
          2482 => x"08848090",
          2483 => x"0482d8d4",
          2484 => x"0c80f4f8",
          2485 => x"2d82d8d4",
          2486 => x"08848090",
          2487 => x"0482d8d4",
          2488 => x"0c80f6ef",
          2489 => x"2d82d8d4",
          2490 => x"08848090",
          2491 => x"0482d8d4",
          2492 => x"0c80f8a2",
          2493 => x"2d82d8d4",
          2494 => x"08848090",
          2495 => x"0482d8d4",
          2496 => x"0c81eec7",
          2497 => x"2d82d8d4",
          2498 => x"08848090",
          2499 => x"0482d8d4",
          2500 => x"0c81fbc6",
          2501 => x"2d82d8d4",
          2502 => x"08848090",
          2503 => x"0482d8d4",
          2504 => x"0c81f3ac",
          2505 => x"2d82d8d4",
          2506 => x"08848090",
          2507 => x"0482d8d4",
          2508 => x"0c81f6ac",
          2509 => x"2d82d8d4",
          2510 => x"08848090",
          2511 => x"0482d8d4",
          2512 => x"0c828184",
          2513 => x"2d82d8d4",
          2514 => x"08848090",
          2515 => x"0482d8d4",
          2516 => x"0c8289ed",
          2517 => x"2d82d8d4",
          2518 => x"08848090",
          2519 => x"0482d8d4",
          2520 => x"0c81faa3",
          2521 => x"2d82d8d4",
          2522 => x"08848090",
          2523 => x"0482d8d4",
          2524 => x"0c8284a7",
          2525 => x"2d82d8d4",
          2526 => x"08848090",
          2527 => x"0482d8d4",
          2528 => x"0c8285c7",
          2529 => x"2d82d8d4",
          2530 => x"08848090",
          2531 => x"0482d8d4",
          2532 => x"0c8285e6",
          2533 => x"2d82d8d4",
          2534 => x"08848090",
          2535 => x"0482d8d4",
          2536 => x"0c828dda",
          2537 => x"2d82d8d4",
          2538 => x"08848090",
          2539 => x"0482d8d4",
          2540 => x"0c828bbc",
          2541 => x"2d82d8d4",
          2542 => x"08848090",
          2543 => x"0482d8d4",
          2544 => x"0c8290b6",
          2545 => x"2d82d8d4",
          2546 => x"08848090",
          2547 => x"0482d8d4",
          2548 => x"0c8286ec",
          2549 => x"2d82d8d4",
          2550 => x"08848090",
          2551 => x"0482d8d4",
          2552 => x"0c8293bb",
          2553 => x"2d82d8d4",
          2554 => x"08848090",
          2555 => x"0482d8d4",
          2556 => x"0c8294bc",
          2557 => x"2d82d8d4",
          2558 => x"08848090",
          2559 => x"0482d8d4",
          2560 => x"0c81fca6",
          2561 => x"2d82d8d4",
          2562 => x"08848090",
          2563 => x"0482d8d4",
          2564 => x"0c81fbff",
          2565 => x"2d82d8d4",
          2566 => x"08848090",
          2567 => x"0482d8d4",
          2568 => x"0c81fdaa",
          2569 => x"2d82d8d4",
          2570 => x"08848090",
          2571 => x"0482d8d4",
          2572 => x"0c8287c3",
          2573 => x"2d82d8d4",
          2574 => x"08848090",
          2575 => x"0482d8d4",
          2576 => x"0c8295ad",
          2577 => x"2d82d8d4",
          2578 => x"08848090",
          2579 => x"0482d8d4",
          2580 => x"0c8297b8",
          2581 => x"2d82d8d4",
          2582 => x"08848090",
          2583 => x"0482d8d4",
          2584 => x"0c829abf",
          2585 => x"2d82d8d4",
          2586 => x"08848090",
          2587 => x"0482d8d4",
          2588 => x"0c81ede6",
          2589 => x"2d82d8d4",
          2590 => x"08848090",
          2591 => x"0482d8d4",
          2592 => x"0c829dab",
          2593 => x"2d82d8d4",
          2594 => x"08848090",
          2595 => x"0482d8d4",
          2596 => x"0c82abe0",
          2597 => x"2d82d8d4",
          2598 => x"08848090",
          2599 => x"0482d8d4",
          2600 => x"0c82a9cc",
          2601 => x"2d82d8d4",
          2602 => x"08848090",
          2603 => x"0482d8d4",
          2604 => x"0c81adee",
          2605 => x"2d82d8d4",
          2606 => x"08848090",
          2607 => x"0482d8d4",
          2608 => x"0c81afd8",
          2609 => x"2d82d8d4",
          2610 => x"08848090",
          2611 => x"0482d8d4",
          2612 => x"0c81b1bc",
          2613 => x"2d82d8d4",
          2614 => x"08848090",
          2615 => x"0482d8d4",
          2616 => x"0c80f5a1",
          2617 => x"2d82d8d4",
          2618 => x"08848090",
          2619 => x"0482d8d4",
          2620 => x"0c80f6c5",
          2621 => x"2d82d8d4",
          2622 => x"08848090",
          2623 => x"0482d8d4",
          2624 => x"0c80faa8",
          2625 => x"2d82d8d4",
          2626 => x"08848090",
          2627 => x"0482d8d4",
          2628 => x"0c80d698",
          2629 => x"2d82d8d4",
          2630 => x"08848090",
          2631 => x"0482d8d4",
          2632 => x"0c81a882",
          2633 => x"2d82d8d4",
          2634 => x"08848090",
          2635 => x"0482d8d4",
          2636 => x"0c81a8aa",
          2637 => x"2d82d8d4",
          2638 => x"08848090",
          2639 => x"0482d8d4",
          2640 => x"0c81aca2",
          2641 => x"2d82d8d4",
          2642 => x"08848090",
          2643 => x"0482d8d4",
          2644 => x"0c81a4ec",
          2645 => x"2d82d8d4",
          2646 => x"08848090",
          2647 => x"043c0400",
          2648 => x"00101010",
          2649 => x"10101010",
          2650 => x"10101010",
          2651 => x"10101010",
          2652 => x"10101010",
          2653 => x"10101010",
          2654 => x"10101010",
          2655 => x"10101010",
          2656 => x"53510400",
          2657 => x"007381ff",
          2658 => x"06738306",
          2659 => x"09810583",
          2660 => x"05101010",
          2661 => x"2b0772fc",
          2662 => x"060c5151",
          2663 => x"04727280",
          2664 => x"728106ff",
          2665 => x"05097206",
          2666 => x"05711052",
          2667 => x"720a100a",
          2668 => x"5372ed38",
          2669 => x"51515351",
          2670 => x"0482d8c8",
          2671 => x"7082f4b4",
          2672 => x"278e3880",
          2673 => x"71708405",
          2674 => x"530c0b0b",
          2675 => x"0b93bc04",
          2676 => x"8c815180",
          2677 => x"f3bb0400",
          2678 => x"82d8d408",
          2679 => x"0282d8d4",
          2680 => x"0cfb3d0d",
          2681 => x"82d8d408",
          2682 => x"8c057082",
          2683 => x"d8d408fc",
          2684 => x"050c82d8",
          2685 => x"d408fc05",
          2686 => x"085482d8",
          2687 => x"d4088805",
          2688 => x"085382f4",
          2689 => x"ac085254",
          2690 => x"849a3f82",
          2691 => x"d8c80870",
          2692 => x"82d8d408",
          2693 => x"f8050c82",
          2694 => x"d8d408f8",
          2695 => x"05087082",
          2696 => x"d8c80c51",
          2697 => x"54873d0d",
          2698 => x"82d8d40c",
          2699 => x"0482d8d4",
          2700 => x"080282d8",
          2701 => x"d40cfb3d",
          2702 => x"0d82d8d4",
          2703 => x"08900508",
          2704 => x"85113370",
          2705 => x"81327081",
          2706 => x"06515151",
          2707 => x"52718f38",
          2708 => x"800b82d8",
          2709 => x"d4088c05",
          2710 => x"08258338",
          2711 => x"8d39800b",
          2712 => x"82d8d408",
          2713 => x"f4050c81",
          2714 => x"c43982d8",
          2715 => x"d4088c05",
          2716 => x"08ff0582",
          2717 => x"d8d4088c",
          2718 => x"050c800b",
          2719 => x"82d8d408",
          2720 => x"f8050c82",
          2721 => x"d8d40888",
          2722 => x"050882d8",
          2723 => x"d408fc05",
          2724 => x"0c82d8d4",
          2725 => x"08f80508",
          2726 => x"8a2e80f6",
          2727 => x"38800b82",
          2728 => x"d8d4088c",
          2729 => x"05082580",
          2730 => x"e93882d8",
          2731 => x"d4089005",
          2732 => x"0851a090",
          2733 => x"3f82d8c8",
          2734 => x"087082d8",
          2735 => x"d408f805",
          2736 => x"0c5282d8",
          2737 => x"d408f805",
          2738 => x"08ff2e09",
          2739 => x"81068d38",
          2740 => x"800b82d8",
          2741 => x"d408f405",
          2742 => x"0c80d239",
          2743 => x"82d8d408",
          2744 => x"fc050882",
          2745 => x"d8d408f8",
          2746 => x"05085353",
          2747 => x"71733482",
          2748 => x"d8d4088c",
          2749 => x"0508ff05",
          2750 => x"82d8d408",
          2751 => x"8c050c82",
          2752 => x"d8d408fc",
          2753 => x"05088105",
          2754 => x"82d8d408",
          2755 => x"fc050cff",
          2756 => x"803982d8",
          2757 => x"d408fc05",
          2758 => x"08528072",
          2759 => x"3482d8d4",
          2760 => x"08880508",
          2761 => x"7082d8d4",
          2762 => x"08f4050c",
          2763 => x"5282d8d4",
          2764 => x"08f40508",
          2765 => x"82d8c80c",
          2766 => x"873d0d82",
          2767 => x"d8d40c04",
          2768 => x"82d8d408",
          2769 => x"0282d8d4",
          2770 => x"0cf43d0d",
          2771 => x"860b82d8",
          2772 => x"d408e505",
          2773 => x"3482d8d4",
          2774 => x"08880508",
          2775 => x"82d8d408",
          2776 => x"e0050cfe",
          2777 => x"0a0b82d8",
          2778 => x"d408e805",
          2779 => x"0c82d8d4",
          2780 => x"08900570",
          2781 => x"82d8d408",
          2782 => x"fc050c82",
          2783 => x"d8d408fc",
          2784 => x"05085482",
          2785 => x"d8d4088c",
          2786 => x"05085382",
          2787 => x"d8d408e0",
          2788 => x"05705351",
          2789 => x"54818d3f",
          2790 => x"82d8c808",
          2791 => x"7082d8d4",
          2792 => x"08dc050c",
          2793 => x"82d8d408",
          2794 => x"ec050882",
          2795 => x"d8d40888",
          2796 => x"05080551",
          2797 => x"54807434",
          2798 => x"82d8d408",
          2799 => x"dc050870",
          2800 => x"82d8c80c",
          2801 => x"548e3d0d",
          2802 => x"82d8d40c",
          2803 => x"0482d8d4",
          2804 => x"080282d8",
          2805 => x"d40cfb3d",
          2806 => x"0d82d8d4",
          2807 => x"08900570",
          2808 => x"82d8d408",
          2809 => x"fc050c82",
          2810 => x"d8d408fc",
          2811 => x"05085482",
          2812 => x"d8d4088c",
          2813 => x"05085382",
          2814 => x"d8d40888",
          2815 => x"05085254",
          2816 => x"a33f82d8",
          2817 => x"c8087082",
          2818 => x"d8d408f8",
          2819 => x"050c82d8",
          2820 => x"d408f805",
          2821 => x"087082d8",
          2822 => x"c80c5154",
          2823 => x"873d0d82",
          2824 => x"d8d40c04",
          2825 => x"82d8d408",
          2826 => x"0282d8d4",
          2827 => x"0ced3d0d",
          2828 => x"800b82d8",
          2829 => x"d408e405",
          2830 => x"2382d8d4",
          2831 => x"08880508",
          2832 => x"53800b8c",
          2833 => x"140c82d8",
          2834 => x"d4088805",
          2835 => x"08851133",
          2836 => x"70812a70",
          2837 => x"81327081",
          2838 => x"06515151",
          2839 => x"51537280",
          2840 => x"2e8d38ff",
          2841 => x"0b82d8d4",
          2842 => x"08e0050c",
          2843 => x"96ac3982",
          2844 => x"d8d4088c",
          2845 => x"05085372",
          2846 => x"33537282",
          2847 => x"d8d408f8",
          2848 => x"05347281",
          2849 => x"ff065372",
          2850 => x"802e95fa",
          2851 => x"3882d8d4",
          2852 => x"088c0508",
          2853 => x"810582d8",
          2854 => x"d4088c05",
          2855 => x"0c82d8d4",
          2856 => x"08e40522",
          2857 => x"70810651",
          2858 => x"5372802e",
          2859 => x"958b3882",
          2860 => x"d8d408f8",
          2861 => x"053353af",
          2862 => x"732781fc",
          2863 => x"3882d8d4",
          2864 => x"08f80533",
          2865 => x"5372b926",
          2866 => x"81ee3882",
          2867 => x"d8d408f8",
          2868 => x"05335372",
          2869 => x"b02e0981",
          2870 => x"0680c538",
          2871 => x"82d8d408",
          2872 => x"e8053370",
          2873 => x"982b7098",
          2874 => x"2c515153",
          2875 => x"72b23882",
          2876 => x"d8d408e4",
          2877 => x"05227083",
          2878 => x"2a708132",
          2879 => x"70810651",
          2880 => x"51515372",
          2881 => x"802e9938",
          2882 => x"82d8d408",
          2883 => x"e4052270",
          2884 => x"82800751",
          2885 => x"537282d8",
          2886 => x"d408e405",
          2887 => x"23fed039",
          2888 => x"82d8d408",
          2889 => x"e8053370",
          2890 => x"982b7098",
          2891 => x"2c707083",
          2892 => x"2b721173",
          2893 => x"11515151",
          2894 => x"53515553",
          2895 => x"7282d8d4",
          2896 => x"08e80534",
          2897 => x"82d8d408",
          2898 => x"e8053354",
          2899 => x"82d8d408",
          2900 => x"f8053370",
          2901 => x"15d01151",
          2902 => x"51537282",
          2903 => x"d8d408e8",
          2904 => x"053482d8",
          2905 => x"d408e805",
          2906 => x"3370982b",
          2907 => x"70982c51",
          2908 => x"51537280",
          2909 => x"258b3880",
          2910 => x"ff0b82d8",
          2911 => x"d408e805",
          2912 => x"3482d8d4",
          2913 => x"08e40522",
          2914 => x"70832a70",
          2915 => x"81065151",
          2916 => x"5372fddb",
          2917 => x"3882d8d4",
          2918 => x"08e80533",
          2919 => x"70882b70",
          2920 => x"902b7090",
          2921 => x"2c70882c",
          2922 => x"51515151",
          2923 => x"537282d8",
          2924 => x"d408ec05",
          2925 => x"23fdb839",
          2926 => x"82d8d408",
          2927 => x"e4052270",
          2928 => x"832a7081",
          2929 => x"06515153",
          2930 => x"72802e9d",
          2931 => x"3882d8d4",
          2932 => x"08e80533",
          2933 => x"70982b70",
          2934 => x"982c5151",
          2935 => x"53728a38",
          2936 => x"810b82d8",
          2937 => x"d408e805",
          2938 => x"3482d8d4",
          2939 => x"08f80533",
          2940 => x"e01182d8",
          2941 => x"d408c405",
          2942 => x"0c5382d8",
          2943 => x"d408c405",
          2944 => x"0880d826",
          2945 => x"92943882",
          2946 => x"d8d408c4",
          2947 => x"05087082",
          2948 => x"2b82b0d4",
          2949 => x"11700851",
          2950 => x"51515372",
          2951 => x"0482d8d4",
          2952 => x"08e40522",
          2953 => x"70900751",
          2954 => x"537282d8",
          2955 => x"d408e405",
          2956 => x"2382d8d4",
          2957 => x"08e40522",
          2958 => x"70a00751",
          2959 => x"537282d8",
          2960 => x"d408e405",
          2961 => x"23fca839",
          2962 => x"82d8d408",
          2963 => x"e4052270",
          2964 => x"81800751",
          2965 => x"537282d8",
          2966 => x"d408e405",
          2967 => x"23fc9039",
          2968 => x"82d8d408",
          2969 => x"e4052270",
          2970 => x"80c00751",
          2971 => x"537282d8",
          2972 => x"d408e405",
          2973 => x"23fbf839",
          2974 => x"82d8d408",
          2975 => x"e4052270",
          2976 => x"88075153",
          2977 => x"7282d8d4",
          2978 => x"08e40523",
          2979 => x"800b82d8",
          2980 => x"d408e805",
          2981 => x"34fbd839",
          2982 => x"82d8d408",
          2983 => x"e4052270",
          2984 => x"84075153",
          2985 => x"7282d8d4",
          2986 => x"08e40523",
          2987 => x"fbc139bf",
          2988 => x"0b82d8d4",
          2989 => x"08fc0534",
          2990 => x"82d8d408",
          2991 => x"ec0522ff",
          2992 => x"11515372",
          2993 => x"82d8d408",
          2994 => x"ec052380",
          2995 => x"e30b82d8",
          2996 => x"d408f805",
          2997 => x"348da839",
          2998 => x"82d8d408",
          2999 => x"90050882",
          3000 => x"d8d40890",
          3001 => x"05088405",
          3002 => x"82d8d408",
          3003 => x"90050c70",
          3004 => x"08515372",
          3005 => x"82d8d408",
          3006 => x"fc053482",
          3007 => x"d8d408ec",
          3008 => x"0522ff11",
          3009 => x"51537282",
          3010 => x"d8d408ec",
          3011 => x"05238cef",
          3012 => x"3982d8d4",
          3013 => x"08900508",
          3014 => x"82d8d408",
          3015 => x"90050884",
          3016 => x"0582d8d4",
          3017 => x"0890050c",
          3018 => x"700882d8",
          3019 => x"d408fc05",
          3020 => x"0c82d8d4",
          3021 => x"08e40522",
          3022 => x"70832a70",
          3023 => x"81065151",
          3024 => x"51537280",
          3025 => x"2eab3882",
          3026 => x"d8d408e8",
          3027 => x"05337098",
          3028 => x"2b537298",
          3029 => x"2c5382d8",
          3030 => x"d408fc05",
          3031 => x"085253a2",
          3032 => x"d83f82d8",
          3033 => x"c8085372",
          3034 => x"82d8d408",
          3035 => x"f4052399",
          3036 => x"3982d8d4",
          3037 => x"08fc0508",
          3038 => x"519d8a3f",
          3039 => x"82d8c808",
          3040 => x"537282d8",
          3041 => x"d408f405",
          3042 => x"2382d8d4",
          3043 => x"08ec0522",
          3044 => x"5382d8d4",
          3045 => x"08f40522",
          3046 => x"73713154",
          3047 => x"547282d8",
          3048 => x"d408ec05",
          3049 => x"238bd839",
          3050 => x"82d8d408",
          3051 => x"90050882",
          3052 => x"d8d40890",
          3053 => x"05088405",
          3054 => x"82d8d408",
          3055 => x"90050c70",
          3056 => x"0882d8d4",
          3057 => x"08fc050c",
          3058 => x"82d8d408",
          3059 => x"e4052270",
          3060 => x"832a7081",
          3061 => x"06515151",
          3062 => x"5372802e",
          3063 => x"ab3882d8",
          3064 => x"d408e805",
          3065 => x"3370982b",
          3066 => x"5372982c",
          3067 => x"5382d8d4",
          3068 => x"08fc0508",
          3069 => x"5253a1c1",
          3070 => x"3f82d8c8",
          3071 => x"08537282",
          3072 => x"d8d408f4",
          3073 => x"05239939",
          3074 => x"82d8d408",
          3075 => x"fc050851",
          3076 => x"9bf33f82",
          3077 => x"d8c80853",
          3078 => x"7282d8d4",
          3079 => x"08f40523",
          3080 => x"82d8d408",
          3081 => x"ec052253",
          3082 => x"82d8d408",
          3083 => x"f4052273",
          3084 => x"71315454",
          3085 => x"7282d8d4",
          3086 => x"08ec0523",
          3087 => x"8ac13982",
          3088 => x"d8d408e4",
          3089 => x"05227082",
          3090 => x"2a708106",
          3091 => x"51515372",
          3092 => x"802ea438",
          3093 => x"82d8d408",
          3094 => x"90050882",
          3095 => x"d8d40890",
          3096 => x"05088405",
          3097 => x"82d8d408",
          3098 => x"90050c70",
          3099 => x"0882d8d4",
          3100 => x"08dc050c",
          3101 => x"53a23982",
          3102 => x"d8d40890",
          3103 => x"050882d8",
          3104 => x"d4089005",
          3105 => x"08840582",
          3106 => x"d8d40890",
          3107 => x"050c7008",
          3108 => x"82d8d408",
          3109 => x"dc050c53",
          3110 => x"82d8d408",
          3111 => x"dc050882",
          3112 => x"d8d408fc",
          3113 => x"050c82d8",
          3114 => x"d408fc05",
          3115 => x"088025a4",
          3116 => x"3882d8d4",
          3117 => x"08e40522",
          3118 => x"70820751",
          3119 => x"537282d8",
          3120 => x"d408e405",
          3121 => x"2382d8d4",
          3122 => x"08fc0508",
          3123 => x"3082d8d4",
          3124 => x"08fc050c",
          3125 => x"82d8d408",
          3126 => x"e4052270",
          3127 => x"ffbf0651",
          3128 => x"537282d8",
          3129 => x"d408e405",
          3130 => x"2381af39",
          3131 => x"880b82d8",
          3132 => x"d408f405",
          3133 => x"23a93982",
          3134 => x"d8d408e4",
          3135 => x"05227080",
          3136 => x"c0075153",
          3137 => x"7282d8d4",
          3138 => x"08e40523",
          3139 => x"80f80b82",
          3140 => x"d8d408f8",
          3141 => x"0534900b",
          3142 => x"82d8d408",
          3143 => x"f4052382",
          3144 => x"d8d408e4",
          3145 => x"05227082",
          3146 => x"2a708106",
          3147 => x"51515372",
          3148 => x"802ea438",
          3149 => x"82d8d408",
          3150 => x"90050882",
          3151 => x"d8d40890",
          3152 => x"05088405",
          3153 => x"82d8d408",
          3154 => x"90050c70",
          3155 => x"0882d8d4",
          3156 => x"08d8050c",
          3157 => x"53a23982",
          3158 => x"d8d40890",
          3159 => x"050882d8",
          3160 => x"d4089005",
          3161 => x"08840582",
          3162 => x"d8d40890",
          3163 => x"050c7008",
          3164 => x"82d8d408",
          3165 => x"d8050c53",
          3166 => x"82d8d408",
          3167 => x"d8050882",
          3168 => x"d8d408fc",
          3169 => x"050c82d8",
          3170 => x"d408e405",
          3171 => x"2270cf06",
          3172 => x"51537282",
          3173 => x"d8d408e4",
          3174 => x"052382d8",
          3175 => x"d80b82d8",
          3176 => x"d408f005",
          3177 => x"0c82d8d4",
          3178 => x"08f00508",
          3179 => x"82d8d408",
          3180 => x"f4052282",
          3181 => x"d8d408fc",
          3182 => x"05087155",
          3183 => x"70545654",
          3184 => x"55a3f33f",
          3185 => x"82d8c808",
          3186 => x"53727534",
          3187 => x"82d8d408",
          3188 => x"f0050882",
          3189 => x"d8d408d4",
          3190 => x"050c82d8",
          3191 => x"d408f005",
          3192 => x"08703351",
          3193 => x"53897327",
          3194 => x"a43882d8",
          3195 => x"d408f005",
          3196 => x"08537233",
          3197 => x"5482d8d4",
          3198 => x"08f80533",
          3199 => x"7015df11",
          3200 => x"51515372",
          3201 => x"82d8d408",
          3202 => x"d0053497",
          3203 => x"3982d8d4",
          3204 => x"08f00508",
          3205 => x"537233b0",
          3206 => x"11515372",
          3207 => x"82d8d408",
          3208 => x"d0053482",
          3209 => x"d8d408d4",
          3210 => x"05085382",
          3211 => x"d8d408d0",
          3212 => x"05337334",
          3213 => x"82d8d408",
          3214 => x"f0050881",
          3215 => x"0582d8d4",
          3216 => x"08f0050c",
          3217 => x"82d8d408",
          3218 => x"f4052270",
          3219 => x"5382d8d4",
          3220 => x"08fc0508",
          3221 => x"5253a2ab",
          3222 => x"3f82d8c8",
          3223 => x"087082d8",
          3224 => x"d408fc05",
          3225 => x"0c5382d8",
          3226 => x"d408fc05",
          3227 => x"08802e84",
          3228 => x"38feb239",
          3229 => x"82d8d408",
          3230 => x"f0050882",
          3231 => x"d8d85455",
          3232 => x"72547470",
          3233 => x"75315153",
          3234 => x"7282d8d4",
          3235 => x"08fc0534",
          3236 => x"82d8d408",
          3237 => x"e4052270",
          3238 => x"b2065153",
          3239 => x"72802e94",
          3240 => x"3882d8d4",
          3241 => x"08ec0522",
          3242 => x"ff115153",
          3243 => x"7282d8d4",
          3244 => x"08ec0523",
          3245 => x"82d8d408",
          3246 => x"e4052270",
          3247 => x"862a7081",
          3248 => x"06515153",
          3249 => x"72802e80",
          3250 => x"e73882d8",
          3251 => x"d408ec05",
          3252 => x"2270902b",
          3253 => x"82d8d408",
          3254 => x"cc050c82",
          3255 => x"d8d408cc",
          3256 => x"0508902c",
          3257 => x"82d8d408",
          3258 => x"cc050c82",
          3259 => x"d8d408f4",
          3260 => x"05225153",
          3261 => x"72902e09",
          3262 => x"81069538",
          3263 => x"82d8d408",
          3264 => x"cc0508fe",
          3265 => x"05537282",
          3266 => x"d8d408c8",
          3267 => x"05239339",
          3268 => x"82d8d408",
          3269 => x"cc0508ff",
          3270 => x"05537282",
          3271 => x"d8d408c8",
          3272 => x"052382d8",
          3273 => x"d408c805",
          3274 => x"2282d8d4",
          3275 => x"08ec0523",
          3276 => x"82d8d408",
          3277 => x"e4052270",
          3278 => x"832a7081",
          3279 => x"06515153",
          3280 => x"72802e80",
          3281 => x"d03882d8",
          3282 => x"d408e805",
          3283 => x"3370982b",
          3284 => x"70982c82",
          3285 => x"d8d408fc",
          3286 => x"05335751",
          3287 => x"51537274",
          3288 => x"24973882",
          3289 => x"d8d408e4",
          3290 => x"052270f7",
          3291 => x"06515372",
          3292 => x"82d8d408",
          3293 => x"e405239d",
          3294 => x"3982d8d4",
          3295 => x"08e80533",
          3296 => x"5382d8d4",
          3297 => x"08fc0533",
          3298 => x"73713154",
          3299 => x"547282d8",
          3300 => x"d408e805",
          3301 => x"3482d8d4",
          3302 => x"08e40522",
          3303 => x"70832a70",
          3304 => x"81065151",
          3305 => x"5372802e",
          3306 => x"b13882d8",
          3307 => x"d408e805",
          3308 => x"3370882b",
          3309 => x"70902b70",
          3310 => x"902c7088",
          3311 => x"2c515151",
          3312 => x"51537254",
          3313 => x"82d8d408",
          3314 => x"ec052270",
          3315 => x"75315153",
          3316 => x"7282d8d4",
          3317 => x"08ec0523",
          3318 => x"af3982d8",
          3319 => x"d408fc05",
          3320 => x"3370882b",
          3321 => x"70902b70",
          3322 => x"902c7088",
          3323 => x"2c515151",
          3324 => x"51537254",
          3325 => x"82d8d408",
          3326 => x"ec052270",
          3327 => x"75315153",
          3328 => x"7282d8d4",
          3329 => x"08ec0523",
          3330 => x"82d8d408",
          3331 => x"e4052270",
          3332 => x"83800651",
          3333 => x"5372b038",
          3334 => x"82d8d408",
          3335 => x"ec0522ff",
          3336 => x"11545472",
          3337 => x"82d8d408",
          3338 => x"ec052373",
          3339 => x"902b7090",
          3340 => x"2c515380",
          3341 => x"73259038",
          3342 => x"82d8d408",
          3343 => x"88050852",
          3344 => x"a0518aee",
          3345 => x"3fd23982",
          3346 => x"d8d408e4",
          3347 => x"05227081",
          3348 => x"2a708106",
          3349 => x"51515372",
          3350 => x"802e9138",
          3351 => x"82d8d408",
          3352 => x"88050852",
          3353 => x"ad518aca",
          3354 => x"3f80c739",
          3355 => x"82d8d408",
          3356 => x"e4052270",
          3357 => x"842a7081",
          3358 => x"06515153",
          3359 => x"72802e90",
          3360 => x"3882d8d4",
          3361 => x"08880508",
          3362 => x"52ab518a",
          3363 => x"a53fa339",
          3364 => x"82d8d408",
          3365 => x"e4052270",
          3366 => x"852a7081",
          3367 => x"06515153",
          3368 => x"72802e8e",
          3369 => x"3882d8d4",
          3370 => x"08880508",
          3371 => x"52a0518a",
          3372 => x"813f82d8",
          3373 => x"d408e405",
          3374 => x"2270862a",
          3375 => x"70810651",
          3376 => x"51537280",
          3377 => x"2eb13882",
          3378 => x"d8d40888",
          3379 => x"050852b0",
          3380 => x"5189df3f",
          3381 => x"82d8d408",
          3382 => x"f4052253",
          3383 => x"72902e09",
          3384 => x"81069438",
          3385 => x"82d8d408",
          3386 => x"88050852",
          3387 => x"82d8d408",
          3388 => x"f8053351",
          3389 => x"89bc3f82",
          3390 => x"d8d408e4",
          3391 => x"05227088",
          3392 => x"2a708106",
          3393 => x"51515372",
          3394 => x"802eb038",
          3395 => x"82d8d408",
          3396 => x"ec0522ff",
          3397 => x"11545472",
          3398 => x"82d8d408",
          3399 => x"ec052373",
          3400 => x"902b7090",
          3401 => x"2c515380",
          3402 => x"73259038",
          3403 => x"82d8d408",
          3404 => x"88050852",
          3405 => x"b05188fa",
          3406 => x"3fd23982",
          3407 => x"d8d408e4",
          3408 => x"05227083",
          3409 => x"2a708106",
          3410 => x"51515372",
          3411 => x"802eb038",
          3412 => x"82d8d408",
          3413 => x"e80533ff",
          3414 => x"11545472",
          3415 => x"82d8d408",
          3416 => x"e8053473",
          3417 => x"982b7098",
          3418 => x"2c515380",
          3419 => x"73259038",
          3420 => x"82d8d408",
          3421 => x"88050852",
          3422 => x"b05188b6",
          3423 => x"3fd23982",
          3424 => x"d8d408e4",
          3425 => x"05227087",
          3426 => x"2a708106",
          3427 => x"51515372",
          3428 => x"b03882d8",
          3429 => x"d408ec05",
          3430 => x"22ff1154",
          3431 => x"547282d8",
          3432 => x"d408ec05",
          3433 => x"2373902b",
          3434 => x"70902c51",
          3435 => x"53807325",
          3436 => x"903882d8",
          3437 => x"d4088805",
          3438 => x"0852a051",
          3439 => x"87f43fd2",
          3440 => x"3982d8d4",
          3441 => x"08f80533",
          3442 => x"537280e3",
          3443 => x"2e098106",
          3444 => x"973882d8",
          3445 => x"d4088805",
          3446 => x"085282d8",
          3447 => x"d408fc05",
          3448 => x"335187ce",
          3449 => x"3f81ee39",
          3450 => x"82d8d408",
          3451 => x"f8053353",
          3452 => x"7280f32e",
          3453 => x"09810680",
          3454 => x"cb3882d8",
          3455 => x"d408f405",
          3456 => x"22ff1151",
          3457 => x"537282d8",
          3458 => x"d408f405",
          3459 => x"237283ff",
          3460 => x"ff065372",
          3461 => x"83ffff2e",
          3462 => x"81bb3882",
          3463 => x"d8d40888",
          3464 => x"05085282",
          3465 => x"d8d408fc",
          3466 => x"05087033",
          3467 => x"5282d8d4",
          3468 => x"08fc0508",
          3469 => x"810582d8",
          3470 => x"d408fc05",
          3471 => x"0c5386f2",
          3472 => x"3fffb739",
          3473 => x"82d8d408",
          3474 => x"f8053353",
          3475 => x"7280d32e",
          3476 => x"09810680",
          3477 => x"cb3882d8",
          3478 => x"d408f405",
          3479 => x"22ff1151",
          3480 => x"537282d8",
          3481 => x"d408f405",
          3482 => x"237283ff",
          3483 => x"ff065372",
          3484 => x"83ffff2e",
          3485 => x"80df3882",
          3486 => x"d8d40888",
          3487 => x"05085282",
          3488 => x"d8d408fc",
          3489 => x"05087033",
          3490 => x"525386a6",
          3491 => x"3f82d8d4",
          3492 => x"08fc0508",
          3493 => x"810582d8",
          3494 => x"d408fc05",
          3495 => x"0cffb739",
          3496 => x"82d8d408",
          3497 => x"f0050882",
          3498 => x"d8d82ea9",
          3499 => x"3882d8d4",
          3500 => x"08880508",
          3501 => x"5282d8d4",
          3502 => x"08f00508",
          3503 => x"ff0582d8",
          3504 => x"d408f005",
          3505 => x"0c82d8d4",
          3506 => x"08f00508",
          3507 => x"70335253",
          3508 => x"85e03fcc",
          3509 => x"3982d8d4",
          3510 => x"08e40522",
          3511 => x"70872a70",
          3512 => x"81065151",
          3513 => x"5372802e",
          3514 => x"80c33882",
          3515 => x"d8d408ec",
          3516 => x"0522ff11",
          3517 => x"54547282",
          3518 => x"d8d408ec",
          3519 => x"05237390",
          3520 => x"2b70902c",
          3521 => x"51538073",
          3522 => x"25a33882",
          3523 => x"d8d40888",
          3524 => x"050852a0",
          3525 => x"51859b3f",
          3526 => x"d23982d8",
          3527 => x"d4088805",
          3528 => x"085282d8",
          3529 => x"d408f805",
          3530 => x"33518586",
          3531 => x"3f800b82",
          3532 => x"d8d408e4",
          3533 => x"0523eab7",
          3534 => x"3982d8d4",
          3535 => x"08f80533",
          3536 => x"5372a52e",
          3537 => x"098106a8",
          3538 => x"38810b82",
          3539 => x"d8d408e4",
          3540 => x"0523800b",
          3541 => x"82d8d408",
          3542 => x"ec052380",
          3543 => x"0b82d8d4",
          3544 => x"08e80534",
          3545 => x"8a0b82d8",
          3546 => x"d408f405",
          3547 => x"23ea8039",
          3548 => x"82d8d408",
          3549 => x"88050852",
          3550 => x"82d8d408",
          3551 => x"f8053351",
          3552 => x"84b03fe9",
          3553 => x"ea3982d8",
          3554 => x"d4088805",
          3555 => x"088c1108",
          3556 => x"7082d8d4",
          3557 => x"08e0050c",
          3558 => x"515382d8",
          3559 => x"d408e005",
          3560 => x"0882d8c8",
          3561 => x"0c953d0d",
          3562 => x"82d8d40c",
          3563 => x"0482d8d4",
          3564 => x"080282d8",
          3565 => x"d40cfd3d",
          3566 => x"0d82f4a8",
          3567 => x"085382d8",
          3568 => x"d4088c05",
          3569 => x"085282d8",
          3570 => x"d4088805",
          3571 => x"0851e4dd",
          3572 => x"3f82d8c8",
          3573 => x"087082d8",
          3574 => x"c80c5485",
          3575 => x"3d0d82d8",
          3576 => x"d40c0482",
          3577 => x"d8d40802",
          3578 => x"82d8d40c",
          3579 => x"fb3d0d80",
          3580 => x"0b82d8d4",
          3581 => x"08f8050c",
          3582 => x"82f4ac08",
          3583 => x"85113370",
          3584 => x"812a7081",
          3585 => x"32708106",
          3586 => x"51515151",
          3587 => x"5372802e",
          3588 => x"8d38ff0b",
          3589 => x"82d8d408",
          3590 => x"f4050c81",
          3591 => x"923982d8",
          3592 => x"d4088805",
          3593 => x"08537233",
          3594 => x"82d8d408",
          3595 => x"88050881",
          3596 => x"0582d8d4",
          3597 => x"0888050c",
          3598 => x"537282d8",
          3599 => x"d408fc05",
          3600 => x"347281ff",
          3601 => x"06537280",
          3602 => x"2eb03882",
          3603 => x"f4ac0882",
          3604 => x"f4ac0853",
          3605 => x"82d8d408",
          3606 => x"fc053352",
          3607 => x"90110851",
          3608 => x"53722d82",
          3609 => x"d8c80853",
          3610 => x"72802eff",
          3611 => x"b138ff0b",
          3612 => x"82d8d408",
          3613 => x"f8050cff",
          3614 => x"a53982f4",
          3615 => x"ac0882f4",
          3616 => x"ac085353",
          3617 => x"8a519013",
          3618 => x"0853722d",
          3619 => x"82d8c808",
          3620 => x"5372802e",
          3621 => x"8a38ff0b",
          3622 => x"82d8d408",
          3623 => x"f8050c82",
          3624 => x"d8d408f8",
          3625 => x"05087082",
          3626 => x"d8d408f4",
          3627 => x"050c5382",
          3628 => x"d8d408f4",
          3629 => x"050882d8",
          3630 => x"c80c873d",
          3631 => x"0d82d8d4",
          3632 => x"0c0482d8",
          3633 => x"d4080282",
          3634 => x"d8d40cfb",
          3635 => x"3d0d800b",
          3636 => x"82d8d408",
          3637 => x"f8050c82",
          3638 => x"d8d4088c",
          3639 => x"05088511",
          3640 => x"3370812a",
          3641 => x"70813270",
          3642 => x"81065151",
          3643 => x"51515372",
          3644 => x"802e8d38",
          3645 => x"ff0b82d8",
          3646 => x"d408f405",
          3647 => x"0c80f339",
          3648 => x"82d8d408",
          3649 => x"88050853",
          3650 => x"723382d8",
          3651 => x"d4088805",
          3652 => x"08810582",
          3653 => x"d8d40888",
          3654 => x"050c5372",
          3655 => x"82d8d408",
          3656 => x"fc053472",
          3657 => x"81ff0653",
          3658 => x"72802eb6",
          3659 => x"3882d8d4",
          3660 => x"088c0508",
          3661 => x"82d8d408",
          3662 => x"8c050853",
          3663 => x"82d8d408",
          3664 => x"fc053352",
          3665 => x"90110851",
          3666 => x"53722d82",
          3667 => x"d8c80853",
          3668 => x"72802eff",
          3669 => x"ab38ff0b",
          3670 => x"82d8d408",
          3671 => x"f8050cff",
          3672 => x"9f3982d8",
          3673 => x"d408f805",
          3674 => x"087082d8",
          3675 => x"d408f405",
          3676 => x"0c5382d8",
          3677 => x"d408f405",
          3678 => x"0882d8c8",
          3679 => x"0c873d0d",
          3680 => x"82d8d40c",
          3681 => x"0482d8d4",
          3682 => x"080282d8",
          3683 => x"d40cfe3d",
          3684 => x"0d82f4ac",
          3685 => x"085282d8",
          3686 => x"d4088805",
          3687 => x"0851933f",
          3688 => x"82d8c808",
          3689 => x"7082d8c8",
          3690 => x"0c53843d",
          3691 => x"0d82d8d4",
          3692 => x"0c0482d8",
          3693 => x"d4080282",
          3694 => x"d8d40cfb",
          3695 => x"3d0d82d8",
          3696 => x"d4088c05",
          3697 => x"08851133",
          3698 => x"70812a70",
          3699 => x"81327081",
          3700 => x"06515151",
          3701 => x"51537280",
          3702 => x"2e8d38ff",
          3703 => x"0b82d8d4",
          3704 => x"08fc050c",
          3705 => x"81cb3982",
          3706 => x"d8d4088c",
          3707 => x"05088511",
          3708 => x"3370822a",
          3709 => x"70810651",
          3710 => x"51515372",
          3711 => x"802e80db",
          3712 => x"3882d8d4",
          3713 => x"088c0508",
          3714 => x"82d8d408",
          3715 => x"8c050854",
          3716 => x"548c1408",
          3717 => x"88140825",
          3718 => x"9f3882d8",
          3719 => x"d4088c05",
          3720 => x"08700870",
          3721 => x"82d8d408",
          3722 => x"88050852",
          3723 => x"57545472",
          3724 => x"75347308",
          3725 => x"8105740c",
          3726 => x"82d8d408",
          3727 => x"8c05088c",
          3728 => x"11088105",
          3729 => x"8c120c82",
          3730 => x"d8d40888",
          3731 => x"05087082",
          3732 => x"d8d408fc",
          3733 => x"050c5153",
          3734 => x"80d73982",
          3735 => x"d8d4088c",
          3736 => x"050882d8",
          3737 => x"d4088c05",
          3738 => x"085382d8",
          3739 => x"d4088805",
          3740 => x"087081ff",
          3741 => x"06539012",
          3742 => x"08515454",
          3743 => x"722d82d8",
          3744 => x"c8085372",
          3745 => x"a33882d8",
          3746 => x"d4088c05",
          3747 => x"088c1108",
          3748 => x"81058c12",
          3749 => x"0c82d8d4",
          3750 => x"08880508",
          3751 => x"7082d8d4",
          3752 => x"08fc050c",
          3753 => x"51538a39",
          3754 => x"ff0b82d8",
          3755 => x"d408fc05",
          3756 => x"0c82d8d4",
          3757 => x"08fc0508",
          3758 => x"82d8c80c",
          3759 => x"873d0d82",
          3760 => x"d8d40c04",
          3761 => x"82d8d408",
          3762 => x"0282d8d4",
          3763 => x"0cf93d0d",
          3764 => x"82d8d408",
          3765 => x"88050885",
          3766 => x"11337081",
          3767 => x"32708106",
          3768 => x"51515152",
          3769 => x"71802e8d",
          3770 => x"38ff0b82",
          3771 => x"d8d408f8",
          3772 => x"050c8394",
          3773 => x"3982d8d4",
          3774 => x"08880508",
          3775 => x"85113370",
          3776 => x"862a7081",
          3777 => x"06515151",
          3778 => x"5271802e",
          3779 => x"80c53882",
          3780 => x"d8d40888",
          3781 => x"050882d8",
          3782 => x"d4088805",
          3783 => x"08535385",
          3784 => x"123370ff",
          3785 => x"bf065152",
          3786 => x"71851434",
          3787 => x"82d8d408",
          3788 => x"8805088c",
          3789 => x"11088105",
          3790 => x"8c120c82",
          3791 => x"d8d40888",
          3792 => x"05088411",
          3793 => x"337082d8",
          3794 => x"d408f805",
          3795 => x"0c515152",
          3796 => x"82b63982",
          3797 => x"d8d40888",
          3798 => x"05088511",
          3799 => x"3370822a",
          3800 => x"70810651",
          3801 => x"51515271",
          3802 => x"802e80d7",
          3803 => x"3882d8d4",
          3804 => x"08880508",
          3805 => x"70087033",
          3806 => x"82d8d408",
          3807 => x"fc050c51",
          3808 => x"5282d8d4",
          3809 => x"08fc0508",
          3810 => x"a93882d8",
          3811 => x"d4088805",
          3812 => x"0882d8d4",
          3813 => x"08880508",
          3814 => x"53538512",
          3815 => x"3370a007",
          3816 => x"51527185",
          3817 => x"1434ff0b",
          3818 => x"82d8d408",
          3819 => x"f8050c81",
          3820 => x"d73982d8",
          3821 => x"d4088805",
          3822 => x"08700881",
          3823 => x"05710c52",
          3824 => x"81a13982",
          3825 => x"d8d40888",
          3826 => x"050882d8",
          3827 => x"d4088805",
          3828 => x"08529411",
          3829 => x"08515271",
          3830 => x"2d82d8c8",
          3831 => x"087082d8",
          3832 => x"d408fc05",
          3833 => x"0c5282d8",
          3834 => x"d408fc05",
          3835 => x"08802580",
          3836 => x"f23882d8",
          3837 => x"d4088805",
          3838 => x"0882d8d4",
          3839 => x"08f4050c",
          3840 => x"82d8d408",
          3841 => x"88050885",
          3842 => x"113382d8",
          3843 => x"d408f005",
          3844 => x"0c5282d8",
          3845 => x"d408fc05",
          3846 => x"08ff2e09",
          3847 => x"81069538",
          3848 => x"82d8d408",
          3849 => x"f0050890",
          3850 => x"07527182",
          3851 => x"d8d408ec",
          3852 => x"05349339",
          3853 => x"82d8d408",
          3854 => x"f00508a0",
          3855 => x"07527182",
          3856 => x"d8d408ec",
          3857 => x"053482d8",
          3858 => x"d408f405",
          3859 => x"085282d8",
          3860 => x"d408ec05",
          3861 => x"33851334",
          3862 => x"ff0b82d8",
          3863 => x"d408f805",
          3864 => x"0ca63982",
          3865 => x"d8d40888",
          3866 => x"05088c11",
          3867 => x"0881058c",
          3868 => x"120c82d8",
          3869 => x"d408fc05",
          3870 => x"087081ff",
          3871 => x"067082d8",
          3872 => x"d408f805",
          3873 => x"0c515152",
          3874 => x"82d8d408",
          3875 => x"f8050882",
          3876 => x"d8c80c89",
          3877 => x"3d0d82d8",
          3878 => x"d40c0482",
          3879 => x"d8d40802",
          3880 => x"82d8d40c",
          3881 => x"fd3d0d82",
          3882 => x"d8d40888",
          3883 => x"050882d8",
          3884 => x"d408fc05",
          3885 => x"0c82d8d4",
          3886 => x"088c0508",
          3887 => x"82d8d408",
          3888 => x"f8050c82",
          3889 => x"d8d40890",
          3890 => x"0508802e",
          3891 => x"82a23882",
          3892 => x"d8d408f8",
          3893 => x"050882d8",
          3894 => x"d408fc05",
          3895 => x"082681ac",
          3896 => x"3882d8d4",
          3897 => x"08f80508",
          3898 => x"82d8d408",
          3899 => x"90050805",
          3900 => x"5182d8d4",
          3901 => x"08fc0508",
          3902 => x"71278190",
          3903 => x"3882d8d4",
          3904 => x"08fc0508",
          3905 => x"82d8d408",
          3906 => x"90050805",
          3907 => x"82d8d408",
          3908 => x"fc050c82",
          3909 => x"d8d408f8",
          3910 => x"050882d8",
          3911 => x"d4089005",
          3912 => x"080582d8",
          3913 => x"d408f805",
          3914 => x"0c82d8d4",
          3915 => x"08900508",
          3916 => x"810582d8",
          3917 => x"d4089005",
          3918 => x"0c82d8d4",
          3919 => x"08900508",
          3920 => x"ff0582d8",
          3921 => x"d4089005",
          3922 => x"0c82d8d4",
          3923 => x"08900508",
          3924 => x"802e819c",
          3925 => x"3882d8d4",
          3926 => x"08fc0508",
          3927 => x"ff0582d8",
          3928 => x"d408fc05",
          3929 => x"0c82d8d4",
          3930 => x"08f80508",
          3931 => x"ff0582d8",
          3932 => x"d408f805",
          3933 => x"0c82d8d4",
          3934 => x"08fc0508",
          3935 => x"82d8d408",
          3936 => x"f8050853",
          3937 => x"51713371",
          3938 => x"34ffae39",
          3939 => x"82d8d408",
          3940 => x"90050881",
          3941 => x"0582d8d4",
          3942 => x"0890050c",
          3943 => x"82d8d408",
          3944 => x"900508ff",
          3945 => x"0582d8d4",
          3946 => x"0890050c",
          3947 => x"82d8d408",
          3948 => x"90050880",
          3949 => x"2eba3882",
          3950 => x"d8d408f8",
          3951 => x"05085170",
          3952 => x"3382d8d4",
          3953 => x"08f80508",
          3954 => x"810582d8",
          3955 => x"d408f805",
          3956 => x"0c82d8d4",
          3957 => x"08fc0508",
          3958 => x"52527171",
          3959 => x"3482d8d4",
          3960 => x"08fc0508",
          3961 => x"810582d8",
          3962 => x"d408fc05",
          3963 => x"0cffad39",
          3964 => x"82d8d408",
          3965 => x"88050870",
          3966 => x"82d8c80c",
          3967 => x"51853d0d",
          3968 => x"82d8d40c",
          3969 => x"0482d8d4",
          3970 => x"080282d8",
          3971 => x"d40cfe3d",
          3972 => x"0d82d8d4",
          3973 => x"08880508",
          3974 => x"82d8d408",
          3975 => x"fc050c82",
          3976 => x"d8d408fc",
          3977 => x"05085271",
          3978 => x"3382d8d4",
          3979 => x"08fc0508",
          3980 => x"810582d8",
          3981 => x"d408fc05",
          3982 => x"0c7081ff",
          3983 => x"06515170",
          3984 => x"802e8338",
          3985 => x"da3982d8",
          3986 => x"d408fc05",
          3987 => x"08ff0582",
          3988 => x"d8d408fc",
          3989 => x"050c82d8",
          3990 => x"d408fc05",
          3991 => x"0882d8d4",
          3992 => x"08880508",
          3993 => x"317082d8",
          3994 => x"c80c5184",
          3995 => x"3d0d82d8",
          3996 => x"d40c0482",
          3997 => x"d8d40802",
          3998 => x"82d8d40c",
          3999 => x"fe3d0d82",
          4000 => x"d8d40888",
          4001 => x"050882d8",
          4002 => x"d408fc05",
          4003 => x"0c82d8d4",
          4004 => x"088c0508",
          4005 => x"52713382",
          4006 => x"d8d4088c",
          4007 => x"05088105",
          4008 => x"82d8d408",
          4009 => x"8c050c82",
          4010 => x"d8d408fc",
          4011 => x"05085351",
          4012 => x"70723482",
          4013 => x"d8d408fc",
          4014 => x"05088105",
          4015 => x"82d8d408",
          4016 => x"fc050c70",
          4017 => x"81ff0651",
          4018 => x"70802e84",
          4019 => x"38ffbe39",
          4020 => x"82d8d408",
          4021 => x"88050870",
          4022 => x"82d8c80c",
          4023 => x"51843d0d",
          4024 => x"82d8d40c",
          4025 => x"0482d8d4",
          4026 => x"080282d8",
          4027 => x"d40cfd3d",
          4028 => x"0d82d8d4",
          4029 => x"08880508",
          4030 => x"82d8d408",
          4031 => x"fc050c82",
          4032 => x"d8d4088c",
          4033 => x"050882d8",
          4034 => x"d408f805",
          4035 => x"0c82d8d4",
          4036 => x"08900508",
          4037 => x"802e80e5",
          4038 => x"3882d8d4",
          4039 => x"08900508",
          4040 => x"810582d8",
          4041 => x"d4089005",
          4042 => x"0c82d8d4",
          4043 => x"08900508",
          4044 => x"ff0582d8",
          4045 => x"d4089005",
          4046 => x"0c82d8d4",
          4047 => x"08900508",
          4048 => x"802eba38",
          4049 => x"82d8d408",
          4050 => x"f8050851",
          4051 => x"703382d8",
          4052 => x"d408f805",
          4053 => x"08810582",
          4054 => x"d8d408f8",
          4055 => x"050c82d8",
          4056 => x"d408fc05",
          4057 => x"08525271",
          4058 => x"713482d8",
          4059 => x"d408fc05",
          4060 => x"08810582",
          4061 => x"d8d408fc",
          4062 => x"050cffad",
          4063 => x"3982d8d4",
          4064 => x"08880508",
          4065 => x"7082d8c8",
          4066 => x"0c51853d",
          4067 => x"0d82d8d4",
          4068 => x"0c0482d8",
          4069 => x"d4080282",
          4070 => x"d8d40cfd",
          4071 => x"3d0d82d8",
          4072 => x"d4089005",
          4073 => x"08802e81",
          4074 => x"f43882d8",
          4075 => x"d4088c05",
          4076 => x"08527133",
          4077 => x"82d8d408",
          4078 => x"8c050881",
          4079 => x"0582d8d4",
          4080 => x"088c050c",
          4081 => x"82d8d408",
          4082 => x"88050870",
          4083 => x"337281ff",
          4084 => x"06535454",
          4085 => x"5171712e",
          4086 => x"843880ce",
          4087 => x"3982d8d4",
          4088 => x"08880508",
          4089 => x"52713382",
          4090 => x"d8d40888",
          4091 => x"05088105",
          4092 => x"82d8d408",
          4093 => x"88050c70",
          4094 => x"81ff0651",
          4095 => x"51708d38",
          4096 => x"800b82d8",
          4097 => x"d408fc05",
          4098 => x"0c819b39",
          4099 => x"82d8d408",
          4100 => x"900508ff",
          4101 => x"0582d8d4",
          4102 => x"0890050c",
          4103 => x"82d8d408",
          4104 => x"90050880",
          4105 => x"2e8438ff",
          4106 => x"813982d8",
          4107 => x"d4089005",
          4108 => x"08802e80",
          4109 => x"e83882d8",
          4110 => x"d4088805",
          4111 => x"08703352",
          4112 => x"53708d38",
          4113 => x"ff0b82d8",
          4114 => x"d408fc05",
          4115 => x"0c80d739",
          4116 => x"82d8d408",
          4117 => x"8c0508ff",
          4118 => x"0582d8d4",
          4119 => x"088c050c",
          4120 => x"82d8d408",
          4121 => x"8c050870",
          4122 => x"33525270",
          4123 => x"8c38810b",
          4124 => x"82d8d408",
          4125 => x"fc050cae",
          4126 => x"3982d8d4",
          4127 => x"08880508",
          4128 => x"703382d8",
          4129 => x"d4088c05",
          4130 => x"08703372",
          4131 => x"71317082",
          4132 => x"d8d408fc",
          4133 => x"050c5355",
          4134 => x"5252538a",
          4135 => x"39800b82",
          4136 => x"d8d408fc",
          4137 => x"050c82d8",
          4138 => x"d408fc05",
          4139 => x"0882d8c8",
          4140 => x"0c853d0d",
          4141 => x"82d8d40c",
          4142 => x"0482d8d4",
          4143 => x"080282d8",
          4144 => x"d40cfd3d",
          4145 => x"0d82d8d4",
          4146 => x"08880508",
          4147 => x"82d8d408",
          4148 => x"f8050c82",
          4149 => x"d8d4088c",
          4150 => x"05088d38",
          4151 => x"800b82d8",
          4152 => x"d408fc05",
          4153 => x"0c80ec39",
          4154 => x"82d8d408",
          4155 => x"f8050852",
          4156 => x"713382d8",
          4157 => x"d408f805",
          4158 => x"08810582",
          4159 => x"d8d408f8",
          4160 => x"050c7081",
          4161 => x"ff065151",
          4162 => x"70802e9f",
          4163 => x"3882d8d4",
          4164 => x"088c0508",
          4165 => x"ff0582d8",
          4166 => x"d4088c05",
          4167 => x"0c82d8d4",
          4168 => x"088c0508",
          4169 => x"ff2e8438",
          4170 => x"ffbe3982",
          4171 => x"d8d408f8",
          4172 => x"0508ff05",
          4173 => x"82d8d408",
          4174 => x"f8050c82",
          4175 => x"d8d408f8",
          4176 => x"050882d8",
          4177 => x"d4088805",
          4178 => x"08317082",
          4179 => x"d8d408fc",
          4180 => x"050c5182",
          4181 => x"d8d408fc",
          4182 => x"050882d8",
          4183 => x"c80c853d",
          4184 => x"0d82d8d4",
          4185 => x"0c0482d8",
          4186 => x"d4080282",
          4187 => x"d8d40cfe",
          4188 => x"3d0d82d8",
          4189 => x"d4088805",
          4190 => x"0882d8d4",
          4191 => x"08fc050c",
          4192 => x"82d8d408",
          4193 => x"90050880",
          4194 => x"2e80d438",
          4195 => x"82d8d408",
          4196 => x"90050881",
          4197 => x"0582d8d4",
          4198 => x"0890050c",
          4199 => x"82d8d408",
          4200 => x"900508ff",
          4201 => x"0582d8d4",
          4202 => x"0890050c",
          4203 => x"82d8d408",
          4204 => x"90050880",
          4205 => x"2ea93882",
          4206 => x"d8d4088c",
          4207 => x"05085170",
          4208 => x"82d8d408",
          4209 => x"fc050852",
          4210 => x"52717134",
          4211 => x"82d8d408",
          4212 => x"fc050881",
          4213 => x"0582d8d4",
          4214 => x"08fc050c",
          4215 => x"ffbe3982",
          4216 => x"d8d40888",
          4217 => x"05087082",
          4218 => x"d8c80c51",
          4219 => x"843d0d82",
          4220 => x"d8d40c04",
          4221 => x"82d8d408",
          4222 => x"0282d8d4",
          4223 => x"0cf93d0d",
          4224 => x"800b82d8",
          4225 => x"d408fc05",
          4226 => x"0c82d8d4",
          4227 => x"08880508",
          4228 => x"8025b938",
          4229 => x"82d8d408",
          4230 => x"88050830",
          4231 => x"82d8d408",
          4232 => x"88050c80",
          4233 => x"0b82d8d4",
          4234 => x"08f4050c",
          4235 => x"82d8d408",
          4236 => x"fc05088a",
          4237 => x"38810b82",
          4238 => x"d8d408f4",
          4239 => x"050c82d8",
          4240 => x"d408f405",
          4241 => x"0882d8d4",
          4242 => x"08fc050c",
          4243 => x"82d8d408",
          4244 => x"8c050880",
          4245 => x"25b93882",
          4246 => x"d8d4088c",
          4247 => x"05083082",
          4248 => x"d8d4088c",
          4249 => x"050c800b",
          4250 => x"82d8d408",
          4251 => x"f0050c82",
          4252 => x"d8d408fc",
          4253 => x"05088a38",
          4254 => x"810b82d8",
          4255 => x"d408f005",
          4256 => x"0c82d8d4",
          4257 => x"08f00508",
          4258 => x"82d8d408",
          4259 => x"fc050c80",
          4260 => x"5382d8d4",
          4261 => x"088c0508",
          4262 => x"5282d8d4",
          4263 => x"08880508",
          4264 => x"5182c53f",
          4265 => x"82d8c808",
          4266 => x"7082d8d4",
          4267 => x"08f8050c",
          4268 => x"5482d8d4",
          4269 => x"08fc0508",
          4270 => x"802e9038",
          4271 => x"82d8d408",
          4272 => x"f8050830",
          4273 => x"82d8d408",
          4274 => x"f8050c82",
          4275 => x"d8d408f8",
          4276 => x"05087082",
          4277 => x"d8c80c54",
          4278 => x"893d0d82",
          4279 => x"d8d40c04",
          4280 => x"82d8d408",
          4281 => x"0282d8d4",
          4282 => x"0cfb3d0d",
          4283 => x"800b82d8",
          4284 => x"d408fc05",
          4285 => x"0c82d8d4",
          4286 => x"08880508",
          4287 => x"80259938",
          4288 => x"82d8d408",
          4289 => x"88050830",
          4290 => x"82d8d408",
          4291 => x"88050c81",
          4292 => x"0b82d8d4",
          4293 => x"08fc050c",
          4294 => x"82d8d408",
          4295 => x"8c050880",
          4296 => x"25903882",
          4297 => x"d8d4088c",
          4298 => x"05083082",
          4299 => x"d8d4088c",
          4300 => x"050c8153",
          4301 => x"82d8d408",
          4302 => x"8c050852",
          4303 => x"82d8d408",
          4304 => x"88050851",
          4305 => x"81a23f82",
          4306 => x"d8c80870",
          4307 => x"82d8d408",
          4308 => x"f8050c54",
          4309 => x"82d8d408",
          4310 => x"fc050880",
          4311 => x"2e903882",
          4312 => x"d8d408f8",
          4313 => x"05083082",
          4314 => x"d8d408f8",
          4315 => x"050c82d8",
          4316 => x"d408f805",
          4317 => x"087082d8",
          4318 => x"c80c5487",
          4319 => x"3d0d82d8",
          4320 => x"d40c0482",
          4321 => x"d8d40802",
          4322 => x"82d8d40c",
          4323 => x"fd3d0d80",
          4324 => x"5382d8d4",
          4325 => x"088c0508",
          4326 => x"5282d8d4",
          4327 => x"08880508",
          4328 => x"5180c53f",
          4329 => x"82d8c808",
          4330 => x"7082d8c8",
          4331 => x"0c54853d",
          4332 => x"0d82d8d4",
          4333 => x"0c0482d8",
          4334 => x"d4080282",
          4335 => x"d8d40cfd",
          4336 => x"3d0d8153",
          4337 => x"82d8d408",
          4338 => x"8c050852",
          4339 => x"82d8d408",
          4340 => x"88050851",
          4341 => x"933f82d8",
          4342 => x"c8087082",
          4343 => x"d8c80c54",
          4344 => x"853d0d82",
          4345 => x"d8d40c04",
          4346 => x"82d8d408",
          4347 => x"0282d8d4",
          4348 => x"0cfd3d0d",
          4349 => x"810b82d8",
          4350 => x"d408fc05",
          4351 => x"0c800b82",
          4352 => x"d8d408f8",
          4353 => x"050c82d8",
          4354 => x"d4088c05",
          4355 => x"0882d8d4",
          4356 => x"08880508",
          4357 => x"27b93882",
          4358 => x"d8d408fc",
          4359 => x"0508802e",
          4360 => x"ae38800b",
          4361 => x"82d8d408",
          4362 => x"8c050824",
          4363 => x"a23882d8",
          4364 => x"d4088c05",
          4365 => x"081082d8",
          4366 => x"d4088c05",
          4367 => x"0c82d8d4",
          4368 => x"08fc0508",
          4369 => x"1082d8d4",
          4370 => x"08fc050c",
          4371 => x"ffb83982",
          4372 => x"d8d408fc",
          4373 => x"0508802e",
          4374 => x"80e13882",
          4375 => x"d8d4088c",
          4376 => x"050882d8",
          4377 => x"d4088805",
          4378 => x"0826ad38",
          4379 => x"82d8d408",
          4380 => x"88050882",
          4381 => x"d8d4088c",
          4382 => x"05083182",
          4383 => x"d8d40888",
          4384 => x"050c82d8",
          4385 => x"d408f805",
          4386 => x"0882d8d4",
          4387 => x"08fc0508",
          4388 => x"0782d8d4",
          4389 => x"08f8050c",
          4390 => x"82d8d408",
          4391 => x"fc050881",
          4392 => x"2a82d8d4",
          4393 => x"08fc050c",
          4394 => x"82d8d408",
          4395 => x"8c050881",
          4396 => x"2a82d8d4",
          4397 => x"088c050c",
          4398 => x"ff953982",
          4399 => x"d8d40890",
          4400 => x"0508802e",
          4401 => x"933882d8",
          4402 => x"d4088805",
          4403 => x"087082d8",
          4404 => x"d408f405",
          4405 => x"0c519139",
          4406 => x"82d8d408",
          4407 => x"f8050870",
          4408 => x"82d8d408",
          4409 => x"f4050c51",
          4410 => x"82d8d408",
          4411 => x"f4050882",
          4412 => x"d8c80c85",
          4413 => x"3d0d82d8",
          4414 => x"d40c0482",
          4415 => x"d8d40802",
          4416 => x"82d8d40c",
          4417 => x"f73d0d80",
          4418 => x"0b82d8d4",
          4419 => x"08f00534",
          4420 => x"82d8d408",
          4421 => x"8c050853",
          4422 => x"80730c82",
          4423 => x"d8d40888",
          4424 => x"05087008",
          4425 => x"51537233",
          4426 => x"537282d8",
          4427 => x"d408f805",
          4428 => x"347281ff",
          4429 => x"065372a0",
          4430 => x"2e098106",
          4431 => x"913882d8",
          4432 => x"d4088805",
          4433 => x"08700881",
          4434 => x"05710c53",
          4435 => x"ce3982d8",
          4436 => x"d408f805",
          4437 => x"335372ad",
          4438 => x"2e098106",
          4439 => x"a438810b",
          4440 => x"82d8d408",
          4441 => x"f0053482",
          4442 => x"d8d40888",
          4443 => x"05087008",
          4444 => x"8105710c",
          4445 => x"70085153",
          4446 => x"723382d8",
          4447 => x"d408f805",
          4448 => x"3482d8d4",
          4449 => x"08f80533",
          4450 => x"5372b02e",
          4451 => x"09810681",
          4452 => x"dc3882d8",
          4453 => x"d4088805",
          4454 => x"08700881",
          4455 => x"05710c70",
          4456 => x"08515372",
          4457 => x"3382d8d4",
          4458 => x"08f80534",
          4459 => x"82d8d408",
          4460 => x"f8053382",
          4461 => x"d8d408e8",
          4462 => x"050c82d8",
          4463 => x"d408e805",
          4464 => x"0880e22e",
          4465 => x"b63882d8",
          4466 => x"d408e805",
          4467 => x"0880f82e",
          4468 => x"843880cd",
          4469 => x"39900b82",
          4470 => x"d8d408f4",
          4471 => x"053482d8",
          4472 => x"d4088805",
          4473 => x"08700881",
          4474 => x"05710c70",
          4475 => x"08515372",
          4476 => x"3382d8d4",
          4477 => x"08f80534",
          4478 => x"81a43982",
          4479 => x"0b82d8d4",
          4480 => x"08f40534",
          4481 => x"82d8d408",
          4482 => x"88050870",
          4483 => x"08810571",
          4484 => x"0c700851",
          4485 => x"53723382",
          4486 => x"d8d408f8",
          4487 => x"053480fe",
          4488 => x"3982d8d4",
          4489 => x"08f80533",
          4490 => x"5372a026",
          4491 => x"8d38810b",
          4492 => x"82d8d408",
          4493 => x"ec050c83",
          4494 => x"803982d8",
          4495 => x"d408f805",
          4496 => x"3353af73",
          4497 => x"27903882",
          4498 => x"d8d408f8",
          4499 => x"05335372",
          4500 => x"b9268338",
          4501 => x"8d39800b",
          4502 => x"82d8d408",
          4503 => x"ec050c82",
          4504 => x"d839880b",
          4505 => x"82d8d408",
          4506 => x"f40534b2",
          4507 => x"3982d8d4",
          4508 => x"08f80533",
          4509 => x"53af7327",
          4510 => x"903882d8",
          4511 => x"d408f805",
          4512 => x"335372b9",
          4513 => x"2683388d",
          4514 => x"39800b82",
          4515 => x"d8d408ec",
          4516 => x"050c82a5",
          4517 => x"398a0b82",
          4518 => x"d8d408f4",
          4519 => x"0534800b",
          4520 => x"82d8d408",
          4521 => x"fc050c82",
          4522 => x"d8d408f8",
          4523 => x"053353a0",
          4524 => x"732781cf",
          4525 => x"3882d8d4",
          4526 => x"08f80533",
          4527 => x"5380e073",
          4528 => x"27943882",
          4529 => x"d8d408f8",
          4530 => x"0533e011",
          4531 => x"51537282",
          4532 => x"d8d408f8",
          4533 => x"053482d8",
          4534 => x"d408f805",
          4535 => x"33d01151",
          4536 => x"537282d8",
          4537 => x"d408f805",
          4538 => x"3482d8d4",
          4539 => x"08f80533",
          4540 => x"53907327",
          4541 => x"ad3882d8",
          4542 => x"d408f805",
          4543 => x"33f91151",
          4544 => x"537282d8",
          4545 => x"d408f805",
          4546 => x"3482d8d4",
          4547 => x"08f80533",
          4548 => x"53728926",
          4549 => x"8d38800b",
          4550 => x"82d8d408",
          4551 => x"ec050c81",
          4552 => x"983982d8",
          4553 => x"d408f805",
          4554 => x"3382d8d4",
          4555 => x"08f40533",
          4556 => x"54547274",
          4557 => x"268d3880",
          4558 => x"0b82d8d4",
          4559 => x"08ec050c",
          4560 => x"80f73982",
          4561 => x"d8d408f4",
          4562 => x"05337082",
          4563 => x"d8d408fc",
          4564 => x"05082982",
          4565 => x"d8d408f8",
          4566 => x"05337012",
          4567 => x"82d8d408",
          4568 => x"fc050c82",
          4569 => x"d8d40888",
          4570 => x"05087008",
          4571 => x"8105710c",
          4572 => x"70085151",
          4573 => x"52555372",
          4574 => x"3382d8d4",
          4575 => x"08f80534",
          4576 => x"fea53982",
          4577 => x"d8d408f0",
          4578 => x"05335372",
          4579 => x"802e9038",
          4580 => x"82d8d408",
          4581 => x"fc050830",
          4582 => x"82d8d408",
          4583 => x"fc050c82",
          4584 => x"d8d4088c",
          4585 => x"050882d8",
          4586 => x"d408fc05",
          4587 => x"08710c53",
          4588 => x"810b82d8",
          4589 => x"d408ec05",
          4590 => x"0c82d8d4",
          4591 => x"08ec0508",
          4592 => x"82d8c80c",
          4593 => x"8b3d0d82",
          4594 => x"d8d40c04",
          4595 => x"82d8d408",
          4596 => x"0282d8d4",
          4597 => x"0cf73d0d",
          4598 => x"800b82d8",
          4599 => x"d408f005",
          4600 => x"3482d8d4",
          4601 => x"088c0508",
          4602 => x"5380730c",
          4603 => x"82d8d408",
          4604 => x"88050870",
          4605 => x"08515372",
          4606 => x"33537282",
          4607 => x"d8d408f8",
          4608 => x"05347281",
          4609 => x"ff065372",
          4610 => x"a02e0981",
          4611 => x"06913882",
          4612 => x"d8d40888",
          4613 => x"05087008",
          4614 => x"8105710c",
          4615 => x"53ce3982",
          4616 => x"d8d408f8",
          4617 => x"05335372",
          4618 => x"ad2e0981",
          4619 => x"06a43881",
          4620 => x"0b82d8d4",
          4621 => x"08f00534",
          4622 => x"82d8d408",
          4623 => x"88050870",
          4624 => x"08810571",
          4625 => x"0c700851",
          4626 => x"53723382",
          4627 => x"d8d408f8",
          4628 => x"053482d8",
          4629 => x"d408f805",
          4630 => x"335372b0",
          4631 => x"2e098106",
          4632 => x"81dc3882",
          4633 => x"d8d40888",
          4634 => x"05087008",
          4635 => x"8105710c",
          4636 => x"70085153",
          4637 => x"723382d8",
          4638 => x"d408f805",
          4639 => x"3482d8d4",
          4640 => x"08f80533",
          4641 => x"82d8d408",
          4642 => x"e8050c82",
          4643 => x"d8d408e8",
          4644 => x"050880e2",
          4645 => x"2eb63882",
          4646 => x"d8d408e8",
          4647 => x"050880f8",
          4648 => x"2e843880",
          4649 => x"cd39900b",
          4650 => x"82d8d408",
          4651 => x"f4053482",
          4652 => x"d8d40888",
          4653 => x"05087008",
          4654 => x"8105710c",
          4655 => x"70085153",
          4656 => x"723382d8",
          4657 => x"d408f805",
          4658 => x"3481a439",
          4659 => x"820b82d8",
          4660 => x"d408f405",
          4661 => x"3482d8d4",
          4662 => x"08880508",
          4663 => x"70088105",
          4664 => x"710c7008",
          4665 => x"51537233",
          4666 => x"82d8d408",
          4667 => x"f8053480",
          4668 => x"fe3982d8",
          4669 => x"d408f805",
          4670 => x"335372a0",
          4671 => x"268d3881",
          4672 => x"0b82d8d4",
          4673 => x"08ec050c",
          4674 => x"83803982",
          4675 => x"d8d408f8",
          4676 => x"053353af",
          4677 => x"73279038",
          4678 => x"82d8d408",
          4679 => x"f8053353",
          4680 => x"72b92683",
          4681 => x"388d3980",
          4682 => x"0b82d8d4",
          4683 => x"08ec050c",
          4684 => x"82d83988",
          4685 => x"0b82d8d4",
          4686 => x"08f40534",
          4687 => x"b23982d8",
          4688 => x"d408f805",
          4689 => x"3353af73",
          4690 => x"27903882",
          4691 => x"d8d408f8",
          4692 => x"05335372",
          4693 => x"b9268338",
          4694 => x"8d39800b",
          4695 => x"82d8d408",
          4696 => x"ec050c82",
          4697 => x"a5398a0b",
          4698 => x"82d8d408",
          4699 => x"f4053480",
          4700 => x"0b82d8d4",
          4701 => x"08fc050c",
          4702 => x"82d8d408",
          4703 => x"f8053353",
          4704 => x"a0732781",
          4705 => x"cf3882d8",
          4706 => x"d408f805",
          4707 => x"335380e0",
          4708 => x"73279438",
          4709 => x"82d8d408",
          4710 => x"f80533e0",
          4711 => x"11515372",
          4712 => x"82d8d408",
          4713 => x"f8053482",
          4714 => x"d8d408f8",
          4715 => x"0533d011",
          4716 => x"51537282",
          4717 => x"d8d408f8",
          4718 => x"053482d8",
          4719 => x"d408f805",
          4720 => x"33539073",
          4721 => x"27ad3882",
          4722 => x"d8d408f8",
          4723 => x"0533f911",
          4724 => x"51537282",
          4725 => x"d8d408f8",
          4726 => x"053482d8",
          4727 => x"d408f805",
          4728 => x"33537289",
          4729 => x"268d3880",
          4730 => x"0b82d8d4",
          4731 => x"08ec050c",
          4732 => x"81983982",
          4733 => x"d8d408f8",
          4734 => x"053382d8",
          4735 => x"d408f405",
          4736 => x"33545472",
          4737 => x"74268d38",
          4738 => x"800b82d8",
          4739 => x"d408ec05",
          4740 => x"0c80f739",
          4741 => x"82d8d408",
          4742 => x"f4053370",
          4743 => x"82d8d408",
          4744 => x"fc050829",
          4745 => x"82d8d408",
          4746 => x"f8053370",
          4747 => x"1282d8d4",
          4748 => x"08fc050c",
          4749 => x"82d8d408",
          4750 => x"88050870",
          4751 => x"08810571",
          4752 => x"0c700851",
          4753 => x"51525553",
          4754 => x"723382d8",
          4755 => x"d408f805",
          4756 => x"34fea539",
          4757 => x"82d8d408",
          4758 => x"f0053353",
          4759 => x"72802e90",
          4760 => x"3882d8d4",
          4761 => x"08fc0508",
          4762 => x"3082d8d4",
          4763 => x"08fc050c",
          4764 => x"82d8d408",
          4765 => x"8c050882",
          4766 => x"d8d408fc",
          4767 => x"0508710c",
          4768 => x"53810b82",
          4769 => x"d8d408ec",
          4770 => x"050c82d8",
          4771 => x"d408ec05",
          4772 => x"0882d8c8",
          4773 => x"0c8b3d0d",
          4774 => x"82d8d40c",
          4775 => x"04f93d0d",
          4776 => x"79700870",
          4777 => x"56565874",
          4778 => x"802e80e3",
          4779 => x"38953975",
          4780 => x"0851e6d1",
          4781 => x"3f82d8c8",
          4782 => x"0815780c",
          4783 => x"85163354",
          4784 => x"80cd3974",
          4785 => x"335473a0",
          4786 => x"2e098106",
          4787 => x"86388115",
          4788 => x"55f13980",
          4789 => x"57769029",
          4790 => x"82d3c805",
          4791 => x"70085256",
          4792 => x"e6a33f82",
          4793 => x"d8c80853",
          4794 => x"74527508",
          4795 => x"51e9a33f",
          4796 => x"82d8c808",
          4797 => x"8b388416",
          4798 => x"33547381",
          4799 => x"2effb038",
          4800 => x"81177081",
          4801 => x"ff065854",
          4802 => x"997727c9",
          4803 => x"38ff5473",
          4804 => x"82d8c80c",
          4805 => x"893d0d04",
          4806 => x"ff3d0d73",
          4807 => x"52719326",
          4808 => x"818e3871",
          4809 => x"842982ae",
          4810 => x"f4055271",
          4811 => x"080482b4",
          4812 => x"e4518180",
          4813 => x"3982b4f0",
          4814 => x"5180f939",
          4815 => x"82b58051",
          4816 => x"80f23982",
          4817 => x"b5905180",
          4818 => x"eb3982b5",
          4819 => x"a05180e4",
          4820 => x"3982b5b0",
          4821 => x"5180dd39",
          4822 => x"82b5c451",
          4823 => x"80d63982",
          4824 => x"b5d45180",
          4825 => x"cf3982b5",
          4826 => x"ec5180c8",
          4827 => x"3982b684",
          4828 => x"5180c139",
          4829 => x"82b69c51",
          4830 => x"bb3982b6",
          4831 => x"b851b539",
          4832 => x"82b6cc51",
          4833 => x"af3982b6",
          4834 => x"f451a939",
          4835 => x"82b78451",
          4836 => x"a33982b7",
          4837 => x"a4519d39",
          4838 => x"82b7b451",
          4839 => x"973982b7",
          4840 => x"cc519139",
          4841 => x"82b7e451",
          4842 => x"8b3982b7",
          4843 => x"fc518539",
          4844 => x"82b88851",
          4845 => x"d8ad3f83",
          4846 => x"3d0d04fb",
          4847 => x"3d0d7779",
          4848 => x"56567487",
          4849 => x"e7268a38",
          4850 => x"74527587",
          4851 => x"e8295190",
          4852 => x"3987e852",
          4853 => x"7451efab",
          4854 => x"3f82d8c8",
          4855 => x"08527551",
          4856 => x"efa13f82",
          4857 => x"d8c80854",
          4858 => x"79537552",
          4859 => x"82b89851",
          4860 => x"ffbbe53f",
          4861 => x"873d0d04",
          4862 => x"ec3d0d66",
          4863 => x"02840580",
          4864 => x"e305335b",
          4865 => x"57806878",
          4866 => x"30707a07",
          4867 => x"73255157",
          4868 => x"59597856",
          4869 => x"7787ff26",
          4870 => x"83388156",
          4871 => x"74760770",
          4872 => x"81ff0651",
          4873 => x"55935674",
          4874 => x"81823881",
          4875 => x"5376528c",
          4876 => x"3d705256",
          4877 => x"8196903f",
          4878 => x"82d8c808",
          4879 => x"5782d8c8",
          4880 => x"08b93882",
          4881 => x"d8c80887",
          4882 => x"c098880c",
          4883 => x"82d8c808",
          4884 => x"59963dd4",
          4885 => x"05548480",
          4886 => x"53775275",
          4887 => x"51819acc",
          4888 => x"3f82d8c8",
          4889 => x"085782d8",
          4890 => x"c8089038",
          4891 => x"7a557480",
          4892 => x"2e893874",
          4893 => x"19751959",
          4894 => x"59d73996",
          4895 => x"3dd80551",
          4896 => x"81a2c33f",
          4897 => x"76307078",
          4898 => x"0780257b",
          4899 => x"30709f2a",
          4900 => x"72065157",
          4901 => x"51567480",
          4902 => x"2e903882",
          4903 => x"b8bc5387",
          4904 => x"c0988808",
          4905 => x"527851fe",
          4906 => x"923f7656",
          4907 => x"7582d8c8",
          4908 => x"0c963d0d",
          4909 => x"04f73d0d",
          4910 => x"7d028405",
          4911 => x"bb053359",
          4912 => x"5aff5980",
          4913 => x"537c527b",
          4914 => x"51fead3f",
          4915 => x"82d8c808",
          4916 => x"80cb3877",
          4917 => x"802e8838",
          4918 => x"77812ebf",
          4919 => x"38bf3982",
          4920 => x"f4a85782",
          4921 => x"f4a85682",
          4922 => x"f4a85582",
          4923 => x"f4b00854",
          4924 => x"82f4ac08",
          4925 => x"5382f4a8",
          4926 => x"085282b8",
          4927 => x"c451ffb9",
          4928 => x"d73f82f4",
          4929 => x"a8566255",
          4930 => x"615482d8",
          4931 => x"c8536052",
          4932 => x"7f51792d",
          4933 => x"82d8c808",
          4934 => x"59833979",
          4935 => x"047882d8",
          4936 => x"c80c8b3d",
          4937 => x"0d04f33d",
          4938 => x"0d7f6163",
          4939 => x"028c0580",
          4940 => x"cf053373",
          4941 => x"73156841",
          4942 => x"5f5c5c5e",
          4943 => x"5e5e7a52",
          4944 => x"82b8f851",
          4945 => x"ffb9913f",
          4946 => x"82b98051",
          4947 => x"ffb9893f",
          4948 => x"80557479",
          4949 => x"27818038",
          4950 => x"7b902e89",
          4951 => x"387ba02e",
          4952 => x"a73880c6",
          4953 => x"39741853",
          4954 => x"727a278e",
          4955 => x"38722252",
          4956 => x"82b98451",
          4957 => x"ffb8e13f",
          4958 => x"893982b9",
          4959 => x"9051ffb8",
          4960 => x"d73f8215",
          4961 => x"5580c339",
          4962 => x"74185372",
          4963 => x"7a278e38",
          4964 => x"72085282",
          4965 => x"b8f851ff",
          4966 => x"b8be3f89",
          4967 => x"3982b98c",
          4968 => x"51ffb8b4",
          4969 => x"3f841555",
          4970 => x"a1397418",
          4971 => x"53727a27",
          4972 => x"8e387233",
          4973 => x"5282b998",
          4974 => x"51ffb89c",
          4975 => x"3f893982",
          4976 => x"b9a051ff",
          4977 => x"b8923f81",
          4978 => x"155582f4",
          4979 => x"ac0852a0",
          4980 => x"51d7df3f",
          4981 => x"fefc3982",
          4982 => x"b9a451ff",
          4983 => x"b7fa3f80",
          4984 => x"55747927",
          4985 => x"80c63874",
          4986 => x"18703355",
          4987 => x"53805672",
          4988 => x"7a278338",
          4989 => x"81568053",
          4990 => x"9f742783",
          4991 => x"38815375",
          4992 => x"73067081",
          4993 => x"ff065153",
          4994 => x"72802e90",
          4995 => x"387380fe",
          4996 => x"268a3882",
          4997 => x"f4ac0852",
          4998 => x"73518839",
          4999 => x"82f4ac08",
          5000 => x"52a051d7",
          5001 => x"8d3f8115",
          5002 => x"55ffb639",
          5003 => x"82b9a851",
          5004 => x"d3b13f78",
          5005 => x"18791c5c",
          5006 => x"58a1803f",
          5007 => x"82d8c808",
          5008 => x"982b7098",
          5009 => x"2c515776",
          5010 => x"a02e0981",
          5011 => x"06aa38a0",
          5012 => x"ea3f82d8",
          5013 => x"c808982b",
          5014 => x"70982c70",
          5015 => x"a0327030",
          5016 => x"729b3270",
          5017 => x"30707207",
          5018 => x"73750706",
          5019 => x"51585859",
          5020 => x"57515780",
          5021 => x"7324d838",
          5022 => x"769b2e09",
          5023 => x"81068538",
          5024 => x"80538c39",
          5025 => x"7c1e5372",
          5026 => x"7826fdb2",
          5027 => x"38ff5372",
          5028 => x"82d8c80c",
          5029 => x"8f3d0d04",
          5030 => x"fc3d0d02",
          5031 => x"9b053382",
          5032 => x"b9ac5382",
          5033 => x"b9b45255",
          5034 => x"ffb6ad3f",
          5035 => x"82d7a022",
          5036 => x"51a9d93f",
          5037 => x"82b9c054",
          5038 => x"82b9cc53",
          5039 => x"82d7a133",
          5040 => x"5282b9d4",
          5041 => x"51ffb690",
          5042 => x"3f74802e",
          5043 => x"8438a58d",
          5044 => x"3f863d0d",
          5045 => x"04fe3d0d",
          5046 => x"87c09680",
          5047 => x"0853aab6",
          5048 => x"3f81519c",
          5049 => x"c33f82b9",
          5050 => x"f0519dd8",
          5051 => x"3f80519c",
          5052 => x"b73f7281",
          5053 => x"2a708106",
          5054 => x"51527180",
          5055 => x"2e923881",
          5056 => x"519ca53f",
          5057 => x"82ba8851",
          5058 => x"9dba3f80",
          5059 => x"519c993f",
          5060 => x"72822a70",
          5061 => x"81065152",
          5062 => x"71802e92",
          5063 => x"3881519c",
          5064 => x"873f82ba",
          5065 => x"98519d9c",
          5066 => x"3f80519b",
          5067 => x"fb3f7283",
          5068 => x"2a708106",
          5069 => x"51527180",
          5070 => x"2e923881",
          5071 => x"519be93f",
          5072 => x"82baa851",
          5073 => x"9cfe3f80",
          5074 => x"519bdd3f",
          5075 => x"72842a70",
          5076 => x"81065152",
          5077 => x"71802e92",
          5078 => x"3881519b",
          5079 => x"cb3f82ba",
          5080 => x"bc519ce0",
          5081 => x"3f80519b",
          5082 => x"bf3f7285",
          5083 => x"2a708106",
          5084 => x"51527180",
          5085 => x"2e923881",
          5086 => x"519bad3f",
          5087 => x"82bad051",
          5088 => x"9cc23f80",
          5089 => x"519ba13f",
          5090 => x"72862a70",
          5091 => x"81065152",
          5092 => x"71802e92",
          5093 => x"3881519b",
          5094 => x"8f3f82ba",
          5095 => x"e4519ca4",
          5096 => x"3f80519b",
          5097 => x"833f7287",
          5098 => x"2a708106",
          5099 => x"51527180",
          5100 => x"2e923881",
          5101 => x"519af13f",
          5102 => x"82baf851",
          5103 => x"9c863f80",
          5104 => x"519ae53f",
          5105 => x"72882a70",
          5106 => x"81065152",
          5107 => x"71802e92",
          5108 => x"3881519a",
          5109 => x"d33f82bb",
          5110 => x"8c519be8",
          5111 => x"3f80519a",
          5112 => x"c73fa8ba",
          5113 => x"3f843d0d",
          5114 => x"04fb3d0d",
          5115 => x"77028405",
          5116 => x"a3053370",
          5117 => x"55565680",
          5118 => x"527551e2",
          5119 => x"e93f0b0b",
          5120 => x"82d3c433",
          5121 => x"5473a938",
          5122 => x"815382bb",
          5123 => x"c85282ef",
          5124 => x"d851818e",
          5125 => x"b23f82d8",
          5126 => x"c8083070",
          5127 => x"82d8c808",
          5128 => x"07802582",
          5129 => x"71315151",
          5130 => x"54730b0b",
          5131 => x"82d3c434",
          5132 => x"0b0b82d3",
          5133 => x"c4335473",
          5134 => x"812e0981",
          5135 => x"06af3882",
          5136 => x"efd85374",
          5137 => x"52755181",
          5138 => x"c9823f82",
          5139 => x"d8c80880",
          5140 => x"2e8b3882",
          5141 => x"d8c80851",
          5142 => x"cf893f91",
          5143 => x"3982efd8",
          5144 => x"51819ae2",
          5145 => x"3f820b0b",
          5146 => x"0b82d3c4",
          5147 => x"340b0b82",
          5148 => x"d3c43354",
          5149 => x"73822e09",
          5150 => x"81068c38",
          5151 => x"82bbd853",
          5152 => x"74527551",
          5153 => x"aeb23f80",
          5154 => x"0b82d8c8",
          5155 => x"0c873d0d",
          5156 => x"04ce3d0d",
          5157 => x"80707182",
          5158 => x"efd40c5f",
          5159 => x"5d81527c",
          5160 => x"5180cbcb",
          5161 => x"3f82d8c8",
          5162 => x"0881ff06",
          5163 => x"59787d2e",
          5164 => x"098106a3",
          5165 => x"38963d59",
          5166 => x"835382bb",
          5167 => x"e4527851",
          5168 => x"dca33f7c",
          5169 => x"53785282",
          5170 => x"d9f45181",
          5171 => x"8c983f82",
          5172 => x"d8c8087d",
          5173 => x"2e883882",
          5174 => x"bbe85191",
          5175 => x"d7398170",
          5176 => x"5f5d82bc",
          5177 => x"a051ffb1",
          5178 => x"ef3f963d",
          5179 => x"70465a80",
          5180 => x"f8527951",
          5181 => x"fdf33fb4",
          5182 => x"3dff8405",
          5183 => x"51f39e3f",
          5184 => x"82d8c808",
          5185 => x"902b7090",
          5186 => x"2c515978",
          5187 => x"80c12e89",
          5188 => x"d4387880",
          5189 => x"c12480d9",
          5190 => x"3878ab2e",
          5191 => x"83b93878",
          5192 => x"ab24a438",
          5193 => x"78822e81",
          5194 => x"b3387882",
          5195 => x"248a3878",
          5196 => x"802effae",
          5197 => x"388f8239",
          5198 => x"78842e82",
          5199 => x"83387894",
          5200 => x"2e82ad38",
          5201 => x"8ef33978",
          5202 => x"bd2e84fc",
          5203 => x"3878bd24",
          5204 => x"903878b0",
          5205 => x"2e83a638",
          5206 => x"78bc2e84",
          5207 => x"84388ed9",
          5208 => x"3978bf2e",
          5209 => x"85c43878",
          5210 => x"80c02e86",
          5211 => x"bd388ec9",
          5212 => x"397880d5",
          5213 => x"2e8da238",
          5214 => x"7880d524",
          5215 => x"b0387880",
          5216 => x"d02e8cd9",
          5217 => x"387880d0",
          5218 => x"24923878",
          5219 => x"80c22e89",
          5220 => x"fc387880",
          5221 => x"c32e8ba5",
          5222 => x"388e9e39",
          5223 => x"7880d12e",
          5224 => x"8cca3878",
          5225 => x"80d42e8c",
          5226 => x"d3388e8d",
          5227 => x"39788182",
          5228 => x"2e8de438",
          5229 => x"78818224",
          5230 => x"92387880",
          5231 => x"f82e8cf6",
          5232 => x"387880f9",
          5233 => x"2e8d9338",
          5234 => x"8def3978",
          5235 => x"81832e8d",
          5236 => x"d5387881",
          5237 => x"852e8ddb",
          5238 => x"388dde39",
          5239 => x"b43dff80",
          5240 => x"1153ff84",
          5241 => x"0551ebe4",
          5242 => x"3f82d8c8",
          5243 => x"08883882",
          5244 => x"bca4518f",
          5245 => x"bf39b43d",
          5246 => x"fefc1153",
          5247 => x"ff840551",
          5248 => x"ebca3f82",
          5249 => x"d8c80880",
          5250 => x"2e883881",
          5251 => x"63258338",
          5252 => x"80430280",
          5253 => x"cb053352",
          5254 => x"0280cf05",
          5255 => x"335180c8",
          5256 => x"ce3f82d8",
          5257 => x"c80881ff",
          5258 => x"0659788d",
          5259 => x"3882bcb4",
          5260 => x"51cbb03f",
          5261 => x"815efdaa",
          5262 => x"3982bcc4",
          5263 => x"518ef539",
          5264 => x"b43dff80",
          5265 => x"1153ff84",
          5266 => x"0551eb80",
          5267 => x"3f82d8c8",
          5268 => x"08802efd",
          5269 => x"8d388053",
          5270 => x"80520280",
          5271 => x"cf053351",
          5272 => x"80ccd93f",
          5273 => x"82d8c808",
          5274 => x"5282bcdc",
          5275 => x"518ca139",
          5276 => x"b43dff80",
          5277 => x"1153ff84",
          5278 => x"0551ead0",
          5279 => x"3f82d8c8",
          5280 => x"08802e87",
          5281 => x"38638926",
          5282 => x"fcd838b4",
          5283 => x"3dfefc11",
          5284 => x"53ff8405",
          5285 => x"51eab53f",
          5286 => x"82d8c808",
          5287 => x"863882d8",
          5288 => x"c8084363",
          5289 => x"5382bce4",
          5290 => x"527951ff",
          5291 => x"b1923f02",
          5292 => x"80cb0533",
          5293 => x"53795263",
          5294 => x"84b82982",
          5295 => x"d9f40551",
          5296 => x"8188a33f",
          5297 => x"82d8c808",
          5298 => x"818c3882",
          5299 => x"bcb451ca",
          5300 => x"923f815d",
          5301 => x"fc8c39b4",
          5302 => x"3dff8405",
          5303 => x"518fc23f",
          5304 => x"82d8c808",
          5305 => x"b53dff84",
          5306 => x"05525b90",
          5307 => x"d83f8153",
          5308 => x"82d8c808",
          5309 => x"527a51f1",
          5310 => x"ff3f80d1",
          5311 => x"39b43dff",
          5312 => x"8405518f",
          5313 => x"9c3f82d8",
          5314 => x"c808b53d",
          5315 => x"ff840552",
          5316 => x"5b90b23f",
          5317 => x"82d8c808",
          5318 => x"b53dff84",
          5319 => x"05525a90",
          5320 => x"a43f82d8",
          5321 => x"c808b53d",
          5322 => x"ff840552",
          5323 => x"5990963f",
          5324 => x"82d6ec58",
          5325 => x"82d8f857",
          5326 => x"80568055",
          5327 => x"82d8c808",
          5328 => x"81ff0654",
          5329 => x"78537952",
          5330 => x"7a51f2e9",
          5331 => x"3f82d8c8",
          5332 => x"08802efb",
          5333 => x"8d3882d8",
          5334 => x"c80851ef",
          5335 => x"bb3ffb82",
          5336 => x"39b43dff",
          5337 => x"801153ff",
          5338 => x"840551e8",
          5339 => x"df3f82d8",
          5340 => x"c808802e",
          5341 => x"faec38b4",
          5342 => x"3dfefc11",
          5343 => x"53ff8405",
          5344 => x"51e8c93f",
          5345 => x"82d8c808",
          5346 => x"802efad6",
          5347 => x"38b43dfe",
          5348 => x"f81153ff",
          5349 => x"840551e8",
          5350 => x"b33f82d8",
          5351 => x"c8088638",
          5352 => x"82d8c808",
          5353 => x"4282bce8",
          5354 => x"51ffacac",
          5355 => x"3f63635c",
          5356 => x"5a797b27",
          5357 => x"81ec3861",
          5358 => x"59787a70",
          5359 => x"84055c0c",
          5360 => x"7a7a26f5",
          5361 => x"3881db39",
          5362 => x"b43dff80",
          5363 => x"1153ff84",
          5364 => x"0551e7f8",
          5365 => x"3f82d8c8",
          5366 => x"08802efa",
          5367 => x"8538b43d",
          5368 => x"fefc1153",
          5369 => x"ff840551",
          5370 => x"e7e23f82",
          5371 => x"d8c80880",
          5372 => x"2ef9ef38",
          5373 => x"b43dfef8",
          5374 => x"1153ff84",
          5375 => x"0551e7cc",
          5376 => x"3f82d8c8",
          5377 => x"08802ef9",
          5378 => x"d93882bc",
          5379 => x"f851ffab",
          5380 => x"c73f635a",
          5381 => x"79632781",
          5382 => x"89386159",
          5383 => x"79708105",
          5384 => x"5b337934",
          5385 => x"61810542",
          5386 => x"eb39b43d",
          5387 => x"ff801153",
          5388 => x"ff840551",
          5389 => x"e7963f82",
          5390 => x"d8c80880",
          5391 => x"2ef9a338",
          5392 => x"b43dfefc",
          5393 => x"1153ff84",
          5394 => x"0551e780",
          5395 => x"3f82d8c8",
          5396 => x"08802ef9",
          5397 => x"8d38b43d",
          5398 => x"fef81153",
          5399 => x"ff840551",
          5400 => x"e6ea3f82",
          5401 => x"d8c80880",
          5402 => x"2ef8f738",
          5403 => x"82bd8451",
          5404 => x"ffaae53f",
          5405 => x"635a7963",
          5406 => x"27a83861",
          5407 => x"70337b33",
          5408 => x"5e5a5b78",
          5409 => x"7c2e9238",
          5410 => x"78557a54",
          5411 => x"79335379",
          5412 => x"5282bd94",
          5413 => x"51ffaac0",
          5414 => x"3f811a62",
          5415 => x"8105435a",
          5416 => x"d5398a51",
          5417 => x"c9df3ff8",
          5418 => x"b939b43d",
          5419 => x"ff801153",
          5420 => x"ff840551",
          5421 => x"e6963f82",
          5422 => x"d8c80880",
          5423 => x"df3882d7",
          5424 => x"b4335978",
          5425 => x"802e8938",
          5426 => x"82d6ec08",
          5427 => x"4480cd39",
          5428 => x"82d7b533",
          5429 => x"5978802e",
          5430 => x"883882d6",
          5431 => x"f40844bc",
          5432 => x"3982d7b6",
          5433 => x"33597880",
          5434 => x"2e883882",
          5435 => x"d6fc0844",
          5436 => x"ab3982d7",
          5437 => x"b7335978",
          5438 => x"802e8838",
          5439 => x"82d78408",
          5440 => x"449a3982",
          5441 => x"d7b23359",
          5442 => x"78802e88",
          5443 => x"3882d78c",
          5444 => x"08448939",
          5445 => x"82d79c08",
          5446 => x"fc800544",
          5447 => x"b43dfefc",
          5448 => x"1153ff84",
          5449 => x"0551e5a4",
          5450 => x"3f82d8c8",
          5451 => x"0880de38",
          5452 => x"82d7b433",
          5453 => x"5978802e",
          5454 => x"893882d6",
          5455 => x"f0084380",
          5456 => x"cc3982d7",
          5457 => x"b5335978",
          5458 => x"802e8838",
          5459 => x"82d6f808",
          5460 => x"43bb3982",
          5461 => x"d7b63359",
          5462 => x"78802e88",
          5463 => x"3882d780",
          5464 => x"0843aa39",
          5465 => x"82d7b733",
          5466 => x"5978802e",
          5467 => x"883882d7",
          5468 => x"88084399",
          5469 => x"3982d7b2",
          5470 => x"33597880",
          5471 => x"2e883882",
          5472 => x"d7900843",
          5473 => x"883982d7",
          5474 => x"9c088805",
          5475 => x"43b43dfe",
          5476 => x"f81153ff",
          5477 => x"840551e4",
          5478 => x"b33f82d8",
          5479 => x"c808802e",
          5480 => x"a7388062",
          5481 => x"5c5c7a88",
          5482 => x"2e833881",
          5483 => x"5c7a9032",
          5484 => x"70307072",
          5485 => x"079f2a70",
          5486 => x"7f065151",
          5487 => x"5a5a7880",
          5488 => x"2e88387a",
          5489 => x"a02e8338",
          5490 => x"884282bd",
          5491 => x"b051c493",
          5492 => x"3fa05563",
          5493 => x"54615362",
          5494 => x"526351ee",
          5495 => x"c93f82bd",
          5496 => x"bc5187d0",
          5497 => x"39b43dff",
          5498 => x"801153ff",
          5499 => x"840551e3",
          5500 => x"db3f82d8",
          5501 => x"c808802e",
          5502 => x"f5e838b4",
          5503 => x"3dfefc11",
          5504 => x"53ff8405",
          5505 => x"51e3c53f",
          5506 => x"82d8c808",
          5507 => x"802ea438",
          5508 => x"63590280",
          5509 => x"cb053379",
          5510 => x"34638105",
          5511 => x"44b43dfe",
          5512 => x"fc1153ff",
          5513 => x"840551e3",
          5514 => x"a33f82d8",
          5515 => x"c808e138",
          5516 => x"f5b03963",
          5517 => x"70335452",
          5518 => x"82bdc851",
          5519 => x"ffa7993f",
          5520 => x"82f4a808",
          5521 => x"5380f852",
          5522 => x"7951ffa7",
          5523 => x"e03f7945",
          5524 => x"79335978",
          5525 => x"ae2ef58a",
          5526 => x"389f7927",
          5527 => x"9f38b43d",
          5528 => x"fefc1153",
          5529 => x"ff840551",
          5530 => x"e2e23f82",
          5531 => x"d8c80880",
          5532 => x"2e913863",
          5533 => x"590280cb",
          5534 => x"05337934",
          5535 => x"63810544",
          5536 => x"ffb13982",
          5537 => x"bdd451c2",
          5538 => x"da3fffa7",
          5539 => x"39b43dfe",
          5540 => x"f41153ff",
          5541 => x"840551dc",
          5542 => x"e23f82d8",
          5543 => x"c808802e",
          5544 => x"f4c038b4",
          5545 => x"3dfef011",
          5546 => x"53ff8405",
          5547 => x"51dccc3f",
          5548 => x"82d8c808",
          5549 => x"802ea538",
          5550 => x"605902be",
          5551 => x"05227970",
          5552 => x"82055b23",
          5553 => x"7841b43d",
          5554 => x"fef01153",
          5555 => x"ff840551",
          5556 => x"dca93f82",
          5557 => x"d8c808e0",
          5558 => x"38f48739",
          5559 => x"60702254",
          5560 => x"5282bdd8",
          5561 => x"51ffa5f0",
          5562 => x"3f82f4a8",
          5563 => x"085380f8",
          5564 => x"527951ff",
          5565 => x"a6b73f79",
          5566 => x"45793359",
          5567 => x"78ae2ef3",
          5568 => x"e138789f",
          5569 => x"26873860",
          5570 => x"820541d0",
          5571 => x"39b43dfe",
          5572 => x"f01153ff",
          5573 => x"840551db",
          5574 => x"e23f82d8",
          5575 => x"c808802e",
          5576 => x"92386059",
          5577 => x"02be0522",
          5578 => x"79708205",
          5579 => x"5b237841",
          5580 => x"ffaa3982",
          5581 => x"bdd451c1",
          5582 => x"aa3fffa0",
          5583 => x"39b43dfe",
          5584 => x"f41153ff",
          5585 => x"840551db",
          5586 => x"b23f82d8",
          5587 => x"c808802e",
          5588 => x"f39038b4",
          5589 => x"3dfef011",
          5590 => x"53ff8405",
          5591 => x"51db9c3f",
          5592 => x"82d8c808",
          5593 => x"802ea038",
          5594 => x"6060710c",
          5595 => x"59608405",
          5596 => x"41b43dfe",
          5597 => x"f01153ff",
          5598 => x"840551da",
          5599 => x"fe3f82d8",
          5600 => x"c808e538",
          5601 => x"f2dc3960",
          5602 => x"70085452",
          5603 => x"82bde451",
          5604 => x"ffa4c53f",
          5605 => x"82f4a808",
          5606 => x"5380f852",
          5607 => x"7951ffa5",
          5608 => x"8c3f7945",
          5609 => x"79335978",
          5610 => x"ae2ef2b6",
          5611 => x"389f7927",
          5612 => x"9b38b43d",
          5613 => x"fef01153",
          5614 => x"ff840551",
          5615 => x"dabd3f82",
          5616 => x"d8c80880",
          5617 => x"2e8d3860",
          5618 => x"60710c59",
          5619 => x"60840541",
          5620 => x"ffb53982",
          5621 => x"bdd451c0",
          5622 => x"8a3fffab",
          5623 => x"3982bdf4",
          5624 => x"51c0803f",
          5625 => x"82519889",
          5626 => x"3ff1f739",
          5627 => x"82be8c51",
          5628 => x"ffbff03f",
          5629 => x"a25197dd",
          5630 => x"3ff1e739",
          5631 => x"82bea051",
          5632 => x"ffbfe03f",
          5633 => x"8480810b",
          5634 => x"87c09484",
          5635 => x"0c848081",
          5636 => x"0b87c094",
          5637 => x"940cf1ca",
          5638 => x"3982beb4",
          5639 => x"51ffbfc3",
          5640 => x"3f8c8083",
          5641 => x"0b87c094",
          5642 => x"840c8c80",
          5643 => x"830b87c0",
          5644 => x"94940cf1",
          5645 => x"ad39b43d",
          5646 => x"ff801153",
          5647 => x"ff840551",
          5648 => x"df8a3f82",
          5649 => x"d8c80880",
          5650 => x"2ef19738",
          5651 => x"635282be",
          5652 => x"c851ffa3",
          5653 => x"833f6359",
          5654 => x"7804b43d",
          5655 => x"ff801153",
          5656 => x"ff840551",
          5657 => x"dee63f82",
          5658 => x"d8c80880",
          5659 => x"2ef0f338",
          5660 => x"635282be",
          5661 => x"e451ffa2",
          5662 => x"df3f6359",
          5663 => x"782d82d8",
          5664 => x"c808802e",
          5665 => x"f0dc3882",
          5666 => x"d8c80852",
          5667 => x"82bf8051",
          5668 => x"ffa2c53f",
          5669 => x"f0cc3982",
          5670 => x"bf9c51ff",
          5671 => x"bec53fff",
          5672 => x"a2973ff0",
          5673 => x"bd3982bf",
          5674 => x"b851ffbe",
          5675 => x"b63f8059",
          5676 => x"ffa63991",
          5677 => x"a83ff0aa",
          5678 => x"39794579",
          5679 => x"33597880",
          5680 => x"2ef09f38",
          5681 => x"7d7d0659",
          5682 => x"78802e81",
          5683 => x"cf38b43d",
          5684 => x"ff840551",
          5685 => x"83cb3f82",
          5686 => x"d8c8085b",
          5687 => x"815c7b82",
          5688 => x"2eb2387b",
          5689 => x"82248938",
          5690 => x"7b812e8c",
          5691 => x"3880ca39",
          5692 => x"7b832ead",
          5693 => x"3880c239",
          5694 => x"82bfcc56",
          5695 => x"7a5582bf",
          5696 => x"d0548053",
          5697 => x"82bfd452",
          5698 => x"b43dffb0",
          5699 => x"0551ffa4",
          5700 => x"af3fb839",
          5701 => x"7a52b43d",
          5702 => x"ffb00551",
          5703 => x"cad53fab",
          5704 => x"397a5582",
          5705 => x"bfd05480",
          5706 => x"5382bfe4",
          5707 => x"52b43dff",
          5708 => x"b00551ff",
          5709 => x"a48a3f93",
          5710 => x"397a5480",
          5711 => x"5382bff0",
          5712 => x"52b43dff",
          5713 => x"b00551ff",
          5714 => x"a3f63f82",
          5715 => x"d6ec5882",
          5716 => x"d8f85780",
          5717 => x"56645580",
          5718 => x"54848080",
          5719 => x"53848080",
          5720 => x"52b43dff",
          5721 => x"b00551e6",
          5722 => x"cc3f82d8",
          5723 => x"c80882d8",
          5724 => x"c8080970",
          5725 => x"30707207",
          5726 => x"8025515b",
          5727 => x"5b5f805a",
          5728 => x"7b832683",
          5729 => x"38815a78",
          5730 => x"7a065978",
          5731 => x"802e8d38",
          5732 => x"811c7081",
          5733 => x"ff065d59",
          5734 => x"7bfec338",
          5735 => x"7d81327d",
          5736 => x"81320759",
          5737 => x"788a387e",
          5738 => x"ff2e0981",
          5739 => x"06eeb338",
          5740 => x"82bff851",
          5741 => x"ffbcac3f",
          5742 => x"eea839f5",
          5743 => x"3d0d800b",
          5744 => x"82d8f834",
          5745 => x"87c0948c",
          5746 => x"70085455",
          5747 => x"87848052",
          5748 => x"7251d3af",
          5749 => x"3f82d8c8",
          5750 => x"08902b75",
          5751 => x"08555387",
          5752 => x"84805273",
          5753 => x"51d39c3f",
          5754 => x"7282d8c8",
          5755 => x"0807750c",
          5756 => x"87c0949c",
          5757 => x"70085455",
          5758 => x"87848052",
          5759 => x"7251d383",
          5760 => x"3f82d8c8",
          5761 => x"08902b75",
          5762 => x"08555387",
          5763 => x"84805273",
          5764 => x"51d2f03f",
          5765 => x"7282d8c8",
          5766 => x"0807750c",
          5767 => x"8c80830b",
          5768 => x"87c09484",
          5769 => x"0c8c8083",
          5770 => x"0b87c094",
          5771 => x"940c80fa",
          5772 => x"c05a80fd",
          5773 => x"ac5b8302",
          5774 => x"84059905",
          5775 => x"34805c82",
          5776 => x"f4a80b87",
          5777 => x"3d708813",
          5778 => x"0c70720c",
          5779 => x"82f4ac0c",
          5780 => x"5489be3f",
          5781 => x"93c03f82",
          5782 => x"c08851ff",
          5783 => x"bb853f82",
          5784 => x"c09451ff",
          5785 => x"bafd3f80",
          5786 => x"ddd55192",
          5787 => x"e33f8151",
          5788 => x"e8a63fec",
          5789 => x"9c3f8004",
          5790 => x"fe3d0d80",
          5791 => x"52835371",
          5792 => x"882b5287",
          5793 => x"d83f82d8",
          5794 => x"c80881ff",
          5795 => x"067207ff",
          5796 => x"14545272",
          5797 => x"8025e838",
          5798 => x"7182d8c8",
          5799 => x"0c843d0d",
          5800 => x"04fc3d0d",
          5801 => x"76700854",
          5802 => x"55807352",
          5803 => x"5472742e",
          5804 => x"818a3872",
          5805 => x"335170a0",
          5806 => x"2e098106",
          5807 => x"86388113",
          5808 => x"53f13972",
          5809 => x"335170a2",
          5810 => x"2e098106",
          5811 => x"86388113",
          5812 => x"53815472",
          5813 => x"5273812e",
          5814 => x"0981069f",
          5815 => x"38843981",
          5816 => x"12528072",
          5817 => x"33525470",
          5818 => x"a22e8338",
          5819 => x"81547080",
          5820 => x"2e9d3873",
          5821 => x"ea389839",
          5822 => x"81125280",
          5823 => x"72335254",
          5824 => x"70a02e83",
          5825 => x"38815470",
          5826 => x"802e8438",
          5827 => x"73ea3880",
          5828 => x"72335254",
          5829 => x"70a02e09",
          5830 => x"81068338",
          5831 => x"815470a2",
          5832 => x"32703070",
          5833 => x"80257607",
          5834 => x"51515170",
          5835 => x"802e8838",
          5836 => x"80727081",
          5837 => x"05543471",
          5838 => x"750c7251",
          5839 => x"7082d8c8",
          5840 => x"0c863d0d",
          5841 => x"04fc3d0d",
          5842 => x"76537208",
          5843 => x"802e9138",
          5844 => x"863dfc05",
          5845 => x"527251d3",
          5846 => x"a23f82d8",
          5847 => x"c8088538",
          5848 => x"80538339",
          5849 => x"74537282",
          5850 => x"d8c80c86",
          5851 => x"3d0d04fc",
          5852 => x"3d0d7682",
          5853 => x"1133ff05",
          5854 => x"52538152",
          5855 => x"708b2681",
          5856 => x"98388313",
          5857 => x"33ff0551",
          5858 => x"8252709e",
          5859 => x"26818a38",
          5860 => x"84133351",
          5861 => x"83527097",
          5862 => x"2680fe38",
          5863 => x"85133351",
          5864 => x"845270bb",
          5865 => x"2680f238",
          5866 => x"86133351",
          5867 => x"855270bb",
          5868 => x"2680e638",
          5869 => x"88132255",
          5870 => x"86527487",
          5871 => x"e72680d9",
          5872 => x"388a1322",
          5873 => x"54875273",
          5874 => x"87e72680",
          5875 => x"cc38810b",
          5876 => x"87c0989c",
          5877 => x"0c722287",
          5878 => x"c098bc0c",
          5879 => x"82133387",
          5880 => x"c098b80c",
          5881 => x"83133387",
          5882 => x"c098b40c",
          5883 => x"84133387",
          5884 => x"c098b00c",
          5885 => x"85133387",
          5886 => x"c098ac0c",
          5887 => x"86133387",
          5888 => x"c098a80c",
          5889 => x"7487c098",
          5890 => x"a40c7387",
          5891 => x"c098a00c",
          5892 => x"800b87c0",
          5893 => x"989c0c80",
          5894 => x"527182d8",
          5895 => x"c80c863d",
          5896 => x"0d04f33d",
          5897 => x"0d7f5b87",
          5898 => x"c0989c5d",
          5899 => x"817d0c87",
          5900 => x"c098bc08",
          5901 => x"5e7d7b23",
          5902 => x"87c098b8",
          5903 => x"085a7982",
          5904 => x"1c3487c0",
          5905 => x"98b4085a",
          5906 => x"79831c34",
          5907 => x"87c098b0",
          5908 => x"085a7984",
          5909 => x"1c3487c0",
          5910 => x"98ac085a",
          5911 => x"79851c34",
          5912 => x"87c098a8",
          5913 => x"085a7986",
          5914 => x"1c3487c0",
          5915 => x"98a4085c",
          5916 => x"7b881c23",
          5917 => x"87c098a0",
          5918 => x"085a798a",
          5919 => x"1c23807d",
          5920 => x"0c7983ff",
          5921 => x"ff06597b",
          5922 => x"83ffff06",
          5923 => x"58861b33",
          5924 => x"57851b33",
          5925 => x"56841b33",
          5926 => x"55831b33",
          5927 => x"54821b33",
          5928 => x"537d83ff",
          5929 => x"ff065282",
          5930 => x"c0ac51ff",
          5931 => x"9aaa3f8f",
          5932 => x"3d0d04fb",
          5933 => x"3d0d029f",
          5934 => x"053382d6",
          5935 => x"e8337081",
          5936 => x"ff065855",
          5937 => x"5587c094",
          5938 => x"84517580",
          5939 => x"2e863887",
          5940 => x"c0949451",
          5941 => x"70087096",
          5942 => x"2a708106",
          5943 => x"53545270",
          5944 => x"802e8c38",
          5945 => x"71912a70",
          5946 => x"81065151",
          5947 => x"70d73872",
          5948 => x"81327081",
          5949 => x"06515170",
          5950 => x"802e8d38",
          5951 => x"71932a70",
          5952 => x"81065151",
          5953 => x"70ffbe38",
          5954 => x"7381ff06",
          5955 => x"5187c094",
          5956 => x"80527080",
          5957 => x"2e863887",
          5958 => x"c0949052",
          5959 => x"74720c74",
          5960 => x"82d8c80c",
          5961 => x"873d0d04",
          5962 => x"ff3d0d02",
          5963 => x"8f053370",
          5964 => x"30709f2a",
          5965 => x"51525270",
          5966 => x"82d6e834",
          5967 => x"833d0d04",
          5968 => x"f93d0d02",
          5969 => x"a7053358",
          5970 => x"778a2e09",
          5971 => x"81068738",
          5972 => x"7a528d51",
          5973 => x"eb3f82d6",
          5974 => x"e8337081",
          5975 => x"ff065856",
          5976 => x"87c09484",
          5977 => x"5376802e",
          5978 => x"863887c0",
          5979 => x"94945372",
          5980 => x"0870962a",
          5981 => x"70810655",
          5982 => x"56547280",
          5983 => x"2e8c3873",
          5984 => x"912a7081",
          5985 => x"06515372",
          5986 => x"d7387481",
          5987 => x"32708106",
          5988 => x"51537280",
          5989 => x"2e8d3873",
          5990 => x"932a7081",
          5991 => x"06515372",
          5992 => x"ffbe3875",
          5993 => x"81ff0653",
          5994 => x"87c09480",
          5995 => x"5472802e",
          5996 => x"863887c0",
          5997 => x"94905477",
          5998 => x"740c800b",
          5999 => x"82d8c80c",
          6000 => x"893d0d04",
          6001 => x"f93d0d79",
          6002 => x"54807433",
          6003 => x"7081ff06",
          6004 => x"53535770",
          6005 => x"772e80fc",
          6006 => x"387181ff",
          6007 => x"06811582",
          6008 => x"d6e83370",
          6009 => x"81ff0659",
          6010 => x"57555887",
          6011 => x"c0948451",
          6012 => x"75802e86",
          6013 => x"3887c094",
          6014 => x"94517008",
          6015 => x"70962a70",
          6016 => x"81065354",
          6017 => x"5270802e",
          6018 => x"8c387191",
          6019 => x"2a708106",
          6020 => x"515170d7",
          6021 => x"38728132",
          6022 => x"70810651",
          6023 => x"5170802e",
          6024 => x"8d387193",
          6025 => x"2a708106",
          6026 => x"515170ff",
          6027 => x"be387481",
          6028 => x"ff065187",
          6029 => x"c0948052",
          6030 => x"70802e86",
          6031 => x"3887c094",
          6032 => x"90527772",
          6033 => x"0c811774",
          6034 => x"337081ff",
          6035 => x"06535357",
          6036 => x"70ff8638",
          6037 => x"7682d8c8",
          6038 => x"0c893d0d",
          6039 => x"04fe3d0d",
          6040 => x"82d6e833",
          6041 => x"7081ff06",
          6042 => x"545287c0",
          6043 => x"94845172",
          6044 => x"802e8638",
          6045 => x"87c09494",
          6046 => x"51700870",
          6047 => x"822a7081",
          6048 => x"06515151",
          6049 => x"70802ee2",
          6050 => x"387181ff",
          6051 => x"065187c0",
          6052 => x"94805270",
          6053 => x"802e8638",
          6054 => x"87c09490",
          6055 => x"52710870",
          6056 => x"81ff0682",
          6057 => x"d8c80c51",
          6058 => x"843d0d04",
          6059 => x"ffaf3f82",
          6060 => x"d8c80881",
          6061 => x"ff0682d8",
          6062 => x"c80c04fe",
          6063 => x"3d0d82d6",
          6064 => x"e8337081",
          6065 => x"ff065253",
          6066 => x"87c09484",
          6067 => x"5270802e",
          6068 => x"863887c0",
          6069 => x"94945271",
          6070 => x"0870822a",
          6071 => x"70810651",
          6072 => x"5151ff52",
          6073 => x"70802ea0",
          6074 => x"387281ff",
          6075 => x"065187c0",
          6076 => x"94805270",
          6077 => x"802e8638",
          6078 => x"87c09490",
          6079 => x"52710870",
          6080 => x"982b7098",
          6081 => x"2c515351",
          6082 => x"7182d8c8",
          6083 => x"0c843d0d",
          6084 => x"04ff3d0d",
          6085 => x"87c09e80",
          6086 => x"08709c2a",
          6087 => x"8a065151",
          6088 => x"70802e84",
          6089 => x"b43887c0",
          6090 => x"9ea40882",
          6091 => x"d6ec0c87",
          6092 => x"c09ea808",
          6093 => x"82d6f00c",
          6094 => x"87c09e94",
          6095 => x"0882d6f4",
          6096 => x"0c87c09e",
          6097 => x"980882d6",
          6098 => x"f80c87c0",
          6099 => x"9e9c0882",
          6100 => x"d6fc0c87",
          6101 => x"c09ea008",
          6102 => x"82d7800c",
          6103 => x"87c09eac",
          6104 => x"0882d784",
          6105 => x"0c87c09e",
          6106 => x"b00882d7",
          6107 => x"880c87c0",
          6108 => x"9eb40882",
          6109 => x"d78c0c87",
          6110 => x"c09eb808",
          6111 => x"82d7900c",
          6112 => x"87c09ebc",
          6113 => x"0882d794",
          6114 => x"0c87c09e",
          6115 => x"c00882d7",
          6116 => x"980c87c0",
          6117 => x"9ec40882",
          6118 => x"d79c0c87",
          6119 => x"c09e8008",
          6120 => x"517082d7",
          6121 => x"a02387c0",
          6122 => x"9e840882",
          6123 => x"d7a40c87",
          6124 => x"c09e8808",
          6125 => x"82d7a80c",
          6126 => x"87c09e8c",
          6127 => x"0882d7ac",
          6128 => x"0c810b82",
          6129 => x"d7b03480",
          6130 => x"0b87c09e",
          6131 => x"90087084",
          6132 => x"800a0651",
          6133 => x"52527080",
          6134 => x"2e833881",
          6135 => x"527182d7",
          6136 => x"b134800b",
          6137 => x"87c09e90",
          6138 => x"08708880",
          6139 => x"0a065152",
          6140 => x"5270802e",
          6141 => x"83388152",
          6142 => x"7182d7b2",
          6143 => x"34800b87",
          6144 => x"c09e9008",
          6145 => x"7090800a",
          6146 => x"06515252",
          6147 => x"70802e83",
          6148 => x"38815271",
          6149 => x"82d7b334",
          6150 => x"800b87c0",
          6151 => x"9e900870",
          6152 => x"88808006",
          6153 => x"51525270",
          6154 => x"802e8338",
          6155 => x"81527182",
          6156 => x"d7b43480",
          6157 => x"0b87c09e",
          6158 => x"900870a0",
          6159 => x"80800651",
          6160 => x"52527080",
          6161 => x"2e833881",
          6162 => x"527182d7",
          6163 => x"b534800b",
          6164 => x"87c09e90",
          6165 => x"08709080",
          6166 => x"80065152",
          6167 => x"5270802e",
          6168 => x"83388152",
          6169 => x"7182d7b6",
          6170 => x"34800b87",
          6171 => x"c09e9008",
          6172 => x"70848080",
          6173 => x"06515252",
          6174 => x"70802e83",
          6175 => x"38815271",
          6176 => x"82d7b734",
          6177 => x"800b87c0",
          6178 => x"9e900870",
          6179 => x"82808006",
          6180 => x"51525270",
          6181 => x"802e8338",
          6182 => x"81527182",
          6183 => x"d7b83480",
          6184 => x"0b87c09e",
          6185 => x"90087081",
          6186 => x"80800651",
          6187 => x"52527080",
          6188 => x"2e833881",
          6189 => x"527182d7",
          6190 => x"b934800b",
          6191 => x"87c09e90",
          6192 => x"087080c0",
          6193 => x"80065152",
          6194 => x"5270802e",
          6195 => x"83388152",
          6196 => x"7182d7ba",
          6197 => x"34800b87",
          6198 => x"c09e9008",
          6199 => x"70a08006",
          6200 => x"51525270",
          6201 => x"802e8338",
          6202 => x"81527182",
          6203 => x"d7bb3487",
          6204 => x"c09e9008",
          6205 => x"70988006",
          6206 => x"708a2a51",
          6207 => x"51517082",
          6208 => x"d7bc3480",
          6209 => x"0b87c09e",
          6210 => x"90087084",
          6211 => x"80065152",
          6212 => x"5270802e",
          6213 => x"83388152",
          6214 => x"7182d7bd",
          6215 => x"3487c09e",
          6216 => x"90087083",
          6217 => x"f0067084",
          6218 => x"2a515151",
          6219 => x"7082d7be",
          6220 => x"34800b87",
          6221 => x"c09e9008",
          6222 => x"70880651",
          6223 => x"52527080",
          6224 => x"2e833881",
          6225 => x"527182d7",
          6226 => x"bf3487c0",
          6227 => x"9e900870",
          6228 => x"87065151",
          6229 => x"7082d7c0",
          6230 => x"34833d0d",
          6231 => x"04fb3d0d",
          6232 => x"82c0c451",
          6233 => x"ff90f13f",
          6234 => x"82d7b033",
          6235 => x"5473802e",
          6236 => x"893882c0",
          6237 => x"d851ff90",
          6238 => x"df3f82c0",
          6239 => x"ec51ffac",
          6240 => x"e23f82d7",
          6241 => x"b2335473",
          6242 => x"802e9438",
          6243 => x"82d78c08",
          6244 => x"82d79008",
          6245 => x"11545282",
          6246 => x"c18451ff",
          6247 => x"90ba3f82",
          6248 => x"d7b73354",
          6249 => x"73802e94",
          6250 => x"3882d784",
          6251 => x"0882d788",
          6252 => x"08115452",
          6253 => x"82c1a051",
          6254 => x"ff909d3f",
          6255 => x"82d7b433",
          6256 => x"5473802e",
          6257 => x"943882d6",
          6258 => x"ec0882d6",
          6259 => x"f0081154",
          6260 => x"5282c1bc",
          6261 => x"51ff9080",
          6262 => x"3f82d7b5",
          6263 => x"33547380",
          6264 => x"2e943882",
          6265 => x"d6f40882",
          6266 => x"d6f80811",
          6267 => x"545282c1",
          6268 => x"d851ff8f",
          6269 => x"e33f82d7",
          6270 => x"b6335473",
          6271 => x"802e9438",
          6272 => x"82d6fc08",
          6273 => x"82d78008",
          6274 => x"11545282",
          6275 => x"c1f451ff",
          6276 => x"8fc63f82",
          6277 => x"d7bb3354",
          6278 => x"73802e8e",
          6279 => x"3882d7bc",
          6280 => x"335282c2",
          6281 => x"9051ff8f",
          6282 => x"af3f82d7",
          6283 => x"bf335473",
          6284 => x"802e8e38",
          6285 => x"82d7c033",
          6286 => x"5282c2b0",
          6287 => x"51ff8f98",
          6288 => x"3f82d7bd",
          6289 => x"33547380",
          6290 => x"2e8e3882",
          6291 => x"d7be3352",
          6292 => x"82c2d051",
          6293 => x"ff8f813f",
          6294 => x"82d7b133",
          6295 => x"5473802e",
          6296 => x"893882c2",
          6297 => x"f051ffaa",
          6298 => x"fa3f82d7",
          6299 => x"b3335473",
          6300 => x"802e8938",
          6301 => x"82c38451",
          6302 => x"ffaae83f",
          6303 => x"82d7b833",
          6304 => x"5473802e",
          6305 => x"893882c3",
          6306 => x"9051ffaa",
          6307 => x"d63f82d7",
          6308 => x"b9335473",
          6309 => x"802e8938",
          6310 => x"82c39c51",
          6311 => x"ffaac43f",
          6312 => x"82d7ba33",
          6313 => x"5473802e",
          6314 => x"893882c3",
          6315 => x"a451ffaa",
          6316 => x"b23f82c3",
          6317 => x"ac51ffaa",
          6318 => x"aa3f82d7",
          6319 => x"94085282",
          6320 => x"c3b851ff",
          6321 => x"8e923f82",
          6322 => x"d7980852",
          6323 => x"82c3e051",
          6324 => x"ff8e853f",
          6325 => x"82d79c08",
          6326 => x"5282c488",
          6327 => x"51ff8df8",
          6328 => x"3f82c4b0",
          6329 => x"51ffa9fb",
          6330 => x"3f82d7a0",
          6331 => x"225282c4",
          6332 => x"b851ff8d",
          6333 => x"e33f82d7",
          6334 => x"a40856bd",
          6335 => x"84c05275",
          6336 => x"51c1803f",
          6337 => x"82d8c808",
          6338 => x"bd84c029",
          6339 => x"76713154",
          6340 => x"5482d8c8",
          6341 => x"085282c4",
          6342 => x"e051ff8d",
          6343 => x"bb3f82d7",
          6344 => x"b7335473",
          6345 => x"802ea938",
          6346 => x"82d7a808",
          6347 => x"56bd84c0",
          6348 => x"527551c0",
          6349 => x"ce3f82d8",
          6350 => x"c808bd84",
          6351 => x"c0297671",
          6352 => x"31545482",
          6353 => x"d8c80852",
          6354 => x"82c58c51",
          6355 => x"ff8d893f",
          6356 => x"82d7b233",
          6357 => x"5473802e",
          6358 => x"a93882d7",
          6359 => x"ac0856bd",
          6360 => x"84c05275",
          6361 => x"51c09c3f",
          6362 => x"82d8c808",
          6363 => x"bd84c029",
          6364 => x"76713154",
          6365 => x"5482d8c8",
          6366 => x"085282c5",
          6367 => x"b851ff8c",
          6368 => x"d73f8a51",
          6369 => x"ffabfe3f",
          6370 => x"873d0d04",
          6371 => x"fe3d0d02",
          6372 => x"920533ff",
          6373 => x"05527184",
          6374 => x"26aa3871",
          6375 => x"842982af",
          6376 => x"c4055271",
          6377 => x"080482c5",
          6378 => x"e4519d39",
          6379 => x"82c5ec51",
          6380 => x"973982c5",
          6381 => x"f4519139",
          6382 => x"82c5fc51",
          6383 => x"8b3982c6",
          6384 => x"80518539",
          6385 => x"82c68851",
          6386 => x"ff8c8d3f",
          6387 => x"843d0d04",
          6388 => x"7188800c",
          6389 => x"04ff3d0d",
          6390 => x"87c09684",
          6391 => x"70085252",
          6392 => x"80720c70",
          6393 => x"74077082",
          6394 => x"d7c40c72",
          6395 => x"0c833d0d",
          6396 => x"04ff3d0d",
          6397 => x"87c09684",
          6398 => x"700882d7",
          6399 => x"c40c5280",
          6400 => x"720c7309",
          6401 => x"7082d7c4",
          6402 => x"08067082",
          6403 => x"d7c40c73",
          6404 => x"0c51833d",
          6405 => x"0d04800b",
          6406 => x"87c09684",
          6407 => x"0c0482d7",
          6408 => x"c40887c0",
          6409 => x"96840c04",
          6410 => x"fd3d0d76",
          6411 => x"982b7098",
          6412 => x"2c79982b",
          6413 => x"70982c72",
          6414 => x"10137082",
          6415 => x"2b515351",
          6416 => x"54515180",
          6417 => x"0b82c694",
          6418 => x"12335553",
          6419 => x"7174259c",
          6420 => x"3882c690",
          6421 => x"11081202",
          6422 => x"84059705",
          6423 => x"33713352",
          6424 => x"52527072",
          6425 => x"2e098106",
          6426 => x"83388153",
          6427 => x"7282d8c8",
          6428 => x"0c853d0d",
          6429 => x"04fb3d0d",
          6430 => x"79028405",
          6431 => x"a3053371",
          6432 => x"33555654",
          6433 => x"72802eb1",
          6434 => x"3882f4ac",
          6435 => x"08528851",
          6436 => x"ffaa9f3f",
          6437 => x"82f4ac08",
          6438 => x"52a051ff",
          6439 => x"aa943f82",
          6440 => x"f4ac0852",
          6441 => x"8851ffaa",
          6442 => x"893f7333",
          6443 => x"ff055372",
          6444 => x"74347281",
          6445 => x"ff0653cc",
          6446 => x"397751ff",
          6447 => x"8a9a3f74",
          6448 => x"7434873d",
          6449 => x"0d04f63d",
          6450 => x"0d7c0284",
          6451 => x"05b70533",
          6452 => x"028805bb",
          6453 => x"053382d8",
          6454 => x"a0337084",
          6455 => x"2982d7c8",
          6456 => x"05700851",
          6457 => x"59595a58",
          6458 => x"5974802e",
          6459 => x"86387451",
          6460 => x"9afa3f82",
          6461 => x"d8a03370",
          6462 => x"842982d7",
          6463 => x"c8058119",
          6464 => x"70545856",
          6465 => x"5a9dfb3f",
          6466 => x"82d8c808",
          6467 => x"750c82d8",
          6468 => x"a0337084",
          6469 => x"2982d7c8",
          6470 => x"05700851",
          6471 => x"565a7480",
          6472 => x"2ea73875",
          6473 => x"53785274",
          6474 => x"51ffb3b9",
          6475 => x"3f82d8a0",
          6476 => x"33810555",
          6477 => x"7482d8a0",
          6478 => x"347481ff",
          6479 => x"06559375",
          6480 => x"27873880",
          6481 => x"0b82d8a0",
          6482 => x"3477802e",
          6483 => x"b63882d8",
          6484 => x"9c085675",
          6485 => x"802eac38",
          6486 => x"82d89833",
          6487 => x"5574a438",
          6488 => x"8c3dfc05",
          6489 => x"54765378",
          6490 => x"52755180",
          6491 => x"ebbe3f82",
          6492 => x"d89c0852",
          6493 => x"8a5181a0",
          6494 => x"e73f82d8",
          6495 => x"9c085180",
          6496 => x"efa13f8c",
          6497 => x"3d0d04fd",
          6498 => x"3d0d82d7",
          6499 => x"c8539354",
          6500 => x"72085271",
          6501 => x"802e8938",
          6502 => x"715199d0",
          6503 => x"3f80730c",
          6504 => x"ff148414",
          6505 => x"54547380",
          6506 => x"25e63880",
          6507 => x"0b82d8a0",
          6508 => x"3482d89c",
          6509 => x"08527180",
          6510 => x"2e953871",
          6511 => x"5180f086",
          6512 => x"3f82d89c",
          6513 => x"085199a4",
          6514 => x"3f800b82",
          6515 => x"d89c0c85",
          6516 => x"3d0d04dc",
          6517 => x"3d0d8157",
          6518 => x"805282d8",
          6519 => x"9c085180",
          6520 => x"f5a23f82",
          6521 => x"d8c80880",
          6522 => x"d33882d8",
          6523 => x"9c085380",
          6524 => x"f852883d",
          6525 => x"70525681",
          6526 => x"9dd23f82",
          6527 => x"d8c80880",
          6528 => x"2eba3875",
          6529 => x"51ffaffd",
          6530 => x"3f82d8c8",
          6531 => x"0855800b",
          6532 => x"82d8c808",
          6533 => x"259d3882",
          6534 => x"d8c808ff",
          6535 => x"05701755",
          6536 => x"55807434",
          6537 => x"75537652",
          6538 => x"811782c9",
          6539 => x"845257ff",
          6540 => x"87a63f74",
          6541 => x"ff2e0981",
          6542 => x"06ffaf38",
          6543 => x"a63d0d04",
          6544 => x"d93d0daa",
          6545 => x"3d08ad3d",
          6546 => x"085a5a81",
          6547 => x"70585880",
          6548 => x"5282d89c",
          6549 => x"085180f4",
          6550 => x"ab3f82d8",
          6551 => x"c8088195",
          6552 => x"38ff0b82",
          6553 => x"d89c0854",
          6554 => x"5580f852",
          6555 => x"8b3d7052",
          6556 => x"56819cd8",
          6557 => x"3f82d8c8",
          6558 => x"08802ea5",
          6559 => x"387551ff",
          6560 => x"af833f82",
          6561 => x"d8c80881",
          6562 => x"18585580",
          6563 => x"0b82d8c8",
          6564 => x"08258e38",
          6565 => x"82d8c808",
          6566 => x"ff057017",
          6567 => x"55558074",
          6568 => x"34740970",
          6569 => x"30707207",
          6570 => x"9f2a5155",
          6571 => x"5578772e",
          6572 => x"853873ff",
          6573 => x"ac3882d8",
          6574 => x"9c088c11",
          6575 => x"08535180",
          6576 => x"f3c23f82",
          6577 => x"d8c80880",
          6578 => x"2e893882",
          6579 => x"c99051ff",
          6580 => x"86863f78",
          6581 => x"772e0981",
          6582 => x"069b3875",
          6583 => x"527951ff",
          6584 => x"af913f79",
          6585 => x"51ffae9d",
          6586 => x"3fab3d08",
          6587 => x"5482d8c8",
          6588 => x"08743480",
          6589 => x"587782d8",
          6590 => x"c80ca93d",
          6591 => x"0d04f63d",
          6592 => x"0d7c7e71",
          6593 => x"5c717233",
          6594 => x"57595a58",
          6595 => x"73a02e09",
          6596 => x"8106a238",
          6597 => x"78337805",
          6598 => x"56777627",
          6599 => x"98388117",
          6600 => x"705b7071",
          6601 => x"33565855",
          6602 => x"73a02e09",
          6603 => x"81068638",
          6604 => x"757526ea",
          6605 => x"38805473",
          6606 => x"882982d8",
          6607 => x"a4057008",
          6608 => x"5255ffad",
          6609 => x"c03f82d8",
          6610 => x"c8085379",
          6611 => x"52740851",
          6612 => x"ffb0bf3f",
          6613 => x"82d8c808",
          6614 => x"80c53884",
          6615 => x"15335574",
          6616 => x"812e8838",
          6617 => x"74822e88",
          6618 => x"38b539fc",
          6619 => x"e63fac39",
          6620 => x"811a5a8c",
          6621 => x"3dfc1153",
          6622 => x"f80551c0",
          6623 => x"cf3f82d8",
          6624 => x"c808802e",
          6625 => x"9a38ff1b",
          6626 => x"53785277",
          6627 => x"51fdb13f",
          6628 => x"82d8c808",
          6629 => x"81ff0655",
          6630 => x"74853874",
          6631 => x"54913981",
          6632 => x"147081ff",
          6633 => x"06515482",
          6634 => x"7427ff8b",
          6635 => x"38805473",
          6636 => x"82d8c80c",
          6637 => x"8c3d0d04",
          6638 => x"d33d0db0",
          6639 => x"3d08b23d",
          6640 => x"08b43d08",
          6641 => x"595f5a80",
          6642 => x"0baf3d34",
          6643 => x"82d8a033",
          6644 => x"82d89c08",
          6645 => x"555b7381",
          6646 => x"cb387382",
          6647 => x"d8983355",
          6648 => x"55738338",
          6649 => x"81557680",
          6650 => x"2e81bc38",
          6651 => x"81707606",
          6652 => x"55567380",
          6653 => x"2e81ad38",
          6654 => x"a8519886",
          6655 => x"3f82d8c8",
          6656 => x"0882d89c",
          6657 => x"0c82d8c8",
          6658 => x"08802e81",
          6659 => x"92389353",
          6660 => x"765282d8",
          6661 => x"c8085180",
          6662 => x"dead3f82",
          6663 => x"d8c80880",
          6664 => x"2e8c3882",
          6665 => x"c9bc51ff",
          6666 => x"9fb93f80",
          6667 => x"f73982d8",
          6668 => x"c8085b82",
          6669 => x"d89c0853",
          6670 => x"80f85290",
          6671 => x"3d705254",
          6672 => x"8199893f",
          6673 => x"82d8c808",
          6674 => x"5682d8c8",
          6675 => x"08742e09",
          6676 => x"810680d0",
          6677 => x"3882d8c8",
          6678 => x"0851ffab",
          6679 => x"a83f82d8",
          6680 => x"c8085580",
          6681 => x"0b82d8c8",
          6682 => x"0825a938",
          6683 => x"82d8c808",
          6684 => x"ff057017",
          6685 => x"55558074",
          6686 => x"34805374",
          6687 => x"81ff0652",
          6688 => x"7551f8c2",
          6689 => x"3f811b70",
          6690 => x"81ff065c",
          6691 => x"54937b27",
          6692 => x"8338805b",
          6693 => x"74ff2e09",
          6694 => x"8106ff97",
          6695 => x"38863975",
          6696 => x"82d89834",
          6697 => x"768c3882",
          6698 => x"d89c0880",
          6699 => x"2e8438f9",
          6700 => x"d63f8f3d",
          6701 => x"5dec843f",
          6702 => x"82d8c808",
          6703 => x"982b7098",
          6704 => x"2c515978",
          6705 => x"ff2eee38",
          6706 => x"7881ff06",
          6707 => x"82f08433",
          6708 => x"70982b70",
          6709 => x"982c82f0",
          6710 => x"80337098",
          6711 => x"2b70972c",
          6712 => x"71982c05",
          6713 => x"70842982",
          6714 => x"c6900570",
          6715 => x"08157033",
          6716 => x"51515151",
          6717 => x"59595159",
          6718 => x"5d588156",
          6719 => x"73782e80",
          6720 => x"e9387774",
          6721 => x"27b43874",
          6722 => x"81800a29",
          6723 => x"81ff0a05",
          6724 => x"70982c51",
          6725 => x"55807524",
          6726 => x"80ce3876",
          6727 => x"53745277",
          6728 => x"51f6853f",
          6729 => x"82d8c808",
          6730 => x"81ff0654",
          6731 => x"73802ed7",
          6732 => x"387482f0",
          6733 => x"80348156",
          6734 => x"b1397481",
          6735 => x"800a2981",
          6736 => x"800a0570",
          6737 => x"982c7081",
          6738 => x"ff065651",
          6739 => x"55739526",
          6740 => x"97387653",
          6741 => x"74527751",
          6742 => x"f5ce3f82",
          6743 => x"d8c80881",
          6744 => x"ff065473",
          6745 => x"cc38d339",
          6746 => x"80567580",
          6747 => x"2e80ca38",
          6748 => x"811c5574",
          6749 => x"82f08434",
          6750 => x"74982b70",
          6751 => x"982c82f0",
          6752 => x"80337098",
          6753 => x"2b70982c",
          6754 => x"70101170",
          6755 => x"822b82c6",
          6756 => x"9411335e",
          6757 => x"51515157",
          6758 => x"58515574",
          6759 => x"772e0981",
          6760 => x"06fe9238",
          6761 => x"82c69814",
          6762 => x"087d0c80",
          6763 => x"0b82f084",
          6764 => x"34800b82",
          6765 => x"f0803492",
          6766 => x"397582f0",
          6767 => x"84347582",
          6768 => x"f0803478",
          6769 => x"af3d3475",
          6770 => x"7d0c7e54",
          6771 => x"739526fd",
          6772 => x"e1387384",
          6773 => x"2982afd8",
          6774 => x"05547308",
          6775 => x"0482f08c",
          6776 => x"3354737e",
          6777 => x"2efdcb38",
          6778 => x"82f08833",
          6779 => x"55737527",
          6780 => x"ab387498",
          6781 => x"2b70982c",
          6782 => x"51557375",
          6783 => x"249e3874",
          6784 => x"1a547333",
          6785 => x"81153474",
          6786 => x"81800a29",
          6787 => x"81ff0a05",
          6788 => x"70982c82",
          6789 => x"f08c3356",
          6790 => x"5155df39",
          6791 => x"82f08c33",
          6792 => x"81115654",
          6793 => x"7482f08c",
          6794 => x"34731a54",
          6795 => x"ae3d3374",
          6796 => x"3482f088",
          6797 => x"3354737e",
          6798 => x"25893881",
          6799 => x"14547382",
          6800 => x"f0883482",
          6801 => x"f08c3370",
          6802 => x"81800a29",
          6803 => x"81ff0a05",
          6804 => x"70982c82",
          6805 => x"f088335a",
          6806 => x"51565674",
          6807 => x"7725a838",
          6808 => x"82f4ac08",
          6809 => x"52741a70",
          6810 => x"335254ff",
          6811 => x"9ec43f74",
          6812 => x"81800a29",
          6813 => x"81800a05",
          6814 => x"70982c82",
          6815 => x"f0883356",
          6816 => x"51557375",
          6817 => x"24da3882",
          6818 => x"f08c3370",
          6819 => x"982b7098",
          6820 => x"2c82f088",
          6821 => x"335a5156",
          6822 => x"56747725",
          6823 => x"fc943882",
          6824 => x"f4ac0852",
          6825 => x"8851ff9e",
          6826 => x"893f7481",
          6827 => x"800a2981",
          6828 => x"800a0570",
          6829 => x"982c82f0",
          6830 => x"88335651",
          6831 => x"55737524",
          6832 => x"de38fbee",
          6833 => x"39837a34",
          6834 => x"800b811b",
          6835 => x"3482f08c",
          6836 => x"53805282",
          6837 => x"b8b851f3",
          6838 => x"9c3f81fd",
          6839 => x"3982f08c",
          6840 => x"337081ff",
          6841 => x"06555573",
          6842 => x"802efbc6",
          6843 => x"3882f088",
          6844 => x"33ff0554",
          6845 => x"7382f088",
          6846 => x"34ff1554",
          6847 => x"7382f08c",
          6848 => x"3482f4ac",
          6849 => x"08528851",
          6850 => x"ff9da73f",
          6851 => x"82f08c33",
          6852 => x"70982b70",
          6853 => x"982c82f0",
          6854 => x"88335751",
          6855 => x"56577474",
          6856 => x"25ad3874",
          6857 => x"1a548114",
          6858 => x"33743482",
          6859 => x"f4ac0852",
          6860 => x"733351ff",
          6861 => x"9cfc3f74",
          6862 => x"81800a29",
          6863 => x"81800a05",
          6864 => x"70982c82",
          6865 => x"f0883358",
          6866 => x"51557575",
          6867 => x"24d53882",
          6868 => x"f4ac0852",
          6869 => x"a051ff9c",
          6870 => x"d93f82f0",
          6871 => x"8c337098",
          6872 => x"2b70982c",
          6873 => x"82f08833",
          6874 => x"57515657",
          6875 => x"747424fa",
          6876 => x"c13882f4",
          6877 => x"ac085288",
          6878 => x"51ff9cb6",
          6879 => x"3f748180",
          6880 => x"0a298180",
          6881 => x"0a057098",
          6882 => x"2c82f088",
          6883 => x"33585155",
          6884 => x"757525de",
          6885 => x"38fa9b39",
          6886 => x"82f08833",
          6887 => x"7a055480",
          6888 => x"743482f4",
          6889 => x"ac08528a",
          6890 => x"51ff9c86",
          6891 => x"3f82f088",
          6892 => x"527951f6",
          6893 => x"c93f82d8",
          6894 => x"c80881ff",
          6895 => x"06547396",
          6896 => x"3882f088",
          6897 => x"33547380",
          6898 => x"2e8f3881",
          6899 => x"53735279",
          6900 => x"51f1f33f",
          6901 => x"8439807a",
          6902 => x"34800b82",
          6903 => x"f08c3480",
          6904 => x"0b82f088",
          6905 => x"347982d8",
          6906 => x"c80caf3d",
          6907 => x"0d0482f0",
          6908 => x"8c335473",
          6909 => x"802ef9ba",
          6910 => x"3882f4ac",
          6911 => x"08528851",
          6912 => x"ff9baf3f",
          6913 => x"82f08c33",
          6914 => x"ff055473",
          6915 => x"82f08c34",
          6916 => x"7381ff06",
          6917 => x"54dd3982",
          6918 => x"f08c3382",
          6919 => x"f0883355",
          6920 => x"5573752e",
          6921 => x"f98c38ff",
          6922 => x"14547382",
          6923 => x"f0883474",
          6924 => x"982b7098",
          6925 => x"2c7581ff",
          6926 => x"06565155",
          6927 => x"747425ad",
          6928 => x"38741a54",
          6929 => x"81143374",
          6930 => x"3482f4ac",
          6931 => x"08527333",
          6932 => x"51ff9ade",
          6933 => x"3f748180",
          6934 => x"0a298180",
          6935 => x"0a057098",
          6936 => x"2c82f088",
          6937 => x"33585155",
          6938 => x"757524d5",
          6939 => x"3882f4ac",
          6940 => x"0852a051",
          6941 => x"ff9abb3f",
          6942 => x"82f08c33",
          6943 => x"70982b70",
          6944 => x"982c82f0",
          6945 => x"88335751",
          6946 => x"56577474",
          6947 => x"24f8a338",
          6948 => x"82f4ac08",
          6949 => x"528851ff",
          6950 => x"9a983f74",
          6951 => x"81800a29",
          6952 => x"81800a05",
          6953 => x"70982c82",
          6954 => x"f0883358",
          6955 => x"51557575",
          6956 => x"25de38f7",
          6957 => x"fd3982f0",
          6958 => x"8c337081",
          6959 => x"ff0682f0",
          6960 => x"88335956",
          6961 => x"54747727",
          6962 => x"f7e83882",
          6963 => x"f4ac0852",
          6964 => x"81145473",
          6965 => x"82f08c34",
          6966 => x"741a7033",
          6967 => x"5254ff99",
          6968 => x"d13f82f0",
          6969 => x"8c337081",
          6970 => x"ff0682f0",
          6971 => x"88335856",
          6972 => x"54757526",
          6973 => x"d638f7ba",
          6974 => x"3982f08c",
          6975 => x"53805282",
          6976 => x"b8b851ee",
          6977 => x"f03f800b",
          6978 => x"82f08c34",
          6979 => x"800b82f0",
          6980 => x"8834f79e",
          6981 => x"397ab038",
          6982 => x"82d89408",
          6983 => x"5574802e",
          6984 => x"a6387451",
          6985 => x"ffa1de3f",
          6986 => x"82d8c808",
          6987 => x"82f08834",
          6988 => x"82d8c808",
          6989 => x"81ff0681",
          6990 => x"05537452",
          6991 => x"7951ffa3",
          6992 => x"a43f935b",
          6993 => x"81c0397a",
          6994 => x"842982d7",
          6995 => x"c805fc11",
          6996 => x"08565474",
          6997 => x"802ea738",
          6998 => x"7451ffa1",
          6999 => x"a83f82d8",
          7000 => x"c80882f0",
          7001 => x"883482d8",
          7002 => x"c80881ff",
          7003 => x"06810553",
          7004 => x"74527951",
          7005 => x"ffa2ee3f",
          7006 => x"ff1b5480",
          7007 => x"fa397308",
          7008 => x"5574802e",
          7009 => x"f6ac3874",
          7010 => x"51ffa0f9",
          7011 => x"3f99397a",
          7012 => x"932e0981",
          7013 => x"06ae3882",
          7014 => x"d7c80855",
          7015 => x"74802ea4",
          7016 => x"387451ff",
          7017 => x"a0df3f82",
          7018 => x"d8c80882",
          7019 => x"f0883482",
          7020 => x"d8c80881",
          7021 => x"ff068105",
          7022 => x"53745279",
          7023 => x"51ffa2a5",
          7024 => x"3f80c339",
          7025 => x"7a842982",
          7026 => x"d7cc0570",
          7027 => x"08565474",
          7028 => x"802eab38",
          7029 => x"7451ffa0",
          7030 => x"ac3f82d8",
          7031 => x"c80882f0",
          7032 => x"883482d8",
          7033 => x"c80881ff",
          7034 => x"06810553",
          7035 => x"74527951",
          7036 => x"ffa1f23f",
          7037 => x"811b5473",
          7038 => x"81ff065b",
          7039 => x"89397482",
          7040 => x"f0883474",
          7041 => x"7a3482f0",
          7042 => x"8c5382f0",
          7043 => x"88335279",
          7044 => x"51ece23f",
          7045 => x"f59c3982",
          7046 => x"f08c3370",
          7047 => x"81ff0682",
          7048 => x"f0883359",
          7049 => x"56547477",
          7050 => x"27f58738",
          7051 => x"82f4ac08",
          7052 => x"52811454",
          7053 => x"7382f08c",
          7054 => x"34741a70",
          7055 => x"335254ff",
          7056 => x"96f03ff4",
          7057 => x"ed3982f0",
          7058 => x"8c335473",
          7059 => x"802ef4e2",
          7060 => x"3882f4ac",
          7061 => x"08528851",
          7062 => x"ff96d73f",
          7063 => x"82f08c33",
          7064 => x"ff055473",
          7065 => x"82f08c34",
          7066 => x"f4c839f9",
          7067 => x"3d0d83c0",
          7068 => x"800b82d8",
          7069 => x"c00c8480",
          7070 => x"0b82d8bc",
          7071 => x"23a08053",
          7072 => x"805283c0",
          7073 => x"8051ffa5",
          7074 => x"dd3f82d8",
          7075 => x"c0085480",
          7076 => x"58777434",
          7077 => x"81577681",
          7078 => x"153482d8",
          7079 => x"c0085477",
          7080 => x"84153476",
          7081 => x"85153482",
          7082 => x"d8c00854",
          7083 => x"77861534",
          7084 => x"76871534",
          7085 => x"82d8c008",
          7086 => x"82d8bc22",
          7087 => x"ff05fe80",
          7088 => x"80077083",
          7089 => x"ffff0670",
          7090 => x"882a5851",
          7091 => x"55567488",
          7092 => x"17347389",
          7093 => x"173482d8",
          7094 => x"bc227088",
          7095 => x"2982d8c0",
          7096 => x"0805f811",
          7097 => x"51555577",
          7098 => x"82153476",
          7099 => x"83153489",
          7100 => x"3d0d04ff",
          7101 => x"3d0d7352",
          7102 => x"81518472",
          7103 => x"278f38fb",
          7104 => x"12832a82",
          7105 => x"117083ff",
          7106 => x"ff065151",
          7107 => x"517082d8",
          7108 => x"c80c833d",
          7109 => x"0d04f93d",
          7110 => x"0d02a605",
          7111 => x"22028405",
          7112 => x"aa052271",
          7113 => x"0582d8c0",
          7114 => x"0871832b",
          7115 => x"71117483",
          7116 => x"2b731170",
          7117 => x"33811233",
          7118 => x"71882b07",
          7119 => x"02a405ae",
          7120 => x"05227181",
          7121 => x"ffff0607",
          7122 => x"70882a53",
          7123 => x"51525954",
          7124 => x"5b5b5753",
          7125 => x"54557177",
          7126 => x"34708118",
          7127 => x"3482d8c0",
          7128 => x"08147588",
          7129 => x"2a525470",
          7130 => x"82153474",
          7131 => x"83153482",
          7132 => x"d8c00870",
          7133 => x"17703381",
          7134 => x"12337188",
          7135 => x"2b077083",
          7136 => x"2b8ffff8",
          7137 => x"06515256",
          7138 => x"52710573",
          7139 => x"83ffff06",
          7140 => x"70882a54",
          7141 => x"54517182",
          7142 => x"12347281",
          7143 => x"ff065372",
          7144 => x"83123482",
          7145 => x"d8c00816",
          7146 => x"56717634",
          7147 => x"72811734",
          7148 => x"893d0d04",
          7149 => x"fb3d0d82",
          7150 => x"d8c00802",
          7151 => x"84059e05",
          7152 => x"2270832b",
          7153 => x"72118611",
          7154 => x"33871233",
          7155 => x"718b2b71",
          7156 => x"832b0758",
          7157 => x"5b595255",
          7158 => x"52720584",
          7159 => x"12338513",
          7160 => x"3371882b",
          7161 => x"0770882a",
          7162 => x"54565652",
          7163 => x"70841334",
          7164 => x"73851334",
          7165 => x"82d8c008",
          7166 => x"70148411",
          7167 => x"33851233",
          7168 => x"718b2b71",
          7169 => x"832b0756",
          7170 => x"59575272",
          7171 => x"05861233",
          7172 => x"87133371",
          7173 => x"882b0770",
          7174 => x"882a5456",
          7175 => x"56527086",
          7176 => x"13347387",
          7177 => x"133482d8",
          7178 => x"c0081370",
          7179 => x"33811233",
          7180 => x"71882b07",
          7181 => x"7081ffff",
          7182 => x"0670882a",
          7183 => x"53515353",
          7184 => x"53717334",
          7185 => x"70811434",
          7186 => x"873d0d04",
          7187 => x"fa3d0d02",
          7188 => x"a2052282",
          7189 => x"d8c00871",
          7190 => x"832b7111",
          7191 => x"70338112",
          7192 => x"3371882b",
          7193 => x"07708829",
          7194 => x"15703381",
          7195 => x"12337198",
          7196 => x"2b71902b",
          7197 => x"07535f53",
          7198 => x"55525a56",
          7199 => x"57535471",
          7200 => x"802580f6",
          7201 => x"387251fe",
          7202 => x"ab3f82d8",
          7203 => x"c0087016",
          7204 => x"70338112",
          7205 => x"33718b2b",
          7206 => x"71832b07",
          7207 => x"74117033",
          7208 => x"81123371",
          7209 => x"882b0770",
          7210 => x"832b8fff",
          7211 => x"f8065152",
          7212 => x"5451535a",
          7213 => x"58537205",
          7214 => x"74882a54",
          7215 => x"52728213",
          7216 => x"34738313",
          7217 => x"3482d8c0",
          7218 => x"08701670",
          7219 => x"33811233",
          7220 => x"718b2b71",
          7221 => x"832b0756",
          7222 => x"59575572",
          7223 => x"05703381",
          7224 => x"12337188",
          7225 => x"2b077081",
          7226 => x"ffff0670",
          7227 => x"882a5751",
          7228 => x"52585272",
          7229 => x"74347181",
          7230 => x"1534883d",
          7231 => x"0d04fb3d",
          7232 => x"0d82d8c0",
          7233 => x"08028405",
          7234 => x"9e052270",
          7235 => x"832b7211",
          7236 => x"82113383",
          7237 => x"1233718b",
          7238 => x"2b71832b",
          7239 => x"07595b59",
          7240 => x"52565273",
          7241 => x"05713381",
          7242 => x"13337188",
          7243 => x"2b07028c",
          7244 => x"05a20522",
          7245 => x"71077088",
          7246 => x"2a535153",
          7247 => x"53537173",
          7248 => x"34708114",
          7249 => x"3482d8c0",
          7250 => x"08701570",
          7251 => x"33811233",
          7252 => x"718b2b71",
          7253 => x"832b0756",
          7254 => x"59575272",
          7255 => x"05821233",
          7256 => x"83133371",
          7257 => x"882b0770",
          7258 => x"882a5455",
          7259 => x"56527082",
          7260 => x"13347283",
          7261 => x"133482d8",
          7262 => x"c0081482",
          7263 => x"11338312",
          7264 => x"3371882b",
          7265 => x"0782d8c8",
          7266 => x"0c525487",
          7267 => x"3d0d04f7",
          7268 => x"3d0d7b82",
          7269 => x"d8c00831",
          7270 => x"832a7083",
          7271 => x"ffff0670",
          7272 => x"535753fd",
          7273 => x"a73f82d8",
          7274 => x"c0087683",
          7275 => x"2b711182",
          7276 => x"11338312",
          7277 => x"33718b2b",
          7278 => x"71832b07",
          7279 => x"75117033",
          7280 => x"81123371",
          7281 => x"982b7190",
          7282 => x"2b075342",
          7283 => x"4051535b",
          7284 => x"58555954",
          7285 => x"7280258d",
          7286 => x"38828080",
          7287 => x"527551fe",
          7288 => x"9d3f8184",
          7289 => x"39841433",
          7290 => x"85153371",
          7291 => x"8b2b7183",
          7292 => x"2b077611",
          7293 => x"79882a53",
          7294 => x"51555855",
          7295 => x"76861434",
          7296 => x"7581ff06",
          7297 => x"56758714",
          7298 => x"3482d8c0",
          7299 => x"08701984",
          7300 => x"12338513",
          7301 => x"3371882b",
          7302 => x"0770882a",
          7303 => x"54575b56",
          7304 => x"53728416",
          7305 => x"34738516",
          7306 => x"3482d8c0",
          7307 => x"08185380",
          7308 => x"0b861434",
          7309 => x"800b8714",
          7310 => x"3482d8c0",
          7311 => x"08537684",
          7312 => x"14347585",
          7313 => x"143482d8",
          7314 => x"c0081870",
          7315 => x"33811233",
          7316 => x"71882b07",
          7317 => x"70828080",
          7318 => x"0770882a",
          7319 => x"53515556",
          7320 => x"54747434",
          7321 => x"72811534",
          7322 => x"8b3d0d04",
          7323 => x"ff3d0d73",
          7324 => x"5282d8c0",
          7325 => x"088438f7",
          7326 => x"f23f7180",
          7327 => x"2e863871",
          7328 => x"51fe8c3f",
          7329 => x"833d0d04",
          7330 => x"f53d0d80",
          7331 => x"7e5258f8",
          7332 => x"e23f82d8",
          7333 => x"c80883ff",
          7334 => x"ff0682d8",
          7335 => x"c0088411",
          7336 => x"33851233",
          7337 => x"71882b07",
          7338 => x"705f5956",
          7339 => x"585a81ff",
          7340 => x"ff597578",
          7341 => x"2e80cb38",
          7342 => x"75882917",
          7343 => x"70338112",
          7344 => x"3371882b",
          7345 => x"077081ff",
          7346 => x"ff067931",
          7347 => x"7083ffff",
          7348 => x"06707f27",
          7349 => x"52535156",
          7350 => x"59557779",
          7351 => x"278a3873",
          7352 => x"802e8538",
          7353 => x"75785a5b",
          7354 => x"84153385",
          7355 => x"16337188",
          7356 => x"2b075754",
          7357 => x"75c23878",
          7358 => x"81ffff2e",
          7359 => x"85387a79",
          7360 => x"59568076",
          7361 => x"832b82d8",
          7362 => x"c0081170",
          7363 => x"33811233",
          7364 => x"71882b07",
          7365 => x"7081ffff",
          7366 => x"0651525a",
          7367 => x"565c5573",
          7368 => x"752e8338",
          7369 => x"81558054",
          7370 => x"79782681",
          7371 => x"cc387454",
          7372 => x"74802e81",
          7373 => x"c438777a",
          7374 => x"2e098106",
          7375 => x"89387551",
          7376 => x"f8f23f81",
          7377 => x"ac398280",
          7378 => x"80537952",
          7379 => x"7551f7c6",
          7380 => x"3f82d8c0",
          7381 => x"08701c86",
          7382 => x"11338712",
          7383 => x"33718b2b",
          7384 => x"71832b07",
          7385 => x"535a5e55",
          7386 => x"74057a17",
          7387 => x"7083ffff",
          7388 => x"0670882a",
          7389 => x"5c595654",
          7390 => x"78841534",
          7391 => x"7681ff06",
          7392 => x"57768515",
          7393 => x"3482d8c0",
          7394 => x"0875832b",
          7395 => x"7111721e",
          7396 => x"86113387",
          7397 => x"12337188",
          7398 => x"2b077088",
          7399 => x"2a535b5e",
          7400 => x"535a5654",
          7401 => x"73861934",
          7402 => x"75871934",
          7403 => x"82d8c008",
          7404 => x"701c8411",
          7405 => x"33851233",
          7406 => x"718b2b71",
          7407 => x"832b0753",
          7408 => x"5d5a5574",
          7409 => x"05547886",
          7410 => x"15347687",
          7411 => x"153482d8",
          7412 => x"c0087016",
          7413 => x"711d8411",
          7414 => x"33851233",
          7415 => x"71882b07",
          7416 => x"70882a53",
          7417 => x"5a5f5256",
          7418 => x"54738416",
          7419 => x"34758516",
          7420 => x"3482d8c0",
          7421 => x"081b8405",
          7422 => x"547382d8",
          7423 => x"c80c8d3d",
          7424 => x"0d04fe3d",
          7425 => x"0d745282",
          7426 => x"d8c00884",
          7427 => x"38f4dc3f",
          7428 => x"71537180",
          7429 => x"2e8b3871",
          7430 => x"51fced3f",
          7431 => x"82d8c808",
          7432 => x"537282d8",
          7433 => x"c80c843d",
          7434 => x"0d04ee3d",
          7435 => x"0d646640",
          7436 => x"5c807042",
          7437 => x"4082d8c0",
          7438 => x"08602e09",
          7439 => x"81068438",
          7440 => x"f4a93f7b",
          7441 => x"8e387e51",
          7442 => x"ffb83f82",
          7443 => x"d8c80854",
          7444 => x"83c7397e",
          7445 => x"8b387b51",
          7446 => x"fc923f7e",
          7447 => x"5483ba39",
          7448 => x"7e51f58f",
          7449 => x"3f82d8c8",
          7450 => x"0883ffff",
          7451 => x"0682d8c0",
          7452 => x"087d7131",
          7453 => x"832a7083",
          7454 => x"ffff0670",
          7455 => x"832b7311",
          7456 => x"70338112",
          7457 => x"3371882b",
          7458 => x"07707531",
          7459 => x"7083ffff",
          7460 => x"06708829",
          7461 => x"fc057388",
          7462 => x"291a7033",
          7463 => x"81123371",
          7464 => x"882b0770",
          7465 => x"902b5344",
          7466 => x"4e534841",
          7467 => x"525c545b",
          7468 => x"415c565b",
          7469 => x"5b738025",
          7470 => x"8f387681",
          7471 => x"ffff0675",
          7472 => x"317083ff",
          7473 => x"ff064254",
          7474 => x"82163383",
          7475 => x"17337188",
          7476 => x"2b077088",
          7477 => x"291c7033",
          7478 => x"81123371",
          7479 => x"982b7190",
          7480 => x"2b075347",
          7481 => x"45525654",
          7482 => x"7380258b",
          7483 => x"38787531",
          7484 => x"7083ffff",
          7485 => x"06415477",
          7486 => x"7b2781fe",
          7487 => x"38601854",
          7488 => x"737b2e09",
          7489 => x"81068f38",
          7490 => x"7851f6c0",
          7491 => x"3f7a83ff",
          7492 => x"ff065881",
          7493 => x"e5397f8e",
          7494 => x"387a7424",
          7495 => x"89387851",
          7496 => x"f6aa3f81",
          7497 => x"a5397f18",
          7498 => x"557a7524",
          7499 => x"80c83879",
          7500 => x"1d821133",
          7501 => x"83123371",
          7502 => x"882b0753",
          7503 => x"5754f4f4",
          7504 => x"3f805278",
          7505 => x"51f7b73f",
          7506 => x"82d8c808",
          7507 => x"83ffff06",
          7508 => x"7e547c53",
          7509 => x"70832b82",
          7510 => x"d8c00811",
          7511 => x"84055355",
          7512 => x"59ff8eb7",
          7513 => x"3f82d8c0",
          7514 => x"08148405",
          7515 => x"7583ffff",
          7516 => x"06595c81",
          7517 => x"85396015",
          7518 => x"547a7424",
          7519 => x"80d43878",
          7520 => x"51f5c93f",
          7521 => x"82d8c008",
          7522 => x"1d821133",
          7523 => x"83123371",
          7524 => x"882b0753",
          7525 => x"4354f49c",
          7526 => x"3f805278",
          7527 => x"51f6df3f",
          7528 => x"82d8c808",
          7529 => x"83ffff06",
          7530 => x"7e547c53",
          7531 => x"70832b82",
          7532 => x"d8c00811",
          7533 => x"84055355",
          7534 => x"59ff8ddf",
          7535 => x"3f82d8c0",
          7536 => x"08148405",
          7537 => x"60620519",
          7538 => x"555c7383",
          7539 => x"ffff0658",
          7540 => x"a9397b7f",
          7541 => x"5254f9b0",
          7542 => x"3f82d8c8",
          7543 => x"085c82d8",
          7544 => x"c808802e",
          7545 => x"93387d53",
          7546 => x"735282d8",
          7547 => x"c80851ff",
          7548 => x"91f33f73",
          7549 => x"51f7983f",
          7550 => x"7a587a78",
          7551 => x"27993880",
          7552 => x"537a5278",
          7553 => x"51f28f3f",
          7554 => x"7a19832b",
          7555 => x"82d8c008",
          7556 => x"05840551",
          7557 => x"f6f93f7b",
          7558 => x"547382d8",
          7559 => x"c80c943d",
          7560 => x"0d04fc3d",
          7561 => x"0d777729",
          7562 => x"705254fb",
          7563 => x"d53f82d8",
          7564 => x"c8085582",
          7565 => x"d8c80880",
          7566 => x"2e8e3873",
          7567 => x"53805282",
          7568 => x"d8c80851",
          7569 => x"ff969f3f",
          7570 => x"7482d8c8",
          7571 => x"0c863d0d",
          7572 => x"04ff3d0d",
          7573 => x"028f0533",
          7574 => x"51815270",
          7575 => x"72268738",
          7576 => x"82d8c411",
          7577 => x"33527182",
          7578 => x"d8c80c83",
          7579 => x"3d0d04fc",
          7580 => x"3d0d029b",
          7581 => x"05330284",
          7582 => x"059f0533",
          7583 => x"56538351",
          7584 => x"72812680",
          7585 => x"e0387284",
          7586 => x"2b87c092",
          7587 => x"8c115351",
          7588 => x"88547480",
          7589 => x"2e843881",
          7590 => x"88547372",
          7591 => x"0c87c092",
          7592 => x"8c115181",
          7593 => x"710c850b",
          7594 => x"87c0988c",
          7595 => x"0c705271",
          7596 => x"08708206",
          7597 => x"51517080",
          7598 => x"2e8a3887",
          7599 => x"c0988c08",
          7600 => x"5170ec38",
          7601 => x"7108fc80",
          7602 => x"80065271",
          7603 => x"923887c0",
          7604 => x"988c0851",
          7605 => x"70802e87",
          7606 => x"387182d8",
          7607 => x"c4143482",
          7608 => x"d8c41333",
          7609 => x"517082d8",
          7610 => x"c80c863d",
          7611 => x"0d04f33d",
          7612 => x"0d606264",
          7613 => x"028c05bf",
          7614 => x"05335740",
          7615 => x"585b8374",
          7616 => x"525afecd",
          7617 => x"3f82d8c8",
          7618 => x"0881067a",
          7619 => x"54527181",
          7620 => x"be387172",
          7621 => x"75842b87",
          7622 => x"c0928011",
          7623 => x"87c0928c",
          7624 => x"1287c092",
          7625 => x"8413415a",
          7626 => x"40575a58",
          7627 => x"850b87c0",
          7628 => x"988c0c76",
          7629 => x"7d0c8476",
          7630 => x"0c750870",
          7631 => x"852a7081",
          7632 => x"06515354",
          7633 => x"71802e8e",
          7634 => x"387b0852",
          7635 => x"717b7081",
          7636 => x"055d3481",
          7637 => x"19598074",
          7638 => x"a2065353",
          7639 => x"71732e83",
          7640 => x"38815378",
          7641 => x"83ff268f",
          7642 => x"3872802e",
          7643 => x"8a3887c0",
          7644 => x"988c0852",
          7645 => x"71c33887",
          7646 => x"c0988c08",
          7647 => x"5271802e",
          7648 => x"87387884",
          7649 => x"802e9938",
          7650 => x"81760c87",
          7651 => x"c0928c15",
          7652 => x"53720870",
          7653 => x"82065152",
          7654 => x"71f738ff",
          7655 => x"1a5a8d39",
          7656 => x"84801781",
          7657 => x"197081ff",
          7658 => x"065a5357",
          7659 => x"79802e90",
          7660 => x"3873fc80",
          7661 => x"80065271",
          7662 => x"87387d78",
          7663 => x"26feed38",
          7664 => x"73fc8080",
          7665 => x"06527180",
          7666 => x"2e833881",
          7667 => x"52715372",
          7668 => x"82d8c80c",
          7669 => x"8f3d0d04",
          7670 => x"f33d0d60",
          7671 => x"6264028c",
          7672 => x"05bf0533",
          7673 => x"5740585b",
          7674 => x"83598074",
          7675 => x"5258fce1",
          7676 => x"3f82d8c8",
          7677 => x"08810679",
          7678 => x"54527178",
          7679 => x"2e098106",
          7680 => x"81b13877",
          7681 => x"74842b87",
          7682 => x"c0928011",
          7683 => x"87c0928c",
          7684 => x"1287c092",
          7685 => x"84134059",
          7686 => x"5f565a85",
          7687 => x"0b87c098",
          7688 => x"8c0c767d",
          7689 => x"0c82760c",
          7690 => x"80587508",
          7691 => x"70842a70",
          7692 => x"81065153",
          7693 => x"5471802e",
          7694 => x"8c387a70",
          7695 => x"81055c33",
          7696 => x"7c0c8118",
          7697 => x"5873812a",
          7698 => x"70810651",
          7699 => x"5271802e",
          7700 => x"8a3887c0",
          7701 => x"988c0852",
          7702 => x"71d03887",
          7703 => x"c0988c08",
          7704 => x"5271802e",
          7705 => x"87387784",
          7706 => x"802e9938",
          7707 => x"81760c87",
          7708 => x"c0928c15",
          7709 => x"53720870",
          7710 => x"82065152",
          7711 => x"71f738ff",
          7712 => x"19598d39",
          7713 => x"811a7081",
          7714 => x"ff068480",
          7715 => x"19595b52",
          7716 => x"78802e90",
          7717 => x"3873fc80",
          7718 => x"80065271",
          7719 => x"87387d7a",
          7720 => x"26fef838",
          7721 => x"73fc8080",
          7722 => x"06527180",
          7723 => x"2e833881",
          7724 => x"52715372",
          7725 => x"82d8c80c",
          7726 => x"8f3d0d04",
          7727 => x"fa3d0d7a",
          7728 => x"028405a3",
          7729 => x"05330288",
          7730 => x"05a70533",
          7731 => x"71545456",
          7732 => x"57fafe3f",
          7733 => x"82d8c808",
          7734 => x"81065383",
          7735 => x"547280fe",
          7736 => x"38850b87",
          7737 => x"c0988c0c",
          7738 => x"81567176",
          7739 => x"2e80dc38",
          7740 => x"71762493",
          7741 => x"3874842b",
          7742 => x"87c0928c",
          7743 => x"11545471",
          7744 => x"802e8d38",
          7745 => x"80d43971",
          7746 => x"832e80c6",
          7747 => x"3880cb39",
          7748 => x"72087081",
          7749 => x"2a708106",
          7750 => x"51515271",
          7751 => x"802e8a38",
          7752 => x"87c0988c",
          7753 => x"085271e8",
          7754 => x"3887c098",
          7755 => x"8c085271",
          7756 => x"96388173",
          7757 => x"0c87c092",
          7758 => x"8c145372",
          7759 => x"08708206",
          7760 => x"515271f7",
          7761 => x"38963980",
          7762 => x"56923988",
          7763 => x"800a770c",
          7764 => x"85398180",
          7765 => x"770c7256",
          7766 => x"83398456",
          7767 => x"75547382",
          7768 => x"d8c80c88",
          7769 => x"3d0d04fe",
          7770 => x"3d0d7481",
          7771 => x"11337133",
          7772 => x"71882b07",
          7773 => x"82d8c80c",
          7774 => x"5351843d",
          7775 => x"0d04fd3d",
          7776 => x"0d758311",
          7777 => x"33821233",
          7778 => x"71902b71",
          7779 => x"882b0781",
          7780 => x"14337072",
          7781 => x"07882b75",
          7782 => x"33710782",
          7783 => x"d8c80c52",
          7784 => x"53545654",
          7785 => x"52853d0d",
          7786 => x"04ff3d0d",
          7787 => x"73028405",
          7788 => x"92052252",
          7789 => x"52707270",
          7790 => x"81055434",
          7791 => x"70882a51",
          7792 => x"70723483",
          7793 => x"3d0d04ff",
          7794 => x"3d0d7375",
          7795 => x"52527072",
          7796 => x"70810554",
          7797 => x"3470882a",
          7798 => x"51707270",
          7799 => x"81055434",
          7800 => x"70882a51",
          7801 => x"70727081",
          7802 => x"05543470",
          7803 => x"882a5170",
          7804 => x"7234833d",
          7805 => x"0d04fe3d",
          7806 => x"0d767577",
          7807 => x"54545170",
          7808 => x"802e9238",
          7809 => x"71708105",
          7810 => x"53337370",
          7811 => x"81055534",
          7812 => x"ff1151eb",
          7813 => x"39843d0d",
          7814 => x"04fe3d0d",
          7815 => x"75777654",
          7816 => x"52537272",
          7817 => x"70810554",
          7818 => x"34ff1151",
          7819 => x"70f43884",
          7820 => x"3d0d04fc",
          7821 => x"3d0d7877",
          7822 => x"79565653",
          7823 => x"74708105",
          7824 => x"56337470",
          7825 => x"81055633",
          7826 => x"717131ff",
          7827 => x"16565252",
          7828 => x"5272802e",
          7829 => x"86387180",
          7830 => x"2ee23871",
          7831 => x"82d8c80c",
          7832 => x"863d0d04",
          7833 => x"fe3d0d74",
          7834 => x"76545189",
          7835 => x"3971732e",
          7836 => x"8a388111",
          7837 => x"51703352",
          7838 => x"71f33870",
          7839 => x"3382d8c8",
          7840 => x"0c843d0d",
          7841 => x"04800b82",
          7842 => x"d8c80c04",
          7843 => x"fb3d0d77",
          7844 => x"70087070",
          7845 => x"81055233",
          7846 => x"70545555",
          7847 => x"56e73fff",
          7848 => x"5582d8c8",
          7849 => x"08a23872",
          7850 => x"802e9838",
          7851 => x"83b55272",
          7852 => x"5180f7b6",
          7853 => x"3f82d8c8",
          7854 => x"0883ffff",
          7855 => x"06537280",
          7856 => x"2e863873",
          7857 => x"760c7255",
          7858 => x"7482d8c8",
          7859 => x"0c873d0d",
          7860 => x"04f73d0d",
          7861 => x"7b56800b",
          7862 => x"83173356",
          7863 => x"5a747a2e",
          7864 => x"80d63881",
          7865 => x"54b41608",
          7866 => x"53b81670",
          7867 => x"53811733",
          7868 => x"5259f9e4",
          7869 => x"3f82d8c8",
          7870 => x"087a2e09",
          7871 => x"8106b738",
          7872 => x"82d8c808",
          7873 => x"831734b4",
          7874 => x"160870a8",
          7875 => x"180831a0",
          7876 => x"18085956",
          7877 => x"58747727",
          7878 => x"9f388216",
          7879 => x"33557482",
          7880 => x"2e098106",
          7881 => x"93388154",
          7882 => x"76185378",
          7883 => x"52811633",
          7884 => x"51f9a53f",
          7885 => x"8339815a",
          7886 => x"7982d8c8",
          7887 => x"0c8b3d0d",
          7888 => x"04fa3d0d",
          7889 => x"787a5656",
          7890 => x"805774b4",
          7891 => x"17082eaf",
          7892 => x"387551fe",
          7893 => x"fc3f82d8",
          7894 => x"c8085782",
          7895 => x"d8c8089f",
          7896 => x"38815474",
          7897 => x"53b81652",
          7898 => x"81163351",
          7899 => x"f7803f82",
          7900 => x"d8c80880",
          7901 => x"2e8538ff",
          7902 => x"55815774",
          7903 => x"b4170c76",
          7904 => x"82d8c80c",
          7905 => x"883d0d04",
          7906 => x"f83d0d7a",
          7907 => x"705257fe",
          7908 => x"c03f82d8",
          7909 => x"c8085882",
          7910 => x"d8c80881",
          7911 => x"91387633",
          7912 => x"5574832e",
          7913 => x"09810680",
          7914 => x"f0388417",
          7915 => x"33597881",
          7916 => x"2e098106",
          7917 => x"80e33884",
          7918 => x"805382d8",
          7919 => x"c80852b8",
          7920 => x"17705256",
          7921 => x"fcd33f82",
          7922 => x"d4d55284",
          7923 => x"b61751fb",
          7924 => x"d83f848b",
          7925 => x"85a4d252",
          7926 => x"7551fbeb",
          7927 => x"3f868a85",
          7928 => x"e4f25284",
          7929 => x"9c1751fb",
          7930 => x"de3f9417",
          7931 => x"085284a0",
          7932 => x"1751fbd3",
          7933 => x"3f901708",
          7934 => x"5284a417",
          7935 => x"51fbc83f",
          7936 => x"a4170881",
          7937 => x"0570b419",
          7938 => x"0c795553",
          7939 => x"75528117",
          7940 => x"3351f7c4",
          7941 => x"3f778418",
          7942 => x"34805380",
          7943 => x"52811733",
          7944 => x"51f9993f",
          7945 => x"82d8c808",
          7946 => x"802e8338",
          7947 => x"81587782",
          7948 => x"d8c80c8a",
          7949 => x"3d0d04fb",
          7950 => x"3d0d77fe",
          7951 => x"1a9c1208",
          7952 => x"fe055556",
          7953 => x"54805674",
          7954 => x"73278d38",
          7955 => x"8a142275",
          7956 => x"7129b016",
          7957 => x"08055753",
          7958 => x"7582d8c8",
          7959 => x"0c873d0d",
          7960 => x"04f93d0d",
          7961 => x"7a7a7008",
          7962 => x"56545781",
          7963 => x"772781df",
          7964 => x"38769c15",
          7965 => x"082781d7",
          7966 => x"38ff7433",
          7967 => x"54587282",
          7968 => x"2e80f538",
          7969 => x"72822489",
          7970 => x"3872812e",
          7971 => x"8d3881bf",
          7972 => x"3972832e",
          7973 => x"818e3881",
          7974 => x"b6397681",
          7975 => x"2a177089",
          7976 => x"2aa81608",
          7977 => x"05537452",
          7978 => x"55fd963f",
          7979 => x"82d8c808",
          7980 => x"819f3874",
          7981 => x"83ff0614",
          7982 => x"b8113381",
          7983 => x"1770892a",
          7984 => x"a8180805",
          7985 => x"55765457",
          7986 => x"5753fcf5",
          7987 => x"3f82d8c8",
          7988 => x"0880fe38",
          7989 => x"7483ff06",
          7990 => x"14b81133",
          7991 => x"70882b78",
          7992 => x"07798106",
          7993 => x"71842a5c",
          7994 => x"52585153",
          7995 => x"7280e238",
          7996 => x"759fff06",
          7997 => x"5880da39",
          7998 => x"76882aa8",
          7999 => x"15080552",
          8000 => x"7351fcbd",
          8001 => x"3f82d8c8",
          8002 => x"0880c638",
          8003 => x"761083fe",
          8004 => x"067405b8",
          8005 => x"0551f8cf",
          8006 => x"3f82d8c8",
          8007 => x"0883ffff",
          8008 => x"0658ae39",
          8009 => x"76872aa8",
          8010 => x"15080552",
          8011 => x"7351fc91",
          8012 => x"3f82d8c8",
          8013 => x"089b3876",
          8014 => x"822b83fc",
          8015 => x"067405b8",
          8016 => x"0551f8ba",
          8017 => x"3f82d8c8",
          8018 => x"08f00a06",
          8019 => x"58833981",
          8020 => x"587782d8",
          8021 => x"c80c893d",
          8022 => x"0d04f83d",
          8023 => x"0d7a7c7e",
          8024 => x"5a585682",
          8025 => x"59817727",
          8026 => x"829e3876",
          8027 => x"9c170827",
          8028 => x"82963875",
          8029 => x"33537279",
          8030 => x"2e819d38",
          8031 => x"72792489",
          8032 => x"3872812e",
          8033 => x"8d388280",
          8034 => x"3972832e",
          8035 => x"81b83881",
          8036 => x"f7397681",
          8037 => x"2a177089",
          8038 => x"2aa81808",
          8039 => x"05537652",
          8040 => x"55fb9e3f",
          8041 => x"82d8c808",
          8042 => x"5982d8c8",
          8043 => x"0881d938",
          8044 => x"7483ff06",
          8045 => x"16b80581",
          8046 => x"16788106",
          8047 => x"59565477",
          8048 => x"5376802e",
          8049 => x"8f387784",
          8050 => x"2b9ff006",
          8051 => x"74338f06",
          8052 => x"71075153",
          8053 => x"72743481",
          8054 => x"0b831734",
          8055 => x"74892aa8",
          8056 => x"17080552",
          8057 => x"7551fad9",
          8058 => x"3f82d8c8",
          8059 => x"085982d8",
          8060 => x"c8088194",
          8061 => x"387483ff",
          8062 => x"0616b805",
          8063 => x"78842a54",
          8064 => x"54768f38",
          8065 => x"77882a74",
          8066 => x"3381f006",
          8067 => x"718f0607",
          8068 => x"51537274",
          8069 => x"3480ec39",
          8070 => x"76882aa8",
          8071 => x"17080552",
          8072 => x"7551fa9d",
          8073 => x"3f82d8c8",
          8074 => x"085982d8",
          8075 => x"c80880d8",
          8076 => x"387783ff",
          8077 => x"ff065276",
          8078 => x"1083fe06",
          8079 => x"7605b805",
          8080 => x"51f6e63f",
          8081 => x"be397687",
          8082 => x"2aa81708",
          8083 => x"05527551",
          8084 => x"f9ef3f82",
          8085 => x"d8c80859",
          8086 => x"82d8c808",
          8087 => x"ab3877f0",
          8088 => x"0a067782",
          8089 => x"2b83fc06",
          8090 => x"7018b805",
          8091 => x"70545154",
          8092 => x"54f68b3f",
          8093 => x"82d8c808",
          8094 => x"8f0a0674",
          8095 => x"07527251",
          8096 => x"f6c53f81",
          8097 => x"0b831734",
          8098 => x"7882d8c8",
          8099 => x"0c8a3d0d",
          8100 => x"04f83d0d",
          8101 => x"7a7c7e72",
          8102 => x"08595656",
          8103 => x"59817527",
          8104 => x"a438749c",
          8105 => x"1708279d",
          8106 => x"3873802e",
          8107 => x"aa38ff53",
          8108 => x"73527551",
          8109 => x"fda43f82",
          8110 => x"d8c80854",
          8111 => x"82d8c808",
          8112 => x"80f23893",
          8113 => x"39825480",
          8114 => x"eb398154",
          8115 => x"80e63982",
          8116 => x"d8c80854",
          8117 => x"80de3974",
          8118 => x"527851fb",
          8119 => x"843f82d8",
          8120 => x"c8085882",
          8121 => x"d8c80880",
          8122 => x"2e80c738",
          8123 => x"82d8c808",
          8124 => x"812ed238",
          8125 => x"82d8c808",
          8126 => x"ff2ecf38",
          8127 => x"80537452",
          8128 => x"7551fcd6",
          8129 => x"3f82d8c8",
          8130 => x"08c5389c",
          8131 => x"1608fe11",
          8132 => x"94180857",
          8133 => x"55577474",
          8134 => x"27903881",
          8135 => x"1594170c",
          8136 => x"84163381",
          8137 => x"07547384",
          8138 => x"17347755",
          8139 => x"767826ff",
          8140 => x"a6388054",
          8141 => x"7382d8c8",
          8142 => x"0c8a3d0d",
          8143 => x"04f63d0d",
          8144 => x"7c7e7108",
          8145 => x"595b5b79",
          8146 => x"95389017",
          8147 => x"08587780",
          8148 => x"2e88389c",
          8149 => x"17087826",
          8150 => x"b2388158",
          8151 => x"ae397952",
          8152 => x"7a51f9fd",
          8153 => x"3f815574",
          8154 => x"82d8c808",
          8155 => x"2782e038",
          8156 => x"82d8c808",
          8157 => x"5582d8c8",
          8158 => x"08ff2e82",
          8159 => x"d2389c17",
          8160 => x"0882d8c8",
          8161 => x"082682c7",
          8162 => x"38795894",
          8163 => x"17087056",
          8164 => x"5473802e",
          8165 => x"82b93877",
          8166 => x"7a2e0981",
          8167 => x"0680e238",
          8168 => x"811a569c",
          8169 => x"17087626",
          8170 => x"83388256",
          8171 => x"75527a51",
          8172 => x"f9af3f80",
          8173 => x"5982d8c8",
          8174 => x"08812e09",
          8175 => x"81068638",
          8176 => x"82d8c808",
          8177 => x"5982d8c8",
          8178 => x"08097030",
          8179 => x"70720780",
          8180 => x"25707c07",
          8181 => x"82d8c808",
          8182 => x"54515155",
          8183 => x"557381ef",
          8184 => x"3882d8c8",
          8185 => x"08802e95",
          8186 => x"38901708",
          8187 => x"54817427",
          8188 => x"9038739c",
          8189 => x"18082789",
          8190 => x"38735885",
          8191 => x"397580db",
          8192 => x"38775681",
          8193 => x"16569c17",
          8194 => x"08762689",
          8195 => x"38825675",
          8196 => x"782681ac",
          8197 => x"3875527a",
          8198 => x"51f8c63f",
          8199 => x"82d8c808",
          8200 => x"802eb838",
          8201 => x"805982d8",
          8202 => x"c808812e",
          8203 => x"09810686",
          8204 => x"3882d8c8",
          8205 => x"085982d8",
          8206 => x"c8080970",
          8207 => x"30707207",
          8208 => x"8025707c",
          8209 => x"07515155",
          8210 => x"557380f8",
          8211 => x"3875782e",
          8212 => x"098106ff",
          8213 => x"ae387355",
          8214 => x"80f539ff",
          8215 => x"53755276",
          8216 => x"51f9f73f",
          8217 => x"82d8c808",
          8218 => x"82d8c808",
          8219 => x"307082d8",
          8220 => x"c8080780",
          8221 => x"25515555",
          8222 => x"79802e94",
          8223 => x"3873802e",
          8224 => x"8f387553",
          8225 => x"79527651",
          8226 => x"f9d03f82",
          8227 => x"d8c80855",
          8228 => x"74a53875",
          8229 => x"90180c9c",
          8230 => x"1708fe05",
          8231 => x"94180856",
          8232 => x"54747426",
          8233 => x"8638ff15",
          8234 => x"94180c84",
          8235 => x"17338107",
          8236 => x"54738418",
          8237 => x"349739ff",
          8238 => x"5674812e",
          8239 => x"90388c39",
          8240 => x"80558c39",
          8241 => x"82d8c808",
          8242 => x"55853981",
          8243 => x"56755574",
          8244 => x"82d8c80c",
          8245 => x"8c3d0d04",
          8246 => x"f83d0d7a",
          8247 => x"705255f3",
          8248 => x"f03f82d8",
          8249 => x"c8085881",
          8250 => x"5682d8c8",
          8251 => x"0880d838",
          8252 => x"7b527451",
          8253 => x"f6c13f82",
          8254 => x"d8c80882",
          8255 => x"d8c808b4",
          8256 => x"170c5984",
          8257 => x"80537752",
          8258 => x"b8157052",
          8259 => x"57f28a3f",
          8260 => x"77568439",
          8261 => x"8116568a",
          8262 => x"15225875",
          8263 => x"78279738",
          8264 => x"81547519",
          8265 => x"53765281",
          8266 => x"153351ed",
          8267 => x"ab3f82d8",
          8268 => x"c808802e",
          8269 => x"df388a15",
          8270 => x"22763270",
          8271 => x"30707207",
          8272 => x"709f2a53",
          8273 => x"51565675",
          8274 => x"82d8c80c",
          8275 => x"8a3d0d04",
          8276 => x"f83d0d7a",
          8277 => x"7c710858",
          8278 => x"565774f0",
          8279 => x"800a2680",
          8280 => x"f138749f",
          8281 => x"06537280",
          8282 => x"e9387490",
          8283 => x"180c8817",
          8284 => x"085473aa",
          8285 => x"38753353",
          8286 => x"82732788",
          8287 => x"38ac1608",
          8288 => x"54739b38",
          8289 => x"74852a53",
          8290 => x"820b8817",
          8291 => x"225a5872",
          8292 => x"792780fe",
          8293 => x"38ac1608",
          8294 => x"98180c80",
          8295 => x"cd398a16",
          8296 => x"2270892b",
          8297 => x"54587275",
          8298 => x"26b23873",
          8299 => x"527651f5",
          8300 => x"b03f82d8",
          8301 => x"c8085482",
          8302 => x"d8c808ff",
          8303 => x"2ebd3881",
          8304 => x"0b82d8c8",
          8305 => x"08278b38",
          8306 => x"9c160882",
          8307 => x"d8c80826",
          8308 => x"85388258",
          8309 => x"bd397473",
          8310 => x"3155cb39",
          8311 => x"73527551",
          8312 => x"f4d53f82",
          8313 => x"d8c80898",
          8314 => x"180c7394",
          8315 => x"180c9817",
          8316 => x"08538258",
          8317 => x"72802e9a",
          8318 => x"38853981",
          8319 => x"58943974",
          8320 => x"892a1398",
          8321 => x"180c7483",
          8322 => x"ff0616b8",
          8323 => x"059c180c",
          8324 => x"80587782",
          8325 => x"d8c80c8a",
          8326 => x"3d0d04f8",
          8327 => x"3d0d7a70",
          8328 => x"08901208",
          8329 => x"a0055957",
          8330 => x"54f0800a",
          8331 => x"77278638",
          8332 => x"800b9815",
          8333 => x"0c981408",
          8334 => x"53845572",
          8335 => x"802e81cb",
          8336 => x"387683ff",
          8337 => x"06587781",
          8338 => x"b5388113",
          8339 => x"98150c94",
          8340 => x"14085574",
          8341 => x"92387685",
          8342 => x"2a881722",
          8343 => x"56537473",
          8344 => x"26819b38",
          8345 => x"80c0398a",
          8346 => x"1622ff05",
          8347 => x"77892a06",
          8348 => x"5372818a",
          8349 => x"38745273",
          8350 => x"51f3e63f",
          8351 => x"82d8c808",
          8352 => x"53825581",
          8353 => x"0b82d8c8",
          8354 => x"082780ff",
          8355 => x"38815582",
          8356 => x"d8c808ff",
          8357 => x"2e80f438",
          8358 => x"9c160882",
          8359 => x"d8c80826",
          8360 => x"80ca387b",
          8361 => x"8a387798",
          8362 => x"150c8455",
          8363 => x"80dd3994",
          8364 => x"14085273",
          8365 => x"51f9863f",
          8366 => x"82d8c808",
          8367 => x"53875582",
          8368 => x"d8c80880",
          8369 => x"2e80c438",
          8370 => x"825582d8",
          8371 => x"c808812e",
          8372 => x"ba388155",
          8373 => x"82d8c808",
          8374 => x"ff2eb038",
          8375 => x"82d8c808",
          8376 => x"527551fb",
          8377 => x"f33f82d8",
          8378 => x"c808a038",
          8379 => x"7294150c",
          8380 => x"72527551",
          8381 => x"f2c13f82",
          8382 => x"d8c80898",
          8383 => x"150c7690",
          8384 => x"150c7716",
          8385 => x"b8059c15",
          8386 => x"0c805574",
          8387 => x"82d8c80c",
          8388 => x"8a3d0d04",
          8389 => x"f73d0d7b",
          8390 => x"7d71085b",
          8391 => x"5b578052",
          8392 => x"7651fcac",
          8393 => x"3f82d8c8",
          8394 => x"085482d8",
          8395 => x"c80880ec",
          8396 => x"3882d8c8",
          8397 => x"08569817",
          8398 => x"08527851",
          8399 => x"f0833f82",
          8400 => x"d8c80854",
          8401 => x"82d8c808",
          8402 => x"80d23882",
          8403 => x"d8c8089c",
          8404 => x"18087033",
          8405 => x"51545872",
          8406 => x"81e52e09",
          8407 => x"81068338",
          8408 => x"815882d8",
          8409 => x"c8085572",
          8410 => x"83388155",
          8411 => x"77750753",
          8412 => x"72802e8e",
          8413 => x"38811656",
          8414 => x"757a2e09",
          8415 => x"81068838",
          8416 => x"a53982d8",
          8417 => x"c8085681",
          8418 => x"527651fd",
          8419 => x"8e3f82d8",
          8420 => x"c8085482",
          8421 => x"d8c80880",
          8422 => x"2eff9b38",
          8423 => x"73842e09",
          8424 => x"81068338",
          8425 => x"87547382",
          8426 => x"d8c80c8b",
          8427 => x"3d0d04fd",
          8428 => x"3d0d769a",
          8429 => x"115254eb",
          8430 => x"ae3f82d8",
          8431 => x"c80883ff",
          8432 => x"ff067670",
          8433 => x"33515353",
          8434 => x"71832e09",
          8435 => x"81069038",
          8436 => x"941451eb",
          8437 => x"923f82d8",
          8438 => x"c808902b",
          8439 => x"73075372",
          8440 => x"82d8c80c",
          8441 => x"853d0d04",
          8442 => x"fc3d0d77",
          8443 => x"797083ff",
          8444 => x"ff06549a",
          8445 => x"12535555",
          8446 => x"ebaf3f76",
          8447 => x"70335153",
          8448 => x"72832e09",
          8449 => x"81068b38",
          8450 => x"73902a52",
          8451 => x"941551eb",
          8452 => x"983f863d",
          8453 => x"0d04fd3d",
          8454 => x"0d755480",
          8455 => x"518b5370",
          8456 => x"812a7181",
          8457 => x"80290574",
          8458 => x"70810556",
          8459 => x"33710570",
          8460 => x"81ff06ff",
          8461 => x"16565151",
          8462 => x"5172e438",
          8463 => x"7082d8c8",
          8464 => x"0c853d0d",
          8465 => x"04f23d0d",
          8466 => x"60624059",
          8467 => x"8479085f",
          8468 => x"5b81ff70",
          8469 => x"5d5d9819",
          8470 => x"08802e83",
          8471 => x"80389819",
          8472 => x"08527d51",
          8473 => x"eddb3f82",
          8474 => x"d8c8085b",
          8475 => x"82d8c808",
          8476 => x"82eb389c",
          8477 => x"19087033",
          8478 => x"55557386",
          8479 => x"38845b82",
          8480 => x"dc398b15",
          8481 => x"33bf0670",
          8482 => x"81ff0658",
          8483 => x"5372861a",
          8484 => x"3482d8c8",
          8485 => x"08567381",
          8486 => x"e52e0981",
          8487 => x"06833881",
          8488 => x"5682d8c8",
          8489 => x"085373ae",
          8490 => x"2e098106",
          8491 => x"83388153",
          8492 => x"75730753",
          8493 => x"72993882",
          8494 => x"d8c80877",
          8495 => x"df065456",
          8496 => x"72882e09",
          8497 => x"81068338",
          8498 => x"8156757f",
          8499 => x"2e873881",
          8500 => x"ff5c81ef",
          8501 => x"39768f2e",
          8502 => x"09810681",
          8503 => x"ca387386",
          8504 => x"2a708106",
          8505 => x"51537280",
          8506 => x"2e92388d",
          8507 => x"15337481",
          8508 => x"bf067090",
          8509 => x"1c08ac1d",
          8510 => x"0c565d5d",
          8511 => x"737c2e09",
          8512 => x"8106819c",
          8513 => x"388d1533",
          8514 => x"537c732e",
          8515 => x"09810681",
          8516 => x"8f388c1e",
          8517 => x"089a1652",
          8518 => x"5ae8cc3f",
          8519 => x"82d8c808",
          8520 => x"83ffff06",
          8521 => x"537280f8",
          8522 => x"38743370",
          8523 => x"81bf068d",
          8524 => x"29f30551",
          8525 => x"54817b58",
          8526 => x"5882cad0",
          8527 => x"17337505",
          8528 => x"51e8a43f",
          8529 => x"82d8c808",
          8530 => x"83ffff06",
          8531 => x"5677802e",
          8532 => x"96387381",
          8533 => x"fe2680c8",
          8534 => x"3873101a",
          8535 => x"76595375",
          8536 => x"73238114",
          8537 => x"548b3975",
          8538 => x"83ffff2e",
          8539 => x"098106b0",
          8540 => x"38811757",
          8541 => x"8c7727c1",
          8542 => x"38743370",
          8543 => x"862a7081",
          8544 => x"06515455",
          8545 => x"72802e8e",
          8546 => x"387381fe",
          8547 => x"26923873",
          8548 => x"101a5380",
          8549 => x"7323ff1c",
          8550 => x"7081ff06",
          8551 => x"51538439",
          8552 => x"81ff5372",
          8553 => x"5c9d397b",
          8554 => x"93387451",
          8555 => x"fce83f82",
          8556 => x"d8c80881",
          8557 => x"ff065372",
          8558 => x"7d2ea738",
          8559 => x"ff0bac1a",
          8560 => x"0ca03980",
          8561 => x"527851f8",
          8562 => x"d23f82d8",
          8563 => x"c8085b82",
          8564 => x"d8c80889",
          8565 => x"38981908",
          8566 => x"fd843886",
          8567 => x"39800b98",
          8568 => x"1a0c7a82",
          8569 => x"d8c80c90",
          8570 => x"3d0d04f2",
          8571 => x"3d0d6070",
          8572 => x"08405980",
          8573 => x"527851f6",
          8574 => x"d73f82d8",
          8575 => x"c8085882",
          8576 => x"d8c80883",
          8577 => x"a43881ff",
          8578 => x"705f5cff",
          8579 => x"0bac1a0c",
          8580 => x"98190852",
          8581 => x"7e51eaa9",
          8582 => x"3f82d8c8",
          8583 => x"085882d8",
          8584 => x"c8088385",
          8585 => x"389c1908",
          8586 => x"70335757",
          8587 => x"75863884",
          8588 => x"5882f639",
          8589 => x"8b1733bf",
          8590 => x"067081ff",
          8591 => x"06565473",
          8592 => x"861a3475",
          8593 => x"81e52e82",
          8594 => x"c3387483",
          8595 => x"2a708106",
          8596 => x"5154748f",
          8597 => x"2e8e3873",
          8598 => x"82b23874",
          8599 => x"8f2e0981",
          8600 => x"0681f738",
          8601 => x"ab193370",
          8602 => x"862a7081",
          8603 => x"06515555",
          8604 => x"7382a138",
          8605 => x"75862a70",
          8606 => x"81065154",
          8607 => x"73802e92",
          8608 => x"388d1733",
          8609 => x"7681bf06",
          8610 => x"70901c08",
          8611 => x"ac1d0c58",
          8612 => x"5d5e757c",
          8613 => x"2e098106",
          8614 => x"81b9388d",
          8615 => x"1733567d",
          8616 => x"762e0981",
          8617 => x"0681ac38",
          8618 => x"8c1f089a",
          8619 => x"18525de5",
          8620 => x"b63f82d8",
          8621 => x"c80883ff",
          8622 => x"ff065574",
          8623 => x"81953876",
          8624 => x"3370bf06",
          8625 => x"8d29f305",
          8626 => x"59568175",
          8627 => x"5c5a82ca",
          8628 => x"d01b3377",
          8629 => x"0551e58f",
          8630 => x"3f82d8c8",
          8631 => x"0883ffff",
          8632 => x"06567980",
          8633 => x"2eb13877",
          8634 => x"81fe2680",
          8635 => x"e6387551",
          8636 => x"80dfb43f",
          8637 => x"82d8c808",
          8638 => x"78101e70",
          8639 => x"22535581",
          8640 => x"19595580",
          8641 => x"dfa13f74",
          8642 => x"82d8c808",
          8643 => x"2e098106",
          8644 => x"80c13875",
          8645 => x"5a8b3975",
          8646 => x"83ffff2e",
          8647 => x"098106b3",
          8648 => x"38811b5b",
          8649 => x"8c7b27ff",
          8650 => x"a5387633",
          8651 => x"70862a70",
          8652 => x"81065155",
          8653 => x"5779802e",
          8654 => x"90387380",
          8655 => x"2e8b3877",
          8656 => x"101d7022",
          8657 => x"5154738b",
          8658 => x"38ff1c70",
          8659 => x"81ff0651",
          8660 => x"54843981",
          8661 => x"ff54735c",
          8662 => x"bb397b93",
          8663 => x"387651f9",
          8664 => x"b53f82d8",
          8665 => x"c80881ff",
          8666 => x"0654737e",
          8667 => x"2ebb38ab",
          8668 => x"19338106",
          8669 => x"54739538",
          8670 => x"8b53a019",
          8671 => x"529c1908",
          8672 => x"51e5b03f",
          8673 => x"82d8c808",
          8674 => x"802e9e38",
          8675 => x"81ff5cff",
          8676 => x"0bac1a0c",
          8677 => x"80527851",
          8678 => x"f5813f82",
          8679 => x"d8c80858",
          8680 => x"82d8c808",
          8681 => x"802efce8",
          8682 => x"387782d8",
          8683 => x"c80c903d",
          8684 => x"0d04ee3d",
          8685 => x"0d647008",
          8686 => x"ab123381",
          8687 => x"a006565d",
          8688 => x"5a865573",
          8689 => x"85b53873",
          8690 => x"8c1d0870",
          8691 => x"2256565d",
          8692 => x"73802e8d",
          8693 => x"38811d70",
          8694 => x"10167022",
          8695 => x"51555df0",
          8696 => x"398c53a0",
          8697 => x"1a705392",
          8698 => x"3d70535f",
          8699 => x"59e4873f",
          8700 => x"0280cb05",
          8701 => x"33810654",
          8702 => x"73802e82",
          8703 => x"a83880c0",
          8704 => x"0bab1b34",
          8705 => x"815b8c1c",
          8706 => x"087b5658",
          8707 => x"8b537d52",
          8708 => x"7851e3e2",
          8709 => x"3f857b27",
          8710 => x"80c6387a",
          8711 => x"56772270",
          8712 => x"83ffff06",
          8713 => x"55557380",
          8714 => x"2eb43874",
          8715 => x"83ffff06",
          8716 => x"82195955",
          8717 => x"8f577481",
          8718 => x"06761007",
          8719 => x"75812a71",
          8720 => x"902a7081",
          8721 => x"06515656",
          8722 => x"5673802e",
          8723 => x"87387584",
          8724 => x"a0a13256",
          8725 => x"ff175776",
          8726 => x"8025db38",
          8727 => x"c0397555",
          8728 => x"87028405",
          8729 => x"bf055757",
          8730 => x"74b007bf",
          8731 => x"0654b974",
          8732 => x"27843887",
          8733 => x"14547376",
          8734 => x"34ff16ff",
          8735 => x"1876842a",
          8736 => x"57585674",
          8737 => x"e338943d",
          8738 => x"ec051754",
          8739 => x"80fe7434",
          8740 => x"807727b5",
          8741 => x"38783354",
          8742 => x"73a02ead",
          8743 => x"38741970",
          8744 => x"335254e3",
          8745 => x"e03f82d8",
          8746 => x"c808802e",
          8747 => x"8c38ff17",
          8748 => x"5474742e",
          8749 => x"94388115",
          8750 => x"55811555",
          8751 => x"74772789",
          8752 => x"38741970",
          8753 => x"335154d0",
          8754 => x"39943d77",
          8755 => x"05eb0554",
          8756 => x"78158116",
          8757 => x"5658a056",
          8758 => x"7687268a",
          8759 => x"38811781",
          8760 => x"15703358",
          8761 => x"55577578",
          8762 => x"34877527",
          8763 => x"e3387951",
          8764 => x"f9f93f82",
          8765 => x"d8c8088b",
          8766 => x"38811b5b",
          8767 => x"80e37b27",
          8768 => x"fe843887",
          8769 => x"557a80e4",
          8770 => x"2e82f038",
          8771 => x"82d8c808",
          8772 => x"5582d8c8",
          8773 => x"08842e09",
          8774 => x"810682df",
          8775 => x"380280cb",
          8776 => x"0533ab1b",
          8777 => x"340280cb",
          8778 => x"05337081",
          8779 => x"2a708106",
          8780 => x"51555e81",
          8781 => x"5973802e",
          8782 => x"90388d52",
          8783 => x"8c1d51fe",
          8784 => x"f4c13f82",
          8785 => x"d8c80819",
          8786 => x"59785279",
          8787 => x"51f3c53f",
          8788 => x"82d8c808",
          8789 => x"5782d8c8",
          8790 => x"08829e38",
          8791 => x"ff195978",
          8792 => x"802e81d4",
          8793 => x"3878852b",
          8794 => x"901b0871",
          8795 => x"31535479",
          8796 => x"51efdd3f",
          8797 => x"82d8c808",
          8798 => x"5782d8c8",
          8799 => x"0881fa38",
          8800 => x"a01a51f5",
          8801 => x"913f82d8",
          8802 => x"c80881ff",
          8803 => x"065d981a",
          8804 => x"08527b51",
          8805 => x"e3ab3f82",
          8806 => x"d8c80857",
          8807 => x"82d8c808",
          8808 => x"81d7388c",
          8809 => x"1c089c1b",
          8810 => x"087a81ff",
          8811 => x"065a575b",
          8812 => x"7c8d1734",
          8813 => x"8f0b8b17",
          8814 => x"3482d8c8",
          8815 => x"088c1734",
          8816 => x"82d8c808",
          8817 => x"529a1651",
          8818 => x"dfdf3f77",
          8819 => x"8d29f305",
          8820 => x"77555573",
          8821 => x"83ffff2e",
          8822 => x"8b387410",
          8823 => x"1b702281",
          8824 => x"17575154",
          8825 => x"735282ca",
          8826 => x"d0173376",
          8827 => x"0551dfb9",
          8828 => x"3f738538",
          8829 => x"83ffff54",
          8830 => x"8117578c",
          8831 => x"7727d438",
          8832 => x"7383ffff",
          8833 => x"2e8b3874",
          8834 => x"101b7022",
          8835 => x"51547386",
          8836 => x"387780c0",
          8837 => x"07587776",
          8838 => x"34810b83",
          8839 => x"1d348052",
          8840 => x"7951eff7",
          8841 => x"3f82d8c8",
          8842 => x"085782d8",
          8843 => x"c80880c9",
          8844 => x"38ff1959",
          8845 => x"78fed738",
          8846 => x"981a0852",
          8847 => x"7b51e281",
          8848 => x"3f82d8c8",
          8849 => x"085782d8",
          8850 => x"c808ae38",
          8851 => x"a05382d8",
          8852 => x"c808529c",
          8853 => x"1a0851df",
          8854 => x"c03f8b53",
          8855 => x"a01a529c",
          8856 => x"1a0851df",
          8857 => x"913f9c1a",
          8858 => x"08ab1b33",
          8859 => x"98065555",
          8860 => x"738c1634",
          8861 => x"810b831d",
          8862 => x"34765574",
          8863 => x"82d8c80c",
          8864 => x"943d0d04",
          8865 => x"fa3d0d78",
          8866 => x"70089012",
          8867 => x"08ac1308",
          8868 => x"56595755",
          8869 => x"72ff2e94",
          8870 => x"38725274",
          8871 => x"51edb13f",
          8872 => x"82d8c808",
          8873 => x"5482d8c8",
          8874 => x"0880c938",
          8875 => x"98150852",
          8876 => x"7551e18d",
          8877 => x"3f82d8c8",
          8878 => x"085482d8",
          8879 => x"c808ab38",
          8880 => x"9c150853",
          8881 => x"e5733481",
          8882 => x"0b831734",
          8883 => x"90150877",
          8884 => x"27a23882",
          8885 => x"d8c80852",
          8886 => x"7451eebf",
          8887 => x"3f82d8c8",
          8888 => x"085482d8",
          8889 => x"c808802e",
          8890 => x"c3387384",
          8891 => x"2e098106",
          8892 => x"83388254",
          8893 => x"7382d8c8",
          8894 => x"0c883d0d",
          8895 => x"04f43d0d",
          8896 => x"7e607108",
          8897 => x"5f595c80",
          8898 => x"0b961934",
          8899 => x"981c0880",
          8900 => x"2e83e238",
          8901 => x"ac1c08ff",
          8902 => x"2e81bb38",
          8903 => x"8070717f",
          8904 => x"8c050870",
          8905 => x"2257575b",
          8906 => x"5c577277",
          8907 => x"2e819d38",
          8908 => x"78101470",
          8909 => x"22811b5b",
          8910 => x"56537a97",
          8911 => x"3880d080",
          8912 => x"157083ff",
          8913 => x"ff065153",
          8914 => x"728fff26",
          8915 => x"8638745b",
          8916 => x"80df3976",
          8917 => x"18961181",
          8918 => x"ff793158",
          8919 => x"5b5483b5",
          8920 => x"527a902b",
          8921 => x"75075180",
          8922 => x"d5983f82",
          8923 => x"d8c80883",
          8924 => x"ffff0655",
          8925 => x"81ff7527",
          8926 => x"95388176",
          8927 => x"27a53874",
          8928 => x"882a5372",
          8929 => x"7a347497",
          8930 => x"15348255",
          8931 => x"9f397430",
          8932 => x"76307078",
          8933 => x"07802572",
          8934 => x"80250752",
          8935 => x"54547380",
          8936 => x"2e853880",
          8937 => x"579a3974",
          8938 => x"7a348155",
          8939 => x"74175780",
          8940 => x"5b8c1d08",
          8941 => x"79101170",
          8942 => x"22515454",
          8943 => x"72fef138",
          8944 => x"7a307080",
          8945 => x"25703079",
          8946 => x"06595153",
          8947 => x"77179405",
          8948 => x"53800b82",
          8949 => x"14348070",
          8950 => x"891a585a",
          8951 => x"579c1c08",
          8952 => x"19703381",
          8953 => x"1b5b5653",
          8954 => x"74a02eb7",
          8955 => x"3874852e",
          8956 => x"09810684",
          8957 => x"3881e555",
          8958 => x"78893270",
          8959 => x"30707207",
          8960 => x"80255154",
          8961 => x"54768b26",
          8962 => x"90387280",
          8963 => x"2e8b38ae",
          8964 => x"76708105",
          8965 => x"58348117",
          8966 => x"57747670",
          8967 => x"81055834",
          8968 => x"8117578a",
          8969 => x"7927ffb5",
          8970 => x"38771788",
          8971 => x"0553800b",
          8972 => x"81143496",
          8973 => x"18335372",
          8974 => x"81873876",
          8975 => x"8b38bf0b",
          8976 => x"96193481",
          8977 => x"5780e139",
          8978 => x"7273891a",
          8979 => x"33555a57",
          8980 => x"72802e80",
          8981 => x"d3389618",
          8982 => x"89195556",
          8983 => x"7333ffbf",
          8984 => x"11545572",
          8985 => x"9926aa38",
          8986 => x"9c1c088c",
          8987 => x"11335153",
          8988 => x"88792787",
          8989 => x"3872842a",
          8990 => x"53853972",
          8991 => x"832a5372",
          8992 => x"81065372",
          8993 => x"802e8a38",
          8994 => x"a0157083",
          8995 => x"ffff0656",
          8996 => x"53747670",
          8997 => x"81055834",
          8998 => x"81198115",
          8999 => x"81197133",
          9000 => x"56595559",
          9001 => x"72ffb538",
          9002 => x"77179405",
          9003 => x"53800b82",
          9004 => x"14349c1c",
          9005 => x"088c1133",
          9006 => x"51537285",
          9007 => x"38728919",
          9008 => x"349c1c08",
          9009 => x"538b1333",
          9010 => x"8819349c",
          9011 => x"1c089c11",
          9012 => x"5253d9aa",
          9013 => x"3f82d8c8",
          9014 => x"08780c96",
          9015 => x"1351d987",
          9016 => x"3f82d8c8",
          9017 => x"08861923",
          9018 => x"981351d8",
          9019 => x"fa3f82d8",
          9020 => x"c8088419",
          9021 => x"238e3d0d",
          9022 => x"04f03d0d",
          9023 => x"62700841",
          9024 => x"5e806470",
          9025 => x"33515555",
          9026 => x"73af2e83",
          9027 => x"38815573",
          9028 => x"80dc2e92",
          9029 => x"3874802e",
          9030 => x"8d387f98",
          9031 => x"0508881f",
          9032 => x"0caa3981",
          9033 => x"15448064",
          9034 => x"70335656",
          9035 => x"5673af2e",
          9036 => x"09810683",
          9037 => x"38815673",
          9038 => x"80dc3270",
          9039 => x"30708025",
          9040 => x"78075151",
          9041 => x"5473dc38",
          9042 => x"73881f0c",
          9043 => x"63703351",
          9044 => x"54739f26",
          9045 => x"9638ff80",
          9046 => x"0bab1f34",
          9047 => x"80527d51",
          9048 => x"e7ee3f82",
          9049 => x"d8c80856",
          9050 => x"87e13963",
          9051 => x"417d088c",
          9052 => x"11085b54",
          9053 => x"8059923d",
          9054 => x"fc0551da",
          9055 => x"8f3f82d8",
          9056 => x"c808ff2e",
          9057 => x"82b13883",
          9058 => x"ffff0b82",
          9059 => x"d8c80827",
          9060 => x"92387810",
          9061 => x"1a82d8c8",
          9062 => x"08902a55",
          9063 => x"55737523",
          9064 => x"81195982",
          9065 => x"d8c80883",
          9066 => x"ffff0670",
          9067 => x"af327030",
          9068 => x"9f732771",
          9069 => x"80250751",
          9070 => x"51555673",
          9071 => x"b4387580",
          9072 => x"dc2eae38",
          9073 => x"7580ff26",
          9074 => x"91387552",
          9075 => x"82c9ec51",
          9076 => x"d9923f82",
          9077 => x"d8c80881",
          9078 => x"de387881",
          9079 => x"fe2681d7",
          9080 => x"3878101a",
          9081 => x"54757423",
          9082 => x"811959ff",
          9083 => x"89398115",
          9084 => x"41806170",
          9085 => x"33565657",
          9086 => x"73af2e09",
          9087 => x"81068338",
          9088 => x"81577380",
          9089 => x"dc327030",
          9090 => x"70802579",
          9091 => x"07515154",
          9092 => x"73dc3874",
          9093 => x"449f7627",
          9094 => x"822b5778",
          9095 => x"812e0981",
          9096 => x"068c3879",
          9097 => x"225473ae",
          9098 => x"2ea53880",
          9099 => x"d2397882",
          9100 => x"2e098106",
          9101 => x"80c93882",
          9102 => x"1a225473",
          9103 => x"ae2e0981",
          9104 => x"0680c138",
          9105 => x"79225473",
          9106 => x"ae2e0981",
          9107 => x"06b63878",
          9108 => x"101a5480",
          9109 => x"7423800b",
          9110 => x"a01f5658",
          9111 => x"ae547878",
          9112 => x"268338a0",
          9113 => x"54737570",
          9114 => x"81055734",
          9115 => x"8118588a",
          9116 => x"7827e938",
          9117 => x"76a00754",
          9118 => x"73ab1f34",
          9119 => x"84c43978",
          9120 => x"802ea838",
          9121 => x"78101afe",
          9122 => x"05557422",
          9123 => x"fe167172",
          9124 => x"a0327030",
          9125 => x"709f2a51",
          9126 => x"51535856",
          9127 => x"5475ae2e",
          9128 => x"84387387",
          9129 => x"38ff1959",
          9130 => x"78e03878",
          9131 => x"197a1155",
          9132 => x"56807423",
          9133 => x"788d3886",
          9134 => x"56859039",
          9135 => x"76830757",
          9136 => x"83993980",
          9137 => x"7a227083",
          9138 => x"ffff0656",
          9139 => x"565d73a0",
          9140 => x"2e098106",
          9141 => x"9338811d",
          9142 => x"70101b70",
          9143 => x"2251555d",
          9144 => x"73a02ef2",
          9145 => x"387c8f38",
          9146 => x"7483ffff",
          9147 => x"065473ae",
          9148 => x"2e098106",
          9149 => x"85387683",
          9150 => x"07577880",
          9151 => x"2eaa3879",
          9152 => x"16fe0570",
          9153 => x"22515473",
          9154 => x"ae2e9d38",
          9155 => x"78101afe",
          9156 => x"0555ff19",
          9157 => x"5978802e",
          9158 => x"8f38fe15",
          9159 => x"70225555",
          9160 => x"73ae2e09",
          9161 => x"8106eb38",
          9162 => x"8b53a052",
          9163 => x"a01e51d5",
          9164 => x"e83f8070",
          9165 => x"595c885f",
          9166 => x"7c101a70",
          9167 => x"22811f5f",
          9168 => x"57547580",
          9169 => x"2e829438",
          9170 => x"75a02e96",
          9171 => x"3875ae32",
          9172 => x"70307080",
          9173 => x"25515154",
          9174 => x"7c792e8c",
          9175 => x"3873802e",
          9176 => x"89387683",
          9177 => x"0757d139",
          9178 => x"8054735b",
          9179 => x"7e782683",
          9180 => x"38815b7c",
          9181 => x"79327030",
          9182 => x"70720780",
          9183 => x"25707e07",
          9184 => x"51515555",
          9185 => x"73802ea6",
          9186 => x"387e8b2e",
          9187 => x"feae387c",
          9188 => x"792e8b38",
          9189 => x"76830757",
          9190 => x"7c792681",
          9191 => x"be38785d",
          9192 => x"88588b7c",
          9193 => x"822b81fc",
          9194 => x"065d5fff",
          9195 => x"8b3980ff",
          9196 => x"7627af38",
          9197 => x"76820757",
          9198 => x"83b55275",
          9199 => x"5180ccc2",
          9200 => x"3f82d8c8",
          9201 => x"0883ffff",
          9202 => x"0670872a",
          9203 => x"70810651",
          9204 => x"55567380",
          9205 => x"2e8c3875",
          9206 => x"80ff0682",
          9207 => x"cae01133",
          9208 => x"575481ff",
          9209 => x"7627a438",
          9210 => x"ff1f5473",
          9211 => x"78268a38",
          9212 => x"7683077f",
          9213 => x"5957fec0",
          9214 => x"397d18a0",
          9215 => x"0576882a",
          9216 => x"55557375",
          9217 => x"34811858",
          9218 => x"80c33975",
          9219 => x"802e9238",
          9220 => x"755282c9",
          9221 => x"f851d4cc",
          9222 => x"3f82d8c8",
          9223 => x"08802e8a",
          9224 => x"3880df77",
          9225 => x"83075856",
          9226 => x"a439ffbf",
          9227 => x"16547399",
          9228 => x"2685387b",
          9229 => x"82075cff",
          9230 => x"9f165473",
          9231 => x"99268e38",
          9232 => x"7b8107e0",
          9233 => x"177083ff",
          9234 => x"ff065855",
          9235 => x"5c7d18a0",
          9236 => x"05547574",
          9237 => x"34811858",
          9238 => x"fdde39a0",
          9239 => x"1e335473",
          9240 => x"81e52e09",
          9241 => x"81068638",
          9242 => x"850ba01f",
          9243 => x"347e882e",
          9244 => x"09810688",
          9245 => x"387b822b",
          9246 => x"81fc065c",
          9247 => x"7b8c0654",
          9248 => x"738c2e8d",
          9249 => x"387b8306",
          9250 => x"5473832e",
          9251 => x"09810685",
          9252 => x"38768207",
          9253 => x"5776812a",
          9254 => x"70810651",
          9255 => x"54739f38",
          9256 => x"7b810654",
          9257 => x"73802e85",
          9258 => x"38769007",
          9259 => x"577b822a",
          9260 => x"70810651",
          9261 => x"5473802e",
          9262 => x"85387688",
          9263 => x"075776ab",
          9264 => x"1f347d51",
          9265 => x"eaa53f82",
          9266 => x"d8c808ab",
          9267 => x"1f335656",
          9268 => x"82d8c808",
          9269 => x"802ebe38",
          9270 => x"82d8c808",
          9271 => x"842e0981",
          9272 => x"0680e838",
          9273 => x"74852a70",
          9274 => x"81067682",
          9275 => x"2a575154",
          9276 => x"73802e96",
          9277 => x"38748106",
          9278 => x"5473802e",
          9279 => x"f8ed38ff",
          9280 => x"800bab1f",
          9281 => x"34805680",
          9282 => x"c2397481",
          9283 => x"065473bb",
          9284 => x"388556b7",
          9285 => x"3974822a",
          9286 => x"70810651",
          9287 => x"5473ac38",
          9288 => x"861e3370",
          9289 => x"842a7081",
          9290 => x"06515555",
          9291 => x"73802ee1",
          9292 => x"38901e08",
          9293 => x"83ff0660",
          9294 => x"05b80552",
          9295 => x"7f51e4ef",
          9296 => x"3f82d8c8",
          9297 => x"08881f0c",
          9298 => x"f8a13975",
          9299 => x"82d8c80c",
          9300 => x"923d0d04",
          9301 => x"f63d0d7c",
          9302 => x"5bff7b08",
          9303 => x"70717355",
          9304 => x"595c5559",
          9305 => x"73802e81",
          9306 => x"c6387570",
          9307 => x"81055733",
          9308 => x"709f2652",
          9309 => x"5271ba2e",
          9310 => x"8d3870ee",
          9311 => x"3871ba2e",
          9312 => x"09810681",
          9313 => x"a5387333",
          9314 => x"d0117081",
          9315 => x"ff065152",
          9316 => x"53708926",
          9317 => x"91388214",
          9318 => x"7381ff06",
          9319 => x"d0055652",
          9320 => x"71762e80",
          9321 => x"f738800b",
          9322 => x"82cac059",
          9323 => x"5577087a",
          9324 => x"55577670",
          9325 => x"81055833",
          9326 => x"74708105",
          9327 => x"5633ff9f",
          9328 => x"12535353",
          9329 => x"70992689",
          9330 => x"38e01370",
          9331 => x"81ff0654",
          9332 => x"51ff9f12",
          9333 => x"51709926",
          9334 => x"8938e012",
          9335 => x"7081ff06",
          9336 => x"53517230",
          9337 => x"709f2a51",
          9338 => x"5172722e",
          9339 => x"09810685",
          9340 => x"3870ffbe",
          9341 => x"38723074",
          9342 => x"77327030",
          9343 => x"7072079f",
          9344 => x"2a739f2a",
          9345 => x"07535454",
          9346 => x"5170802e",
          9347 => x"8f388115",
          9348 => x"84195955",
          9349 => x"837525ff",
          9350 => x"94388b39",
          9351 => x"74832486",
          9352 => x"3874767c",
          9353 => x"0c597851",
          9354 => x"863982f0",
          9355 => x"a4335170",
          9356 => x"82d8c80c",
          9357 => x"8c3d0d04",
          9358 => x"fa3d0d78",
          9359 => x"56800b83",
          9360 => x"1734ff0b",
          9361 => x"b4170c79",
          9362 => x"527551d1",
          9363 => x"f43f8455",
          9364 => x"82d8c808",
          9365 => x"81803884",
          9366 => x"b61651ce",
          9367 => x"8a3f82d8",
          9368 => x"c80883ff",
          9369 => x"ff065483",
          9370 => x"557382d4",
          9371 => x"d52e0981",
          9372 => x"0680e338",
          9373 => x"800bb817",
          9374 => x"33565774",
          9375 => x"81e92e09",
          9376 => x"81068338",
          9377 => x"81577481",
          9378 => x"eb327030",
          9379 => x"70802579",
          9380 => x"07515154",
          9381 => x"738a3874",
          9382 => x"81e82e09",
          9383 => x"8106b538",
          9384 => x"835382ca",
          9385 => x"805280ee",
          9386 => x"1651cf87",
          9387 => x"3f82d8c8",
          9388 => x"085582d8",
          9389 => x"c808802e",
          9390 => x"9d388553",
          9391 => x"82ca8452",
          9392 => x"818a1651",
          9393 => x"ceed3f82",
          9394 => x"d8c80855",
          9395 => x"82d8c808",
          9396 => x"802e8338",
          9397 => x"82557482",
          9398 => x"d8c80c88",
          9399 => x"3d0d04f2",
          9400 => x"3d0d6102",
          9401 => x"840580cb",
          9402 => x"05335855",
          9403 => x"80750c60",
          9404 => x"51fce13f",
          9405 => x"82d8c808",
          9406 => x"588b5680",
          9407 => x"0b82d8c8",
          9408 => x"08248784",
          9409 => x"3882d8c8",
          9410 => x"08842982",
          9411 => x"f0900570",
          9412 => x"0855538c",
          9413 => x"5673802e",
          9414 => x"86ee3873",
          9415 => x"750c7681",
          9416 => x"fe067433",
          9417 => x"54577280",
          9418 => x"2eae3881",
          9419 => x"143351c6",
          9420 => x"a03f82d8",
          9421 => x"c80881ff",
          9422 => x"06708106",
          9423 => x"54557298",
          9424 => x"3876802e",
          9425 => x"86c03874",
          9426 => x"822a7081",
          9427 => x"0651538a",
          9428 => x"567286b4",
          9429 => x"3886af39",
          9430 => x"80743477",
          9431 => x"81153481",
          9432 => x"52811433",
          9433 => x"51c6883f",
          9434 => x"82d8c808",
          9435 => x"81ff0670",
          9436 => x"81065455",
          9437 => x"83567286",
          9438 => x"8f387680",
          9439 => x"2e8f3874",
          9440 => x"822a7081",
          9441 => x"0651538a",
          9442 => x"567285fc",
          9443 => x"38807053",
          9444 => x"74525bfd",
          9445 => x"a33f82d8",
          9446 => x"c80881ff",
          9447 => x"06577682",
          9448 => x"2e098106",
          9449 => x"80e2388c",
          9450 => x"3d745658",
          9451 => x"835683fa",
          9452 => x"15337058",
          9453 => x"5372802e",
          9454 => x"8d3883fe",
          9455 => x"1551cbbe",
          9456 => x"3f82d8c8",
          9457 => x"08577678",
          9458 => x"7084055a",
          9459 => x"0cff1690",
          9460 => x"16565675",
          9461 => x"8025d738",
          9462 => x"800b8d3d",
          9463 => x"54567270",
          9464 => x"84055408",
          9465 => x"5b83577a",
          9466 => x"802e9538",
          9467 => x"7a527351",
          9468 => x"fcc63f82",
          9469 => x"d8c80881",
          9470 => x"ff065781",
          9471 => x"77278938",
          9472 => x"81165683",
          9473 => x"7627d738",
          9474 => x"81567684",
          9475 => x"2e84f938",
          9476 => x"8d567681",
          9477 => x"2684f138",
          9478 => x"80c31451",
          9479 => x"cac93f82",
          9480 => x"d8c80883",
          9481 => x"ffff0653",
          9482 => x"7284802e",
          9483 => x"09810684",
          9484 => x"d73880ce",
          9485 => x"1451caaf",
          9486 => x"3f82d8c8",
          9487 => x"0883ffff",
          9488 => x"0658778d",
          9489 => x"3880dc14",
          9490 => x"51cab33f",
          9491 => x"82d8c808",
          9492 => x"5877a015",
          9493 => x"0c80c814",
          9494 => x"33821534",
          9495 => x"80c81433",
          9496 => x"ff117081",
          9497 => x"ff065154",
          9498 => x"558d5672",
          9499 => x"81268498",
          9500 => x"387481ff",
          9501 => x"06787129",
          9502 => x"80c51633",
          9503 => x"52595372",
          9504 => x"8a152372",
          9505 => x"802e8b38",
          9506 => x"ff137306",
          9507 => x"5372802e",
          9508 => x"86388d56",
          9509 => x"83f23980",
          9510 => x"c91451c9",
          9511 => x"ca3f82d8",
          9512 => x"c8085382",
          9513 => x"d8c80888",
          9514 => x"1523728f",
          9515 => x"06578d56",
          9516 => x"7683d538",
          9517 => x"80cb1451",
          9518 => x"c9ad3f82",
          9519 => x"d8c80883",
          9520 => x"ffff0655",
          9521 => x"748d3880",
          9522 => x"d81451c9",
          9523 => x"b13f82d8",
          9524 => x"c8085580",
          9525 => x"c61451c9",
          9526 => x"8e3f82d8",
          9527 => x"c80883ff",
          9528 => x"ff06538d",
          9529 => x"5672802e",
          9530 => x"839e3888",
          9531 => x"14227814",
          9532 => x"71842a05",
          9533 => x"5a5a7875",
          9534 => x"26838d38",
          9535 => x"8a142252",
          9536 => x"74793151",
          9537 => x"fedcfc3f",
          9538 => x"82d8c808",
          9539 => x"5582d8c8",
          9540 => x"08802e82",
          9541 => x"f33882d8",
          9542 => x"c80880ff",
          9543 => x"fffff526",
          9544 => x"83388357",
          9545 => x"7483fff5",
          9546 => x"26833882",
          9547 => x"57749ff5",
          9548 => x"26853881",
          9549 => x"5789398d",
          9550 => x"5676802e",
          9551 => x"82ca3882",
          9552 => x"15709c16",
          9553 => x"0c7ba416",
          9554 => x"0c731c70",
          9555 => x"a8170c7a",
          9556 => x"1db0170c",
          9557 => x"54557683",
          9558 => x"2e098106",
          9559 => x"af3880e2",
          9560 => x"1451c883",
          9561 => x"3f82d8c8",
          9562 => x"0883ffff",
          9563 => x"06538d56",
          9564 => x"72829538",
          9565 => x"79829138",
          9566 => x"80e41451",
          9567 => x"c8803f82",
          9568 => x"d8c808ac",
          9569 => x"150c7482",
          9570 => x"2b53a239",
          9571 => x"8d567980",
          9572 => x"2e81f538",
          9573 => x"7713ac15",
          9574 => x"0c741553",
          9575 => x"76822e8d",
          9576 => x"38741015",
          9577 => x"70812a76",
          9578 => x"81060551",
          9579 => x"5383ff13",
          9580 => x"892a538d",
          9581 => x"5672a015",
          9582 => x"082681cc",
          9583 => x"38ff0b94",
          9584 => x"150cff0b",
          9585 => x"90150cff",
          9586 => x"800b8415",
          9587 => x"3476832e",
          9588 => x"09810681",
          9589 => x"923880e8",
          9590 => x"1451c78b",
          9591 => x"3f82d8c8",
          9592 => x"0883ffff",
          9593 => x"06537281",
          9594 => x"2e098106",
          9595 => x"80f93881",
          9596 => x"1b527351",
          9597 => x"cacb3f82",
          9598 => x"d8c80880",
          9599 => x"ea3882d8",
          9600 => x"c8088415",
          9601 => x"3484b614",
          9602 => x"51c6dc3f",
          9603 => x"82d8c808",
          9604 => x"83ffff06",
          9605 => x"537282d4",
          9606 => x"d52e0981",
          9607 => x"0680c838",
          9608 => x"b81451c6",
          9609 => x"d93f82d8",
          9610 => x"c808848b",
          9611 => x"85a4d22e",
          9612 => x"098106b3",
          9613 => x"38849c14",
          9614 => x"51c6c33f",
          9615 => x"82d8c808",
          9616 => x"868a85e4",
          9617 => x"f22e0981",
          9618 => x"069d3884",
          9619 => x"a01451c6",
          9620 => x"ad3f82d8",
          9621 => x"c8089415",
          9622 => x"0c84a414",
          9623 => x"51c69f3f",
          9624 => x"82d8c808",
          9625 => x"90150c76",
          9626 => x"743482f0",
          9627 => x"a0228105",
          9628 => x"537282f0",
          9629 => x"a0237286",
          9630 => x"152382f0",
          9631 => x"a80b8c15",
          9632 => x"0c800b98",
          9633 => x"150c8056",
          9634 => x"7582d8c8",
          9635 => x"0c903d0d",
          9636 => x"04fb3d0d",
          9637 => x"77548955",
          9638 => x"73802eba",
          9639 => x"38730853",
          9640 => x"72802eb2",
          9641 => x"38723352",
          9642 => x"71802eaa",
          9643 => x"38861322",
          9644 => x"84152257",
          9645 => x"5271762e",
          9646 => x"0981069a",
          9647 => x"38811333",
          9648 => x"51ffbf8d",
          9649 => x"3f82d8c8",
          9650 => x"08810652",
          9651 => x"71883871",
          9652 => x"74085455",
          9653 => x"83398053",
          9654 => x"7873710c",
          9655 => x"527482d8",
          9656 => x"c80c873d",
          9657 => x"0d04fa3d",
          9658 => x"0d02ab05",
          9659 => x"337a5889",
          9660 => x"3dfc0552",
          9661 => x"56f4dd3f",
          9662 => x"8b54800b",
          9663 => x"82d8c808",
          9664 => x"24bc3882",
          9665 => x"d8c80884",
          9666 => x"2982f090",
          9667 => x"05700855",
          9668 => x"5573802e",
          9669 => x"84388074",
          9670 => x"34785473",
          9671 => x"802e8438",
          9672 => x"80743478",
          9673 => x"750c7554",
          9674 => x"75802e92",
          9675 => x"38805389",
          9676 => x"3d705384",
          9677 => x"0551f7a7",
          9678 => x"3f82d8c8",
          9679 => x"08547382",
          9680 => x"d8c80c88",
          9681 => x"3d0d04ea",
          9682 => x"3d0d6802",
          9683 => x"840580eb",
          9684 => x"05335959",
          9685 => x"89547880",
          9686 => x"2e84c838",
          9687 => x"77bf0670",
          9688 => x"54993dcc",
          9689 => x"05539a3d",
          9690 => x"84055258",
          9691 => x"f6f13f82",
          9692 => x"d8c80855",
          9693 => x"82d8c808",
          9694 => x"84a4387a",
          9695 => x"5c69528c",
          9696 => x"3d705256",
          9697 => x"eaf33f82",
          9698 => x"d8c80855",
          9699 => x"82d8c808",
          9700 => x"92380280",
          9701 => x"d7053370",
          9702 => x"982b5557",
          9703 => x"73802583",
          9704 => x"38865577",
          9705 => x"9c065473",
          9706 => x"802e81ab",
          9707 => x"3874802e",
          9708 => x"95387484",
          9709 => x"2e098106",
          9710 => x"aa387551",
          9711 => x"dff43f82",
          9712 => x"d8c80855",
          9713 => x"9e3902b2",
          9714 => x"05339106",
          9715 => x"547381b8",
          9716 => x"3877822a",
          9717 => x"70810651",
          9718 => x"5473802e",
          9719 => x"8e388855",
          9720 => x"83bc3977",
          9721 => x"88075874",
          9722 => x"83b43877",
          9723 => x"832a7081",
          9724 => x"06515473",
          9725 => x"802e81af",
          9726 => x"3862527a",
          9727 => x"51d7b03f",
          9728 => x"82d8c808",
          9729 => x"568288b2",
          9730 => x"0a52628e",
          9731 => x"0551c3b7",
          9732 => x"3f6254a0",
          9733 => x"0b8b1534",
          9734 => x"80536252",
          9735 => x"7a51d7c8",
          9736 => x"3f805262",
          9737 => x"9c0551c3",
          9738 => x"9e3f7a54",
          9739 => x"810b8315",
          9740 => x"3475802e",
          9741 => x"80f1387a",
          9742 => x"b4110851",
          9743 => x"54805375",
          9744 => x"52983dd0",
          9745 => x"0551ccc9",
          9746 => x"3f82d8c8",
          9747 => x"085582d8",
          9748 => x"c80882ca",
          9749 => x"38b73974",
          9750 => x"82c43802",
          9751 => x"b2053370",
          9752 => x"842a7081",
          9753 => x"06515556",
          9754 => x"73802e86",
          9755 => x"38845582",
          9756 => x"ad397781",
          9757 => x"2a708106",
          9758 => x"51547380",
          9759 => x"2ea93875",
          9760 => x"81065473",
          9761 => x"802ea038",
          9762 => x"87558292",
          9763 => x"3973527a",
          9764 => x"51c5ae3f",
          9765 => x"82d8c808",
          9766 => x"7bff1890",
          9767 => x"120c5555",
          9768 => x"82d8c808",
          9769 => x"81f83877",
          9770 => x"832a7081",
          9771 => x"06515473",
          9772 => x"802e8638",
          9773 => x"7780c007",
          9774 => x"587ab411",
          9775 => x"08a01b0c",
          9776 => x"63a41b0c",
          9777 => x"63537052",
          9778 => x"57d5e43f",
          9779 => x"82d8c808",
          9780 => x"82d8c808",
          9781 => x"881b0c63",
          9782 => x"9c05525a",
          9783 => x"c1a03f82",
          9784 => x"d8c80882",
          9785 => x"d8c8088c",
          9786 => x"1b0c777a",
          9787 => x"0c568617",
          9788 => x"22841a23",
          9789 => x"77901a34",
          9790 => x"800b911a",
          9791 => x"34800b9c",
          9792 => x"1a0c800b",
          9793 => x"941a0c77",
          9794 => x"852a7081",
          9795 => x"06515473",
          9796 => x"802e818d",
          9797 => x"3882d8c8",
          9798 => x"08802e81",
          9799 => x"843882d8",
          9800 => x"c808941a",
          9801 => x"0c8a1722",
          9802 => x"70892b7b",
          9803 => x"525957a8",
          9804 => x"39765278",
          9805 => x"51c6aa3f",
          9806 => x"82d8c808",
          9807 => x"5782d8c8",
          9808 => x"08812683",
          9809 => x"38825582",
          9810 => x"d8c808ff",
          9811 => x"2e098106",
          9812 => x"83387955",
          9813 => x"75783156",
          9814 => x"74307076",
          9815 => x"07802551",
          9816 => x"54777627",
          9817 => x"8a388170",
          9818 => x"7506555a",
          9819 => x"73c33876",
          9820 => x"981a0c74",
          9821 => x"a9387583",
          9822 => x"ff065473",
          9823 => x"802ea238",
          9824 => x"76527a51",
          9825 => x"c5b13f82",
          9826 => x"d8c80885",
          9827 => x"3882558e",
          9828 => x"3975892a",
          9829 => x"82d8c808",
          9830 => x"059c1a0c",
          9831 => x"84398079",
          9832 => x"0c745473",
          9833 => x"82d8c80c",
          9834 => x"983d0d04",
          9835 => x"f23d0d60",
          9836 => x"63656440",
          9837 => x"405d5980",
          9838 => x"7e0c903d",
          9839 => x"fc055278",
          9840 => x"51f9ce3f",
          9841 => x"82d8c808",
          9842 => x"5582d8c8",
          9843 => x"088a3891",
          9844 => x"19335574",
          9845 => x"802e8638",
          9846 => x"745682c7",
          9847 => x"39901933",
          9848 => x"81065587",
          9849 => x"5674802e",
          9850 => x"82b93895",
          9851 => x"39820b91",
          9852 => x"1a348256",
          9853 => x"82ad3981",
          9854 => x"0b911a34",
          9855 => x"815682a3",
          9856 => x"398c1908",
          9857 => x"941a0831",
          9858 => x"55747c27",
          9859 => x"8338745c",
          9860 => x"7b802e82",
          9861 => x"8c389419",
          9862 => x"087083ff",
          9863 => x"06565674",
          9864 => x"81b4387e",
          9865 => x"8a1122ff",
          9866 => x"0577892a",
          9867 => x"065b5579",
          9868 => x"a8387587",
          9869 => x"38881908",
          9870 => x"558f3998",
          9871 => x"19085278",
          9872 => x"51c49e3f",
          9873 => x"82d8c808",
          9874 => x"55817527",
          9875 => x"ff9f3874",
          9876 => x"ff2effa3",
          9877 => x"3874981a",
          9878 => x"0c981908",
          9879 => x"527e51c3",
          9880 => x"d63f82d8",
          9881 => x"c808802e",
          9882 => x"ff833882",
          9883 => x"d8c8081a",
          9884 => x"7c892a59",
          9885 => x"5777802e",
          9886 => x"80d83877",
          9887 => x"1a7f8a11",
          9888 => x"22585c55",
          9889 => x"75752785",
          9890 => x"38757a31",
          9891 => x"58775476",
          9892 => x"537c5281",
          9893 => x"1b3351ff",
          9894 => x"b8d43f82",
          9895 => x"d8c808fe",
          9896 => x"d6387e83",
          9897 => x"11335656",
          9898 => x"74802ea0",
          9899 => x"38b41608",
          9900 => x"77315574",
          9901 => x"78279538",
          9902 => x"848053b8",
          9903 => x"1652b416",
          9904 => x"08773189",
          9905 => x"2b7d0551",
          9906 => x"ffbeab3f",
          9907 => x"77892b56",
          9908 => x"ba39769c",
          9909 => x"1a0c9419",
          9910 => x"0883ff06",
          9911 => x"84807131",
          9912 => x"57557b76",
          9913 => x"2783387b",
          9914 => x"569c1908",
          9915 => x"527e51c0",
          9916 => x"d03f82d8",
          9917 => x"c808fdff",
          9918 => x"38755394",
          9919 => x"190883ff",
          9920 => x"061fb805",
          9921 => x"527c51ff",
          9922 => x"bdec3f7b",
          9923 => x"76317e08",
          9924 => x"177f0c76",
          9925 => x"1e941b08",
          9926 => x"18941c0c",
          9927 => x"5e5cfdf0",
          9928 => x"39805675",
          9929 => x"82d8c80c",
          9930 => x"903d0d04",
          9931 => x"f23d0d60",
          9932 => x"63656440",
          9933 => x"405d5880",
          9934 => x"7e0c903d",
          9935 => x"fc055277",
          9936 => x"51f6ce3f",
          9937 => x"82d8c808",
          9938 => x"5582d8c8",
          9939 => x"088a3891",
          9940 => x"18335574",
          9941 => x"802e8638",
          9942 => x"745683be",
          9943 => x"39901833",
          9944 => x"70812a70",
          9945 => x"81065156",
          9946 => x"56875674",
          9947 => x"802e83aa",
          9948 => x"38953982",
          9949 => x"0b911934",
          9950 => x"8256839e",
          9951 => x"39810b91",
          9952 => x"19348156",
          9953 => x"83943994",
          9954 => x"18087c11",
          9955 => x"56567476",
          9956 => x"27843875",
          9957 => x"095c7b80",
          9958 => x"2e82f238",
          9959 => x"94180870",
          9960 => x"83ff0656",
          9961 => x"56748281",
          9962 => x"387e8a11",
          9963 => x"22ff0577",
          9964 => x"892a065c",
          9965 => x"557abf38",
          9966 => x"758c3888",
          9967 => x"18085574",
          9968 => x"9c387a52",
          9969 => x"85399818",
          9970 => x"08527751",
          9971 => x"c6ef3f82",
          9972 => x"d8c80855",
          9973 => x"82d8c808",
          9974 => x"802e82b1",
          9975 => x"3874812e",
          9976 => x"ff913874",
          9977 => x"ff2eff95",
          9978 => x"38749819",
          9979 => x"0c881808",
          9980 => x"85387488",
          9981 => x"190c7e55",
          9982 => x"b415089c",
          9983 => x"19082e09",
          9984 => x"81068e38",
          9985 => x"7451ffbd",
          9986 => x"c83f82d8",
          9987 => x"c808feed",
          9988 => x"38981808",
          9989 => x"527e51c0",
          9990 => x"9e3f82d8",
          9991 => x"c808802e",
          9992 => x"fed13882",
          9993 => x"d8c8081b",
          9994 => x"7c892a5a",
          9995 => x"5778802e",
          9996 => x"80d73878",
          9997 => x"1b7f8a11",
          9998 => x"22585b55",
          9999 => x"75752785",
         10000 => x"38757b31",
         10001 => x"59785476",
         10002 => x"537c5281",
         10003 => x"1a3351ff",
         10004 => x"b7863f82",
         10005 => x"d8c808fe",
         10006 => x"a4387eb4",
         10007 => x"11087831",
         10008 => x"56567479",
         10009 => x"279c3884",
         10010 => x"8053b416",
         10011 => x"08773189",
         10012 => x"2b7d0552",
         10013 => x"b81651ff",
         10014 => x"bafc3f7e",
         10015 => x"55800b83",
         10016 => x"16347889",
         10017 => x"2b5680de",
         10018 => x"398c1808",
         10019 => x"94190826",
         10020 => x"94387e51",
         10021 => x"ffbcba3f",
         10022 => x"82d8c808",
         10023 => x"fddf387e",
         10024 => x"77b4120c",
         10025 => x"55769c19",
         10026 => x"0c941808",
         10027 => x"83ff0684",
         10028 => x"80713157",
         10029 => x"557b7627",
         10030 => x"83387b56",
         10031 => x"9c180852",
         10032 => x"7e51ffbc",
         10033 => x"fc3f82d8",
         10034 => x"c808fdb1",
         10035 => x"3875537c",
         10036 => x"52941808",
         10037 => x"83ff061f",
         10038 => x"b80551ff",
         10039 => x"ba983f7e",
         10040 => x"55810b83",
         10041 => x"16347b76",
         10042 => x"317e0817",
         10043 => x"7f0c761e",
         10044 => x"941a0818",
         10045 => x"70941c0c",
         10046 => x"8c1b0858",
         10047 => x"585e5c74",
         10048 => x"76278338",
         10049 => x"7555748c",
         10050 => x"190cfd8a",
         10051 => x"39901833",
         10052 => x"80c00755",
         10053 => x"74901934",
         10054 => x"80567582",
         10055 => x"d8c80c90",
         10056 => x"3d0d04f8",
         10057 => x"3d0d7a8b",
         10058 => x"3dfc0553",
         10059 => x"705256f2",
         10060 => x"e03f82d8",
         10061 => x"c8085782",
         10062 => x"d8c80881",
         10063 => x"80389016",
         10064 => x"3370862a",
         10065 => x"70810651",
         10066 => x"55557380",
         10067 => x"2e80ee38",
         10068 => x"a0160852",
         10069 => x"7851ffbb",
         10070 => x"e83f82d8",
         10071 => x"c8085782",
         10072 => x"d8c80880",
         10073 => x"d838a416",
         10074 => x"088b1133",
         10075 => x"a0075555",
         10076 => x"738b1634",
         10077 => x"88160853",
         10078 => x"74527508",
         10079 => x"51cce93f",
         10080 => x"8c160852",
         10081 => x"9c1551ff",
         10082 => x"b8bd3f82",
         10083 => x"88b20a52",
         10084 => x"961551ff",
         10085 => x"b8b13f76",
         10086 => x"52921551",
         10087 => x"ffb88a3f",
         10088 => x"7854810b",
         10089 => x"83153478",
         10090 => x"51ffbbdc",
         10091 => x"3f82d8c8",
         10092 => x"08901733",
         10093 => x"81bf0655",
         10094 => x"57739017",
         10095 => x"347682d8",
         10096 => x"c80c8a3d",
         10097 => x"0d04fc3d",
         10098 => x"0d767052",
         10099 => x"54fed43f",
         10100 => x"82d8c808",
         10101 => x"5382d8c8",
         10102 => x"089c3886",
         10103 => x"3dfc0552",
         10104 => x"7351f1ad",
         10105 => x"3f82d8c8",
         10106 => x"085382d8",
         10107 => x"c8088738",
         10108 => x"82d8c808",
         10109 => x"740c7282",
         10110 => x"d8c80c86",
         10111 => x"3d0d04ff",
         10112 => x"3d0d843d",
         10113 => x"51e6cd3f",
         10114 => x"8b52800b",
         10115 => x"82d8c808",
         10116 => x"248b3882",
         10117 => x"d8c80882",
         10118 => x"f0a43480",
         10119 => x"527182d8",
         10120 => x"c80c833d",
         10121 => x"0d04ee3d",
         10122 => x"0d805394",
         10123 => x"3dcc0552",
         10124 => x"953d51e9",
         10125 => x"aa3f82d8",
         10126 => x"c8085582",
         10127 => x"d8c80880",
         10128 => x"e0387658",
         10129 => x"6452943d",
         10130 => x"d00551dd",
         10131 => x"ac3f82d8",
         10132 => x"c8085582",
         10133 => x"d8c808bc",
         10134 => x"380280c7",
         10135 => x"05337098",
         10136 => x"2b555673",
         10137 => x"80258938",
         10138 => x"767a9812",
         10139 => x"0c54b239",
         10140 => x"02a20533",
         10141 => x"70842a70",
         10142 => x"81065155",
         10143 => x"5673802e",
         10144 => x"9e38767f",
         10145 => x"53705254",
         10146 => x"caa53f82",
         10147 => x"d8c80898",
         10148 => x"150c8e39",
         10149 => x"82d8c808",
         10150 => x"842e0981",
         10151 => x"06833885",
         10152 => x"557482d8",
         10153 => x"c80c943d",
         10154 => x"0d04ffa3",
         10155 => x"3d0d80e1",
         10156 => x"3d0880e1",
         10157 => x"3d085b5b",
         10158 => x"807a3480",
         10159 => x"5380df3d",
         10160 => x"fdb40552",
         10161 => x"80e03d51",
         10162 => x"e8953f82",
         10163 => x"d8c80857",
         10164 => x"82d8c808",
         10165 => x"83a1387b",
         10166 => x"80d43d0c",
         10167 => x"7a7c9811",
         10168 => x"0880d83d",
         10169 => x"0c555880",
         10170 => x"d53d0854",
         10171 => x"73802e82",
         10172 => x"8338a052",
         10173 => x"80d33d70",
         10174 => x"5255c4d4",
         10175 => x"3f82d8c8",
         10176 => x"085782d8",
         10177 => x"c80882ef",
         10178 => x"3880d93d",
         10179 => x"08527b51",
         10180 => x"ffb8ae3f",
         10181 => x"82d8c808",
         10182 => x"5782d8c8",
         10183 => x"0882d838",
         10184 => x"80da3d08",
         10185 => x"527b51c9",
         10186 => x"863f82d8",
         10187 => x"c80880d6",
         10188 => x"3d0c7652",
         10189 => x"7451c498",
         10190 => x"3f82d8c8",
         10191 => x"085782d8",
         10192 => x"c80882b3",
         10193 => x"38805274",
         10194 => x"51c9fa3f",
         10195 => x"82d8c808",
         10196 => x"5782d8c8",
         10197 => x"08a73880",
         10198 => x"da3d0852",
         10199 => x"7b51c8cf",
         10200 => x"3f7382d8",
         10201 => x"c8082ea6",
         10202 => x"38765274",
         10203 => x"51c5ac3f",
         10204 => x"82d8c808",
         10205 => x"5782d8c8",
         10206 => x"08802ec9",
         10207 => x"3876842e",
         10208 => x"09810686",
         10209 => x"38825781",
         10210 => x"ee397681",
         10211 => x"ea3880df",
         10212 => x"3dfdb805",
         10213 => x"527451d6",
         10214 => x"e43f7693",
         10215 => x"3d781182",
         10216 => x"11335156",
         10217 => x"5a567380",
         10218 => x"2e923802",
         10219 => x"80c60555",
         10220 => x"81168116",
         10221 => x"70335656",
         10222 => x"5673f538",
         10223 => x"81165473",
         10224 => x"78268199",
         10225 => x"3875802e",
         10226 => x"9c387816",
         10227 => x"820555ff",
         10228 => x"1880e13d",
         10229 => x"0811ff18",
         10230 => x"ff185858",
         10231 => x"55587433",
         10232 => x"743475eb",
         10233 => x"38ff1880",
         10234 => x"e13d0811",
         10235 => x"5558af74",
         10236 => x"34fdf439",
         10237 => x"777b2e09",
         10238 => x"81068d38",
         10239 => x"ff1880e1",
         10240 => x"3d081155",
         10241 => x"58af7434",
         10242 => x"800b82f0",
         10243 => x"a4337084",
         10244 => x"2982cac0",
         10245 => x"05700870",
         10246 => x"33525c56",
         10247 => x"56567376",
         10248 => x"2e8d3881",
         10249 => x"16701a70",
         10250 => x"33515556",
         10251 => x"73f53882",
         10252 => x"16547378",
         10253 => x"26a73880",
         10254 => x"55747627",
         10255 => x"91387419",
         10256 => x"5473337a",
         10257 => x"7081055c",
         10258 => x"34811555",
         10259 => x"ec39ba7a",
         10260 => x"7081055c",
         10261 => x"3474ff2e",
         10262 => x"09810685",
         10263 => x"38915797",
         10264 => x"3980e03d",
         10265 => x"08188119",
         10266 => x"59547333",
         10267 => x"7a708105",
         10268 => x"5c347a78",
         10269 => x"26eb3880",
         10270 => x"7a347682",
         10271 => x"d8c80c80",
         10272 => x"df3d0d04",
         10273 => x"f73d0d7b",
         10274 => x"7d8d3dfc",
         10275 => x"05547153",
         10276 => x"5755ebfd",
         10277 => x"3f82d8c8",
         10278 => x"085382d8",
         10279 => x"c80882fe",
         10280 => x"38911533",
         10281 => x"537282f6",
         10282 => x"388c1508",
         10283 => x"54737627",
         10284 => x"92389015",
         10285 => x"3370812a",
         10286 => x"70810651",
         10287 => x"54577283",
         10288 => x"38735694",
         10289 => x"15085480",
         10290 => x"7094170c",
         10291 => x"5875782e",
         10292 => x"829b3879",
         10293 => x"8a112270",
         10294 => x"892b5951",
         10295 => x"5373782e",
         10296 => x"b7387652",
         10297 => x"ff1651fe",
         10298 => x"c5993f82",
         10299 => x"d8c808ff",
         10300 => x"15785470",
         10301 => x"535553fe",
         10302 => x"c5893f82",
         10303 => x"d8c80873",
         10304 => x"26963876",
         10305 => x"30707506",
         10306 => x"7094180c",
         10307 => x"77713198",
         10308 => x"18085758",
         10309 => x"5153b239",
         10310 => x"88150854",
         10311 => x"73a73873",
         10312 => x"527451ff",
         10313 => x"bc973f82",
         10314 => x"d8c80854",
         10315 => x"82d8c808",
         10316 => x"812e819d",
         10317 => x"3882d8c8",
         10318 => x"08ff2e81",
         10319 => x"9e3882d8",
         10320 => x"c8088816",
         10321 => x"0c739816",
         10322 => x"0c73802e",
         10323 => x"819f3876",
         10324 => x"762780de",
         10325 => x"38757731",
         10326 => x"94160818",
         10327 => x"94170c90",
         10328 => x"16337081",
         10329 => x"2a708106",
         10330 => x"51555a56",
         10331 => x"72802e9b",
         10332 => x"38735274",
         10333 => x"51ffbbc5",
         10334 => x"3f82d8c8",
         10335 => x"085482d8",
         10336 => x"c8089538",
         10337 => x"82d8c808",
         10338 => x"56a83973",
         10339 => x"527451ff",
         10340 => x"b5cf3f82",
         10341 => x"d8c80854",
         10342 => x"73ff2ebf",
         10343 => x"38817427",
         10344 => x"b0387953",
         10345 => x"739c1408",
         10346 => x"27a73873",
         10347 => x"98160cff",
         10348 => x"9e399415",
         10349 => x"08169416",
         10350 => x"0c7583ff",
         10351 => x"06537280",
         10352 => x"2eab3873",
         10353 => x"527951ff",
         10354 => x"b4ed3f82",
         10355 => x"d8c80894",
         10356 => x"38820b91",
         10357 => x"16348253",
         10358 => x"80c43981",
         10359 => x"0b911634",
         10360 => x"8153bb39",
         10361 => x"75892a82",
         10362 => x"d8c80805",
         10363 => x"58941508",
         10364 => x"548c1508",
         10365 => x"74279038",
         10366 => x"738c160c",
         10367 => x"90153380",
         10368 => x"c0075372",
         10369 => x"90163473",
         10370 => x"83ff0653",
         10371 => x"72802e8c",
         10372 => x"38779c16",
         10373 => x"082e8538",
         10374 => x"779c160c",
         10375 => x"80537282",
         10376 => x"d8c80c8b",
         10377 => x"3d0d04f9",
         10378 => x"3d0d7956",
         10379 => x"89547580",
         10380 => x"2e818b38",
         10381 => x"8053893d",
         10382 => x"fc05528a",
         10383 => x"3d840551",
         10384 => x"e19d3f82",
         10385 => x"d8c80855",
         10386 => x"82d8c808",
         10387 => x"80eb3877",
         10388 => x"760c7a52",
         10389 => x"7551d5a1",
         10390 => x"3f82d8c8",
         10391 => x"085582d8",
         10392 => x"c80880c4",
         10393 => x"38ab1633",
         10394 => x"70982b55",
         10395 => x"57807424",
         10396 => x"a2388616",
         10397 => x"3370842a",
         10398 => x"70810651",
         10399 => x"55577380",
         10400 => x"2eae389c",
         10401 => x"16085277",
         10402 => x"51c2a43f",
         10403 => x"82d8c808",
         10404 => x"88170c77",
         10405 => x"54861422",
         10406 => x"84172374",
         10407 => x"527551ff",
         10408 => x"bdae3f82",
         10409 => x"d8c80855",
         10410 => x"74842e09",
         10411 => x"81068538",
         10412 => x"85558639",
         10413 => x"74802e84",
         10414 => x"3880760c",
         10415 => x"74547382",
         10416 => x"d8c80c89",
         10417 => x"3d0d04fc",
         10418 => x"3d0d7687",
         10419 => x"3dfc0553",
         10420 => x"705253e7",
         10421 => x"bc3f82d8",
         10422 => x"c8088738",
         10423 => x"82d8c808",
         10424 => x"730c863d",
         10425 => x"0d04fb3d",
         10426 => x"0d777989",
         10427 => x"3dfc0554",
         10428 => x"71535654",
         10429 => x"e79b3f82",
         10430 => x"d8c80853",
         10431 => x"82d8c808",
         10432 => x"80e13874",
         10433 => x"943882d8",
         10434 => x"c8085273",
         10435 => x"51ffbcc0",
         10436 => x"3f82d8c8",
         10437 => x"085380cb",
         10438 => x"3982d8c8",
         10439 => x"08527351",
         10440 => x"c2a33f82",
         10441 => x"d8c80853",
         10442 => x"82d8c808",
         10443 => x"842e0981",
         10444 => x"06853880",
         10445 => x"53873982",
         10446 => x"d8c808a7",
         10447 => x"38745273",
         10448 => x"51cfba3f",
         10449 => x"72527351",
         10450 => x"ffbdd03f",
         10451 => x"82d8c808",
         10452 => x"84327030",
         10453 => x"7072079f",
         10454 => x"2c7082d8",
         10455 => x"c8080651",
         10456 => x"51545472",
         10457 => x"82d8c80c",
         10458 => x"873d0d04",
         10459 => x"ed3d0d66",
         10460 => x"57805389",
         10461 => x"3d705397",
         10462 => x"3d5256de",
         10463 => x"e23f82d8",
         10464 => x"c8085582",
         10465 => x"d8c808b2",
         10466 => x"38655275",
         10467 => x"51d2ea3f",
         10468 => x"82d8c808",
         10469 => x"5582d8c8",
         10470 => x"08a03802",
         10471 => x"80cb0533",
         10472 => x"70982b55",
         10473 => x"58738025",
         10474 => x"85388655",
         10475 => x"8d397680",
         10476 => x"2e883876",
         10477 => x"527551ce",
         10478 => x"c43f7482",
         10479 => x"d8c80c95",
         10480 => x"3d0d04f0",
         10481 => x"3d0d6365",
         10482 => x"555c8053",
         10483 => x"923dec05",
         10484 => x"52933d51",
         10485 => x"de893f82",
         10486 => x"d8c8085b",
         10487 => x"82d8c808",
         10488 => x"8282387c",
         10489 => x"740c7308",
         10490 => x"9c1108fe",
         10491 => x"11941308",
         10492 => x"59565855",
         10493 => x"75742691",
         10494 => x"38757c0c",
         10495 => x"81e63981",
         10496 => x"5b81ce39",
         10497 => x"825b81c9",
         10498 => x"3982d8c8",
         10499 => x"08753355",
         10500 => x"5973812e",
         10501 => x"09810680",
         10502 => x"c0388275",
         10503 => x"5f577652",
         10504 => x"923df005",
         10505 => x"51ffb0b9",
         10506 => x"3f82d8c8",
         10507 => x"08ff2ecf",
         10508 => x"3882d8c8",
         10509 => x"08812ecc",
         10510 => x"3882d8c8",
         10511 => x"08307082",
         10512 => x"d8c80807",
         10513 => x"80257a05",
         10514 => x"81197f53",
         10515 => x"595a549c",
         10516 => x"14087726",
         10517 => x"c93880f9",
         10518 => x"39a81508",
         10519 => x"82d8c808",
         10520 => x"57587598",
         10521 => x"38775281",
         10522 => x"187d5258",
         10523 => x"ffadd23f",
         10524 => x"82d8c808",
         10525 => x"5b82d8c8",
         10526 => x"0880d638",
         10527 => x"7c703377",
         10528 => x"12ff1a5d",
         10529 => x"52565474",
         10530 => x"822e0981",
         10531 => x"069e38b8",
         10532 => x"1451ffa9",
         10533 => x"d23f82d8",
         10534 => x"c80883ff",
         10535 => x"ff067030",
         10536 => x"7080251b",
         10537 => x"8219595b",
         10538 => x"51549b39",
         10539 => x"b81451ff",
         10540 => x"a9cc3f82",
         10541 => x"d8c808f0",
         10542 => x"0a067030",
         10543 => x"7080251b",
         10544 => x"8419595b",
         10545 => x"51547583",
         10546 => x"ff067a58",
         10547 => x"5679ff92",
         10548 => x"38787c0c",
         10549 => x"7c799412",
         10550 => x"0c841133",
         10551 => x"81075654",
         10552 => x"74841534",
         10553 => x"7a82d8c8",
         10554 => x"0c923d0d",
         10555 => x"04f93d0d",
         10556 => x"798a3dfc",
         10557 => x"05537052",
         10558 => x"57e3963f",
         10559 => x"82d8c808",
         10560 => x"5682d8c8",
         10561 => x"0881aa38",
         10562 => x"91173356",
         10563 => x"7581a238",
         10564 => x"90173370",
         10565 => x"812a7081",
         10566 => x"06515555",
         10567 => x"87557380",
         10568 => x"2e819038",
         10569 => x"94170854",
         10570 => x"738c1808",
         10571 => x"27818238",
         10572 => x"739c3882",
         10573 => x"d8c80853",
         10574 => x"88170852",
         10575 => x"7651ffb2",
         10576 => x"d03f82d8",
         10577 => x"c8087488",
         10578 => x"190c5680",
         10579 => x"ca399817",
         10580 => x"08527651",
         10581 => x"ffae8a3f",
         10582 => x"82d8c808",
         10583 => x"ff2e0981",
         10584 => x"06833881",
         10585 => x"5682d8c8",
         10586 => x"08812e09",
         10587 => x"81068538",
         10588 => x"8256a439",
         10589 => x"75a13877",
         10590 => x"5482d8c8",
         10591 => x"089c1508",
         10592 => x"27953898",
         10593 => x"17085382",
         10594 => x"d8c80852",
         10595 => x"7651ffb2",
         10596 => x"803f82d8",
         10597 => x"c8085694",
         10598 => x"17088c18",
         10599 => x"0c901733",
         10600 => x"80c00754",
         10601 => x"73901834",
         10602 => x"75802e85",
         10603 => x"38759118",
         10604 => x"34755574",
         10605 => x"82d8c80c",
         10606 => x"893d0d04",
         10607 => x"e03d0d82",
         10608 => x"53a23dff",
         10609 => x"9c0552a3",
         10610 => x"3d51da93",
         10611 => x"3f82d8c8",
         10612 => x"085582d8",
         10613 => x"c80881f9",
         10614 => x"387846a3",
         10615 => x"3d085296",
         10616 => x"3d705258",
         10617 => x"ce933f82",
         10618 => x"d8c80855",
         10619 => x"82d8c808",
         10620 => x"81df3802",
         10621 => x"80ff0533",
         10622 => x"70852a70",
         10623 => x"81065155",
         10624 => x"56865573",
         10625 => x"81cb3875",
         10626 => x"982b5480",
         10627 => x"742481c1",
         10628 => x"380280da",
         10629 => x"05337081",
         10630 => x"06585487",
         10631 => x"557681b1",
         10632 => x"386c5278",
         10633 => x"51ffbb87",
         10634 => x"3f82d8c8",
         10635 => x"0874842a",
         10636 => x"70810651",
         10637 => x"55567380",
         10638 => x"2e80d638",
         10639 => x"785482d8",
         10640 => x"c8089815",
         10641 => x"082e8189",
         10642 => x"38735a82",
         10643 => x"d8c8085c",
         10644 => x"76528a3d",
         10645 => x"705254ff",
         10646 => x"b5f63f82",
         10647 => x"d8c80855",
         10648 => x"82d8c808",
         10649 => x"80eb3882",
         10650 => x"d8c80852",
         10651 => x"7351ffbb",
         10652 => x"d43f82d8",
         10653 => x"c8085582",
         10654 => x"d8c80886",
         10655 => x"38875580",
         10656 => x"d03982d8",
         10657 => x"c808842e",
         10658 => x"883882d8",
         10659 => x"c80880c1",
         10660 => x"387751c7",
         10661 => x"ef3f82d8",
         10662 => x"c80882d8",
         10663 => x"c8083070",
         10664 => x"82d8c808",
         10665 => x"07802551",
         10666 => x"55557580",
         10667 => x"2e953873",
         10668 => x"802e9038",
         10669 => x"80537552",
         10670 => x"7751ffaf",
         10671 => x"d43f82d8",
         10672 => x"c8085574",
         10673 => x"8c387851",
         10674 => x"ffa9bd3f",
         10675 => x"82d8c808",
         10676 => x"557482d8",
         10677 => x"c80ca23d",
         10678 => x"0d04e83d",
         10679 => x"0d82539a",
         10680 => x"3dffbc05",
         10681 => x"529b3d51",
         10682 => x"d7f53f82",
         10683 => x"d8c80854",
         10684 => x"82d8c808",
         10685 => x"82b73878",
         10686 => x"5e6a528e",
         10687 => x"3d705258",
         10688 => x"cbf73f82",
         10689 => x"d8c80854",
         10690 => x"82d8c808",
         10691 => x"86388854",
         10692 => x"829b3982",
         10693 => x"d8c80884",
         10694 => x"2e098106",
         10695 => x"828f3802",
         10696 => x"80df0533",
         10697 => x"70852a81",
         10698 => x"06515586",
         10699 => x"547481fd",
         10700 => x"38785a74",
         10701 => x"528a3d70",
         10702 => x"5257ffb0",
         10703 => x"803f82d8",
         10704 => x"c8087555",
         10705 => x"5682d8c8",
         10706 => x"08833887",
         10707 => x"5482d8c8",
         10708 => x"08812e09",
         10709 => x"81068338",
         10710 => x"825482d8",
         10711 => x"c808ff2e",
         10712 => x"09810686",
         10713 => x"38815481",
         10714 => x"ba397381",
         10715 => x"b63882d8",
         10716 => x"c8085278",
         10717 => x"51ffb2e0",
         10718 => x"3f82d8c8",
         10719 => x"085482d8",
         10720 => x"c808819f",
         10721 => x"388b53a0",
         10722 => x"52b81951",
         10723 => x"ffa58a3f",
         10724 => x"7854ae0b",
         10725 => x"b8153478",
         10726 => x"54900b80",
         10727 => x"c3153482",
         10728 => x"88b20a52",
         10729 => x"80ce1951",
         10730 => x"ffa49c3f",
         10731 => x"755378b8",
         10732 => x"115351ff",
         10733 => x"b8b23fa0",
         10734 => x"5378b811",
         10735 => x"5380d805",
         10736 => x"51ffa4b2",
         10737 => x"3f7854ae",
         10738 => x"0b80d915",
         10739 => x"347f5378",
         10740 => x"80d81153",
         10741 => x"51ffb890",
         10742 => x"3f785481",
         10743 => x"0b831534",
         10744 => x"7751ffbf",
         10745 => x"cd3f82d8",
         10746 => x"c8085482",
         10747 => x"d8c808b3",
         10748 => x"388288b2",
         10749 => x"0a526496",
         10750 => x"0551ffa3",
         10751 => x"ca3f7553",
         10752 => x"64527851",
         10753 => x"ffb7e13f",
         10754 => x"6454900b",
         10755 => x"8b153478",
         10756 => x"54810b83",
         10757 => x"15347851",
         10758 => x"ffa6ed3f",
         10759 => x"82d8c808",
         10760 => x"548b3980",
         10761 => x"53755276",
         10762 => x"51fface5",
         10763 => x"3f7382d8",
         10764 => x"c80c9a3d",
         10765 => x"0d04d83d",
         10766 => x"0dab3d84",
         10767 => x"0551d294",
         10768 => x"3f8253aa",
         10769 => x"3dfefc05",
         10770 => x"52ab3d51",
         10771 => x"d5913f82",
         10772 => x"d8c80855",
         10773 => x"82d8c808",
         10774 => x"82d83878",
         10775 => x"4eab3d08",
         10776 => x"529e3d70",
         10777 => x"5258c991",
         10778 => x"3f82d8c8",
         10779 => x"085582d8",
         10780 => x"c80882be",
         10781 => x"3802819f",
         10782 => x"053381a0",
         10783 => x"06548655",
         10784 => x"7382af38",
         10785 => x"a053a53d",
         10786 => x"0852aa3d",
         10787 => x"ff800551",
         10788 => x"ffa2e33f",
         10789 => x"b0537752",
         10790 => x"923d7052",
         10791 => x"54ffa2d6",
         10792 => x"3fac3d08",
         10793 => x"527351c8",
         10794 => x"d03f82d8",
         10795 => x"c8085582",
         10796 => x"d8c80897",
         10797 => x"3863a13d",
         10798 => x"082e0981",
         10799 => x"06883865",
         10800 => x"a33d082e",
         10801 => x"92388855",
         10802 => x"81e83982",
         10803 => x"d8c80884",
         10804 => x"2e098106",
         10805 => x"81bb3873",
         10806 => x"51ffbdd6",
         10807 => x"3f82d8c8",
         10808 => x"085582d8",
         10809 => x"c80881ca",
         10810 => x"38685693",
         10811 => x"53aa3dff",
         10812 => x"8d05528d",
         10813 => x"1651ffa1",
         10814 => x"fd3f02af",
         10815 => x"05338b17",
         10816 => x"348b1633",
         10817 => x"70842a70",
         10818 => x"81065155",
         10819 => x"55738938",
         10820 => x"74a00754",
         10821 => x"738b1734",
         10822 => x"7854810b",
         10823 => x"8315348b",
         10824 => x"16337084",
         10825 => x"2a708106",
         10826 => x"51555573",
         10827 => x"802e80e7",
         10828 => x"386f642e",
         10829 => x"80e13875",
         10830 => x"527851ff",
         10831 => x"b4f13f82",
         10832 => x"d8c80852",
         10833 => x"7851ffa5",
         10834 => x"ee3f8255",
         10835 => x"82d8c808",
         10836 => x"802e80de",
         10837 => x"3882d8c8",
         10838 => x"08527851",
         10839 => x"ffa3e23f",
         10840 => x"82d8c808",
         10841 => x"7980d811",
         10842 => x"58585582",
         10843 => x"d8c80880",
         10844 => x"c1388116",
         10845 => x"335473ae",
         10846 => x"2e098106",
         10847 => x"9a386353",
         10848 => x"75527651",
         10849 => x"ffb4e13f",
         10850 => x"7854810b",
         10851 => x"83153487",
         10852 => x"3982d8c8",
         10853 => x"089c3877",
         10854 => x"51c1e93f",
         10855 => x"82d8c808",
         10856 => x"5582d8c8",
         10857 => x"088c3878",
         10858 => x"51ffa3dc",
         10859 => x"3f82d8c8",
         10860 => x"08557482",
         10861 => x"d8c80caa",
         10862 => x"3d0d04ec",
         10863 => x"3d0d0280",
         10864 => x"df053302",
         10865 => x"840580e3",
         10866 => x"05335757",
         10867 => x"8253963d",
         10868 => x"cc055297",
         10869 => x"3d51d287",
         10870 => x"3f82d8c8",
         10871 => x"085582d8",
         10872 => x"c80880cf",
         10873 => x"38785a66",
         10874 => x"52963dd0",
         10875 => x"0551c689",
         10876 => x"3f82d8c8",
         10877 => x"085582d8",
         10878 => x"c808b838",
         10879 => x"0280cf05",
         10880 => x"3381a006",
         10881 => x"54865573",
         10882 => x"aa3875a7",
         10883 => x"06617109",
         10884 => x"8b123371",
         10885 => x"067a7406",
         10886 => x"07515755",
         10887 => x"56748b15",
         10888 => x"34785481",
         10889 => x"0b831534",
         10890 => x"7851ffa2",
         10891 => x"db3f82d8",
         10892 => x"c8085574",
         10893 => x"82d8c80c",
         10894 => x"963d0d04",
         10895 => x"ee3d0d65",
         10896 => x"56825394",
         10897 => x"3dcc0552",
         10898 => x"953d51d1",
         10899 => x"923f82d8",
         10900 => x"c8085582",
         10901 => x"d8c80880",
         10902 => x"cb387658",
         10903 => x"6452943d",
         10904 => x"d00551c5",
         10905 => x"943f82d8",
         10906 => x"c8085582",
         10907 => x"d8c808b4",
         10908 => x"380280c7",
         10909 => x"053381a0",
         10910 => x"06548655",
         10911 => x"73a63884",
         10912 => x"16228617",
         10913 => x"2271902b",
         10914 => x"07535496",
         10915 => x"1f51ff9e",
         10916 => x"b63f7654",
         10917 => x"810b8315",
         10918 => x"347651ff",
         10919 => x"a1ea3f82",
         10920 => x"d8c80855",
         10921 => x"7482d8c8",
         10922 => x"0c943d0d",
         10923 => x"04e93d0d",
         10924 => x"6a6c5c5a",
         10925 => x"8053993d",
         10926 => x"cc05529a",
         10927 => x"3d51d09f",
         10928 => x"3f82d8c8",
         10929 => x"0882d8c8",
         10930 => x"08307082",
         10931 => x"d8c80807",
         10932 => x"80255155",
         10933 => x"5779802e",
         10934 => x"81863881",
         10935 => x"70750655",
         10936 => x"5573802e",
         10937 => x"80fa387b",
         10938 => x"5d805f80",
         10939 => x"528d3d70",
         10940 => x"5254ffac",
         10941 => x"db3f82d8",
         10942 => x"c8085782",
         10943 => x"d8c80880",
         10944 => x"d2387452",
         10945 => x"7351ffb2",
         10946 => x"bc3f82d8",
         10947 => x"c8085782",
         10948 => x"d8c808bf",
         10949 => x"3882d8c8",
         10950 => x"0882d8c8",
         10951 => x"08655b59",
         10952 => x"56781881",
         10953 => x"197b1856",
         10954 => x"59557433",
         10955 => x"74348116",
         10956 => x"568a7827",
         10957 => x"ec388b56",
         10958 => x"751a5480",
         10959 => x"74347580",
         10960 => x"2e9e38ff",
         10961 => x"16701b70",
         10962 => x"33515556",
         10963 => x"73a02ee8",
         10964 => x"388e3976",
         10965 => x"842e0981",
         10966 => x"06863880",
         10967 => x"7a348057",
         10968 => x"76307078",
         10969 => x"07802551",
         10970 => x"547a802e",
         10971 => x"80c13873",
         10972 => x"802ebc38",
         10973 => x"7ba41108",
         10974 => x"5351ff9f",
         10975 => x"c43f82d8",
         10976 => x"c8085782",
         10977 => x"d8c808a7",
         10978 => x"387b7033",
         10979 => x"555580c3",
         10980 => x"5673832e",
         10981 => x"8b3880e4",
         10982 => x"5673842e",
         10983 => x"8338a756",
         10984 => x"7515b805",
         10985 => x"51ff9bd6",
         10986 => x"3f82d8c8",
         10987 => x"087b0c76",
         10988 => x"82d8c80c",
         10989 => x"993d0d04",
         10990 => x"e63d0d82",
         10991 => x"539c3dff",
         10992 => x"b405529d",
         10993 => x"3d51ce97",
         10994 => x"3f82d8c8",
         10995 => x"0882d8c8",
         10996 => x"08565482",
         10997 => x"d8c80882",
         10998 => x"dd388b53",
         10999 => x"a0528a3d",
         11000 => x"705258ff",
         11001 => x"9cb33f73",
         11002 => x"6d703351",
         11003 => x"55569f74",
         11004 => x"27818638",
         11005 => x"77579d3d",
         11006 => x"51ff9d90",
         11007 => x"3f82d8c8",
         11008 => x"0883ffff",
         11009 => x"2680c438",
         11010 => x"82d8c808",
         11011 => x"5195983f",
         11012 => x"83b55282",
         11013 => x"d8c80851",
         11014 => x"93e83f82",
         11015 => x"d8c80883",
         11016 => x"ffff0655",
         11017 => x"74802ea3",
         11018 => x"38745282",
         11019 => x"cbe051ff",
         11020 => x"9cb23f82",
         11021 => x"d8c80893",
         11022 => x"3881ff75",
         11023 => x"27883875",
         11024 => x"89268838",
         11025 => x"8b398a76",
         11026 => x"27863886",
         11027 => x"5581e739",
         11028 => x"81ff7527",
         11029 => x"8f387488",
         11030 => x"2a547377",
         11031 => x"70810559",
         11032 => x"34811656",
         11033 => x"74777081",
         11034 => x"05593481",
         11035 => x"166d7033",
         11036 => x"51555673",
         11037 => x"9f26fefe",
         11038 => x"388a3d33",
         11039 => x"54865573",
         11040 => x"81e52e81",
         11041 => x"b1387580",
         11042 => x"2e993802",
         11043 => x"a3055575",
         11044 => x"15703351",
         11045 => x"5473a02e",
         11046 => x"09810687",
         11047 => x"38ff1656",
         11048 => x"75ed3878",
         11049 => x"40804280",
         11050 => x"52903d70",
         11051 => x"5255ffa9",
         11052 => x"9f3f82d8",
         11053 => x"c8085482",
         11054 => x"d8c80880",
         11055 => x"f7388152",
         11056 => x"7451ffaf",
         11057 => x"803f82d8",
         11058 => x"c8085482",
         11059 => x"d8c8088d",
         11060 => x"387580c4",
         11061 => x"386654e5",
         11062 => x"743480c6",
         11063 => x"3982d8c8",
         11064 => x"08842e09",
         11065 => x"810680cc",
         11066 => x"38805475",
         11067 => x"742e80c4",
         11068 => x"38815274",
         11069 => x"51ffac9c",
         11070 => x"3f82d8c8",
         11071 => x"085482d8",
         11072 => x"c808b138",
         11073 => x"a05382d8",
         11074 => x"c8085266",
         11075 => x"51ff9a89",
         11076 => x"3f665488",
         11077 => x"0b8b1534",
         11078 => x"8b537752",
         11079 => x"6651ff99",
         11080 => x"d53f7854",
         11081 => x"810b8315",
         11082 => x"347851ff",
         11083 => x"9cda3f82",
         11084 => x"d8c80854",
         11085 => x"73557482",
         11086 => x"d8c80c9c",
         11087 => x"3d0d04f2",
         11088 => x"3d0d6062",
         11089 => x"02880580",
         11090 => x"cb053393",
         11091 => x"3dfc0555",
         11092 => x"7254405e",
         11093 => x"5ad2ba3f",
         11094 => x"82d8c808",
         11095 => x"5882d8c8",
         11096 => x"0882bd38",
         11097 => x"911a3358",
         11098 => x"7782b538",
         11099 => x"7c802e97",
         11100 => x"388c1a08",
         11101 => x"59789038",
         11102 => x"901a3370",
         11103 => x"812a7081",
         11104 => x"06515555",
         11105 => x"73903887",
         11106 => x"54829739",
         11107 => x"82588290",
         11108 => x"39815882",
         11109 => x"8b397e8a",
         11110 => x"11227089",
         11111 => x"2b70557f",
         11112 => x"54565656",
         11113 => x"feabdc3f",
         11114 => x"ff147d06",
         11115 => x"70307072",
         11116 => x"079f2a82",
         11117 => x"d8c80805",
         11118 => x"9019087c",
         11119 => x"405a5d55",
         11120 => x"55817727",
         11121 => x"88389c16",
         11122 => x"08772683",
         11123 => x"38825776",
         11124 => x"77565980",
         11125 => x"56745279",
         11126 => x"51ff9d85",
         11127 => x"3f81157f",
         11128 => x"55559c14",
         11129 => x"08752683",
         11130 => x"38825582",
         11131 => x"d8c80881",
         11132 => x"2eff9938",
         11133 => x"82d8c808",
         11134 => x"ff2eff95",
         11135 => x"3882d8c8",
         11136 => x"088e3881",
         11137 => x"1656757b",
         11138 => x"2e098106",
         11139 => x"87389339",
         11140 => x"74598056",
         11141 => x"74772e09",
         11142 => x"8106ffb9",
         11143 => x"38875880",
         11144 => x"ff397d80",
         11145 => x"2eba3878",
         11146 => x"7b55557a",
         11147 => x"802eb438",
         11148 => x"81155673",
         11149 => x"812e0981",
         11150 => x"068338ff",
         11151 => x"56755374",
         11152 => x"527e51ff",
         11153 => x"9e943f82",
         11154 => x"d8c80858",
         11155 => x"82d8c808",
         11156 => x"80ce3874",
         11157 => x"8116ff16",
         11158 => x"56565c73",
         11159 => x"d3388439",
         11160 => x"ff195c7e",
         11161 => x"7c90120c",
         11162 => x"557d802e",
         11163 => x"b3387888",
         11164 => x"1b0c7c8c",
         11165 => x"1b0c901a",
         11166 => x"3380c007",
         11167 => x"5473901b",
         11168 => x"349c1508",
         11169 => x"fe059416",
         11170 => x"08575475",
         11171 => x"74269138",
         11172 => x"757b3194",
         11173 => x"160c8415",
         11174 => x"33810754",
         11175 => x"73841634",
         11176 => x"77547382",
         11177 => x"d8c80c90",
         11178 => x"3d0d04e9",
         11179 => x"3d0d6b6d",
         11180 => x"02880580",
         11181 => x"eb05339d",
         11182 => x"3d545a5c",
         11183 => x"59c5953f",
         11184 => x"8b56800b",
         11185 => x"82d8c808",
         11186 => x"248bf838",
         11187 => x"82d8c808",
         11188 => x"842982f0",
         11189 => x"90057008",
         11190 => x"51557480",
         11191 => x"2e843880",
         11192 => x"753482d8",
         11193 => x"c80881ff",
         11194 => x"065f8152",
         11195 => x"7e51ff8e",
         11196 => x"fe3f82d8",
         11197 => x"c80881ff",
         11198 => x"06708106",
         11199 => x"56578356",
         11200 => x"748bc038",
         11201 => x"76822a70",
         11202 => x"81065155",
         11203 => x"8a56748b",
         11204 => x"b238993d",
         11205 => x"fc055383",
         11206 => x"527e51ff",
         11207 => x"939e3f82",
         11208 => x"d8c80899",
         11209 => x"38675574",
         11210 => x"802e9238",
         11211 => x"74828080",
         11212 => x"268b38ff",
         11213 => x"15750655",
         11214 => x"74802e83",
         11215 => x"38814878",
         11216 => x"802e8738",
         11217 => x"84807926",
         11218 => x"92387881",
         11219 => x"800a268b",
         11220 => x"38ff1979",
         11221 => x"06557480",
         11222 => x"2e863893",
         11223 => x"568ae439",
         11224 => x"78892a6e",
         11225 => x"892a7089",
         11226 => x"2b775948",
         11227 => x"43597a83",
         11228 => x"38815661",
         11229 => x"30708025",
         11230 => x"77075155",
         11231 => x"9156748a",
         11232 => x"c238993d",
         11233 => x"f8055381",
         11234 => x"527e51ff",
         11235 => x"92ae3f81",
         11236 => x"5682d8c8",
         11237 => x"088aac38",
         11238 => x"77832a70",
         11239 => x"770682d8",
         11240 => x"c8084356",
         11241 => x"45748338",
         11242 => x"bf416655",
         11243 => x"8e566075",
         11244 => x"268a9038",
         11245 => x"74613170",
         11246 => x"485580ff",
         11247 => x"75278a83",
         11248 => x"38935678",
         11249 => x"81802689",
         11250 => x"fa387781",
         11251 => x"2a708106",
         11252 => x"56437480",
         11253 => x"2e953877",
         11254 => x"87065574",
         11255 => x"822e838d",
         11256 => x"38778106",
         11257 => x"5574802e",
         11258 => x"83833877",
         11259 => x"81065593",
         11260 => x"56825e74",
         11261 => x"802e89cb",
         11262 => x"38785a7d",
         11263 => x"832e0981",
         11264 => x"0680e138",
         11265 => x"78ae3866",
         11266 => x"912a5781",
         11267 => x"0b82cc84",
         11268 => x"22565a74",
         11269 => x"802e9d38",
         11270 => x"74772698",
         11271 => x"3882cc84",
         11272 => x"56791082",
         11273 => x"17702257",
         11274 => x"575a7480",
         11275 => x"2e863876",
         11276 => x"7527ee38",
         11277 => x"79526651",
         11278 => x"fea6c83f",
         11279 => x"82d8c808",
         11280 => x"84298487",
         11281 => x"0570892a",
         11282 => x"5e55a05c",
         11283 => x"800b82d8",
         11284 => x"c808fc80",
         11285 => x"8a055644",
         11286 => x"fdfff00a",
         11287 => x"752780ec",
         11288 => x"3888d339",
         11289 => x"78ae3866",
         11290 => x"8c2a5781",
         11291 => x"0b82cbf4",
         11292 => x"22565a74",
         11293 => x"802e9d38",
         11294 => x"74772698",
         11295 => x"3882cbf4",
         11296 => x"56791082",
         11297 => x"17702257",
         11298 => x"575a7480",
         11299 => x"2e863876",
         11300 => x"7527ee38",
         11301 => x"79526651",
         11302 => x"fea5e83f",
         11303 => x"82d8c808",
         11304 => x"10840557",
         11305 => x"82d8c808",
         11306 => x"9ff52696",
         11307 => x"38810b82",
         11308 => x"d8c80810",
         11309 => x"82d8c808",
         11310 => x"05711172",
         11311 => x"2a830559",
         11312 => x"565e83ff",
         11313 => x"17892a5d",
         11314 => x"815ca044",
         11315 => x"601c7d11",
         11316 => x"65056970",
         11317 => x"12ff0571",
         11318 => x"30707206",
         11319 => x"74315c52",
         11320 => x"59575940",
         11321 => x"7d832e09",
         11322 => x"81068938",
         11323 => x"761c6018",
         11324 => x"415c8439",
         11325 => x"761d5d79",
         11326 => x"90291870",
         11327 => x"62316858",
         11328 => x"51557476",
         11329 => x"2687af38",
         11330 => x"757c317d",
         11331 => x"317a5370",
         11332 => x"65315255",
         11333 => x"fea4ec3f",
         11334 => x"82d8c808",
         11335 => x"587d832e",
         11336 => x"0981069b",
         11337 => x"3882d8c8",
         11338 => x"0883fff5",
         11339 => x"2680dd38",
         11340 => x"78878338",
         11341 => x"79812a59",
         11342 => x"78fdbe38",
         11343 => x"86f8397d",
         11344 => x"822e0981",
         11345 => x"0680c538",
         11346 => x"83fff50b",
         11347 => x"82d8c808",
         11348 => x"27a03878",
         11349 => x"8f38791a",
         11350 => x"557480c0",
         11351 => x"26863874",
         11352 => x"59fd9639",
         11353 => x"62810655",
         11354 => x"74802e8f",
         11355 => x"38835efd",
         11356 => x"883982d8",
         11357 => x"c8089ff5",
         11358 => x"26923878",
         11359 => x"86b83879",
         11360 => x"1a598180",
         11361 => x"7927fcf1",
         11362 => x"3886ab39",
         11363 => x"80557d81",
         11364 => x"2e098106",
         11365 => x"83387d55",
         11366 => x"9ff57827",
         11367 => x"8b387481",
         11368 => x"06558e56",
         11369 => x"74869c38",
         11370 => x"84805380",
         11371 => x"527a51ff",
         11372 => x"90e73f8b",
         11373 => x"5382ca8c",
         11374 => x"527a51ff",
         11375 => x"90b83f84",
         11376 => x"80528b1b",
         11377 => x"51ff8fe1",
         11378 => x"3f798d1c",
         11379 => x"347b83ff",
         11380 => x"ff06528e",
         11381 => x"1b51ff8f",
         11382 => x"d03f810b",
         11383 => x"901c347d",
         11384 => x"83327030",
         11385 => x"70962a84",
         11386 => x"80065451",
         11387 => x"55911b51",
         11388 => x"ff8fb63f",
         11389 => x"66557483",
         11390 => x"ffff2690",
         11391 => x"387483ff",
         11392 => x"ff065293",
         11393 => x"1b51ff8f",
         11394 => x"a03f8a39",
         11395 => x"7452a01b",
         11396 => x"51ff8fb3",
         11397 => x"3ff80b95",
         11398 => x"1c34bf52",
         11399 => x"981b51ff",
         11400 => x"8f873f81",
         11401 => x"ff529a1b",
         11402 => x"51ff8efd",
         11403 => x"3f60529c",
         11404 => x"1b51ff8f",
         11405 => x"923f7d83",
         11406 => x"2e098106",
         11407 => x"80cb3882",
         11408 => x"88b20a52",
         11409 => x"80c31b51",
         11410 => x"ff8efc3f",
         11411 => x"7c52a41b",
         11412 => x"51ff8ef3",
         11413 => x"3f8252ac",
         11414 => x"1b51ff8e",
         11415 => x"ea3f8152",
         11416 => x"b01b51ff",
         11417 => x"8ec33f86",
         11418 => x"52b21b51",
         11419 => x"ff8eba3f",
         11420 => x"ff800b80",
         11421 => x"c01c34a9",
         11422 => x"0b80c21c",
         11423 => x"34935382",
         11424 => x"ca985280",
         11425 => x"c71b51ae",
         11426 => x"398288b2",
         11427 => x"0a52a71b",
         11428 => x"51ff8eb3",
         11429 => x"3f7c83ff",
         11430 => x"ff065296",
         11431 => x"1b51ff8e",
         11432 => x"883fff80",
         11433 => x"0ba41c34",
         11434 => x"a90ba61c",
         11435 => x"34935382",
         11436 => x"caac52ab",
         11437 => x"1b51ff8e",
         11438 => x"bd3f82d4",
         11439 => x"d55283fe",
         11440 => x"1b705259",
         11441 => x"ff8de23f",
         11442 => x"81546053",
         11443 => x"7a527e51",
         11444 => x"ff8a853f",
         11445 => x"815682d8",
         11446 => x"c80883e7",
         11447 => x"387d832e",
         11448 => x"09810680",
         11449 => x"ee387554",
         11450 => x"60860553",
         11451 => x"7a527e51",
         11452 => x"ff89e53f",
         11453 => x"84805380",
         11454 => x"527a51ff",
         11455 => x"8e9b3f84",
         11456 => x"8b85a4d2",
         11457 => x"527a51ff",
         11458 => x"8dbd3f86",
         11459 => x"8a85e4f2",
         11460 => x"5283e41b",
         11461 => x"51ff8daf",
         11462 => x"3fff1852",
         11463 => x"83e81b51",
         11464 => x"ff8da43f",
         11465 => x"825283ec",
         11466 => x"1b51ff8d",
         11467 => x"9a3f82d4",
         11468 => x"d5527851",
         11469 => x"ff8cf23f",
         11470 => x"75546087",
         11471 => x"05537a52",
         11472 => x"7e51ff89",
         11473 => x"933f7554",
         11474 => x"6016537a",
         11475 => x"527e51ff",
         11476 => x"89863f65",
         11477 => x"5380527a",
         11478 => x"51ff8dbd",
         11479 => x"3f7f5680",
         11480 => x"587d832e",
         11481 => x"0981069a",
         11482 => x"38f8527a",
         11483 => x"51ff8cd7",
         11484 => x"3fff5284",
         11485 => x"1b51ff8c",
         11486 => x"ce3ff00a",
         11487 => x"52881b51",
         11488 => x"913987ff",
         11489 => x"fff8557d",
         11490 => x"812e8338",
         11491 => x"f8557452",
         11492 => x"7a51ff8c",
         11493 => x"b23f7c55",
         11494 => x"61577462",
         11495 => x"26833874",
         11496 => x"57765475",
         11497 => x"537a527e",
         11498 => x"51ff88ac",
         11499 => x"3f82d8c8",
         11500 => x"08828738",
         11501 => x"84805382",
         11502 => x"d8c80852",
         11503 => x"7a51ff8c",
         11504 => x"d83f7616",
         11505 => x"75783156",
         11506 => x"5674cd38",
         11507 => x"81185877",
         11508 => x"802eff8d",
         11509 => x"3879557d",
         11510 => x"832e8338",
         11511 => x"63556157",
         11512 => x"74622683",
         11513 => x"38745776",
         11514 => x"5475537a",
         11515 => x"527e51ff",
         11516 => x"87e63f82",
         11517 => x"d8c80881",
         11518 => x"c1387616",
         11519 => x"75783156",
         11520 => x"5674db38",
         11521 => x"8c567d83",
         11522 => x"2e933886",
         11523 => x"566683ff",
         11524 => x"ff268a38",
         11525 => x"84567d82",
         11526 => x"2e833881",
         11527 => x"56648106",
         11528 => x"587780fe",
         11529 => x"38848053",
         11530 => x"77527a51",
         11531 => x"ff8bea3f",
         11532 => x"82d4d552",
         11533 => x"7851ff8a",
         11534 => x"f03f83be",
         11535 => x"1b557775",
         11536 => x"34810b81",
         11537 => x"1634810b",
         11538 => x"82163477",
         11539 => x"83163475",
         11540 => x"84163460",
         11541 => x"67055680",
         11542 => x"fdc15275",
         11543 => x"51fe9ea3",
         11544 => x"3ffe0b85",
         11545 => x"163482d8",
         11546 => x"c808822a",
         11547 => x"bf075675",
         11548 => x"86163482",
         11549 => x"d8c80887",
         11550 => x"16346052",
         11551 => x"83c61b51",
         11552 => x"ff8ac43f",
         11553 => x"665283ca",
         11554 => x"1b51ff8a",
         11555 => x"ba3f8154",
         11556 => x"77537a52",
         11557 => x"7e51ff86",
         11558 => x"bf3f8156",
         11559 => x"82d8c808",
         11560 => x"a2388053",
         11561 => x"80527e51",
         11562 => x"ff88913f",
         11563 => x"815682d8",
         11564 => x"c8089038",
         11565 => x"89398e56",
         11566 => x"8a398156",
         11567 => x"863982d8",
         11568 => x"c8085675",
         11569 => x"82d8c80c",
         11570 => x"993d0d04",
         11571 => x"f53d0d7d",
         11572 => x"605b5980",
         11573 => x"7960ff05",
         11574 => x"5a575776",
         11575 => x"7825b438",
         11576 => x"8d3df811",
         11577 => x"55558153",
         11578 => x"fc155279",
         11579 => x"51c9bd3f",
         11580 => x"7a812e09",
         11581 => x"81069c38",
         11582 => x"8c3d3355",
         11583 => x"748d2edb",
         11584 => x"38747670",
         11585 => x"81055834",
         11586 => x"81175774",
         11587 => x"8a2e0981",
         11588 => x"06c93880",
         11589 => x"76347855",
         11590 => x"76833876",
         11591 => x"557482d8",
         11592 => x"c80c8d3d",
         11593 => x"0d04f73d",
         11594 => x"0d7b0284",
         11595 => x"05b30533",
         11596 => x"5957778a",
         11597 => x"2e098106",
         11598 => x"87388d52",
         11599 => x"7651e73f",
         11600 => x"84170856",
         11601 => x"807624be",
         11602 => x"38881708",
         11603 => x"77178c05",
         11604 => x"56597775",
         11605 => x"34811656",
         11606 => x"bb7625a1",
         11607 => x"388b3dfc",
         11608 => x"05547553",
         11609 => x"8c175276",
         11610 => x"0851cbc0",
         11611 => x"3f797632",
         11612 => x"70307072",
         11613 => x"079f2a70",
         11614 => x"30535156",
         11615 => x"56758418",
         11616 => x"0c811988",
         11617 => x"180c8b3d",
         11618 => x"0d04f93d",
         11619 => x"0d798411",
         11620 => x"08565680",
         11621 => x"7524a738",
         11622 => x"893dfc05",
         11623 => x"5474538c",
         11624 => x"16527508",
         11625 => x"51cb853f",
         11626 => x"82d8c808",
         11627 => x"91388416",
         11628 => x"08782e09",
         11629 => x"81068738",
         11630 => x"88160855",
         11631 => x"8339ff55",
         11632 => x"7482d8c8",
         11633 => x"0c893d0d",
         11634 => x"04fd3d0d",
         11635 => x"755480cc",
         11636 => x"53805273",
         11637 => x"51ff88c1",
         11638 => x"3f76740c",
         11639 => x"853d0d04",
         11640 => x"ea3d0d02",
         11641 => x"80e30533",
         11642 => x"6a53863d",
         11643 => x"70535454",
         11644 => x"d83f7352",
         11645 => x"7251feae",
         11646 => x"3f7251ff",
         11647 => x"8d3f983d",
         11648 => x"0d04fd3d",
         11649 => x"0d750284",
         11650 => x"059a0522",
         11651 => x"55538052",
         11652 => x"7280ff26",
         11653 => x"8a387283",
         11654 => x"ffff0652",
         11655 => x"80c33983",
         11656 => x"ffff7327",
         11657 => x"517383b5",
         11658 => x"2e098106",
         11659 => x"b4387080",
         11660 => x"2eaf3882",
         11661 => x"cc942251",
         11662 => x"72712e9c",
         11663 => x"38811270",
         11664 => x"83ffff06",
         11665 => x"53517180",
         11666 => x"ff268d38",
         11667 => x"711082cc",
         11668 => x"94057022",
         11669 => x"5151e139",
         11670 => x"81801270",
         11671 => x"81ff0653",
         11672 => x"517182d8",
         11673 => x"c80c853d",
         11674 => x"0d04fe3d",
         11675 => x"0d029205",
         11676 => x"22028405",
         11677 => x"96052253",
         11678 => x"51805370",
         11679 => x"80ff2685",
         11680 => x"3870539a",
         11681 => x"397183b5",
         11682 => x"2e098106",
         11683 => x"91387081",
         11684 => x"ff268b38",
         11685 => x"701082ca",
         11686 => x"94057022",
         11687 => x"54517282",
         11688 => x"d8c80c84",
         11689 => x"3d0d04fb",
         11690 => x"3d0d7751",
         11691 => x"7083ffff",
         11692 => x"2681a738",
         11693 => x"7083ffff",
         11694 => x"0682ce94",
         11695 => x"57529fff",
         11696 => x"72278538",
         11697 => x"82d28856",
         11698 => x"75708205",
         11699 => x"57227030",
         11700 => x"70802572",
         11701 => x"75260751",
         11702 => x"52557080",
         11703 => x"fb387570",
         11704 => x"82055722",
         11705 => x"70882a71",
         11706 => x"81ff0670",
         11707 => x"18545255",
         11708 => x"53717125",
         11709 => x"80d73873",
         11710 => x"882680dc",
         11711 => x"38738429",
         11712 => x"82b0b005",
         11713 => x"51700804",
         11714 => x"71753110",
         11715 => x"76117022",
         11716 => x"54515180",
         11717 => x"c3397175",
         11718 => x"31810672",
         11719 => x"71315151",
         11720 => x"a439f012",
         11721 => x"519f39e0",
         11722 => x"12519a39",
         11723 => x"d0125195",
         11724 => x"39e61251",
         11725 => x"90398812",
         11726 => x"518b39ff",
         11727 => x"b0125185",
         11728 => x"39c7a012",
         11729 => x"517083ff",
         11730 => x"ff06528c",
         11731 => x"3973fef8",
         11732 => x"38721016",
         11733 => x"56fef139",
         11734 => x"71517082",
         11735 => x"d8c80c87",
         11736 => x"3d0d0400",
         11737 => x"00ffffff",
         11738 => x"ff00ffff",
         11739 => x"ffff00ff",
         11740 => x"ffffff00",
         11741 => x"00002baa",
         11742 => x"00002b2e",
         11743 => x"00002b35",
         11744 => x"00002b3c",
         11745 => x"00002b43",
         11746 => x"00002b4a",
         11747 => x"00002b51",
         11748 => x"00002b58",
         11749 => x"00002b5f",
         11750 => x"00002b66",
         11751 => x"00002b6d",
         11752 => x"00002b74",
         11753 => x"00002b7a",
         11754 => x"00002b80",
         11755 => x"00002b86",
         11756 => x"00002b8c",
         11757 => x"00002b92",
         11758 => x"00002b98",
         11759 => x"00002b9e",
         11760 => x"00002ba4",
         11761 => x"000043a6",
         11762 => x"000043ac",
         11763 => x"000043b2",
         11764 => x"000043b8",
         11765 => x"000043be",
         11766 => x"000049dd",
         11767 => x"00004add",
         11768 => x"00004bee",
         11769 => x"00004e46",
         11770 => x"00004ac5",
         11771 => x"000048b2",
         11772 => x"00004cb6",
         11773 => x"00004e17",
         11774 => x"00004cf9",
         11775 => x"00004d8f",
         11776 => x"00004d15",
         11777 => x"00004b98",
         11778 => x"000048b2",
         11779 => x"00004bee",
         11780 => x"00004c17",
         11781 => x"00004cb6",
         11782 => x"000048b2",
         11783 => x"000048b2",
         11784 => x"00004d15",
         11785 => x"00004d8f",
         11786 => x"00004e17",
         11787 => x"00004e46",
         11788 => x"00009708",
         11789 => x"00009716",
         11790 => x"00009722",
         11791 => x"00009727",
         11792 => x"0000972c",
         11793 => x"00009731",
         11794 => x"00009736",
         11795 => x"0000973b",
         11796 => x"00009741",
         11797 => x"00000e31",
         11798 => x"0000171a",
         11799 => x"0000171a",
         11800 => x"00000e60",
         11801 => x"0000171a",
         11802 => x"0000171a",
         11803 => x"0000171a",
         11804 => x"0000171a",
         11805 => x"0000171a",
         11806 => x"0000171a",
         11807 => x"0000171a",
         11808 => x"00000e1d",
         11809 => x"0000171a",
         11810 => x"00000e48",
         11811 => x"00000e78",
         11812 => x"0000171a",
         11813 => x"0000171a",
         11814 => x"0000171a",
         11815 => x"0000171a",
         11816 => x"0000171a",
         11817 => x"0000171a",
         11818 => x"0000171a",
         11819 => x"0000171a",
         11820 => x"0000171a",
         11821 => x"0000171a",
         11822 => x"0000171a",
         11823 => x"0000171a",
         11824 => x"0000171a",
         11825 => x"0000171a",
         11826 => x"0000171a",
         11827 => x"0000171a",
         11828 => x"0000171a",
         11829 => x"0000171a",
         11830 => x"0000171a",
         11831 => x"0000171a",
         11832 => x"0000171a",
         11833 => x"0000171a",
         11834 => x"0000171a",
         11835 => x"0000171a",
         11836 => x"0000171a",
         11837 => x"0000171a",
         11838 => x"0000171a",
         11839 => x"0000171a",
         11840 => x"0000171a",
         11841 => x"0000171a",
         11842 => x"0000171a",
         11843 => x"0000171a",
         11844 => x"0000171a",
         11845 => x"0000171a",
         11846 => x"0000171a",
         11847 => x"0000171a",
         11848 => x"00000fa8",
         11849 => x"0000171a",
         11850 => x"0000171a",
         11851 => x"0000171a",
         11852 => x"0000171a",
         11853 => x"00001116",
         11854 => x"0000171a",
         11855 => x"0000171a",
         11856 => x"0000171a",
         11857 => x"0000171a",
         11858 => x"0000171a",
         11859 => x"0000171a",
         11860 => x"0000171a",
         11861 => x"0000171a",
         11862 => x"0000171a",
         11863 => x"0000171a",
         11864 => x"00000ed8",
         11865 => x"0000103f",
         11866 => x"00000eaf",
         11867 => x"00000eaf",
         11868 => x"00000eaf",
         11869 => x"0000171a",
         11870 => x"0000103f",
         11871 => x"0000171a",
         11872 => x"0000171a",
         11873 => x"00000e98",
         11874 => x"0000171a",
         11875 => x"0000171a",
         11876 => x"000010ec",
         11877 => x"000010f7",
         11878 => x"0000171a",
         11879 => x"0000171a",
         11880 => x"00000f11",
         11881 => x"0000171a",
         11882 => x"0000111f",
         11883 => x"0000171a",
         11884 => x"0000171a",
         11885 => x"00001116",
         11886 => x"64696e69",
         11887 => x"74000000",
         11888 => x"64696f63",
         11889 => x"746c0000",
         11890 => x"66696e69",
         11891 => x"74000000",
         11892 => x"666c6f61",
         11893 => x"64000000",
         11894 => x"66657865",
         11895 => x"63000000",
         11896 => x"6d636c65",
         11897 => x"61720000",
         11898 => x"6d636f70",
         11899 => x"79000000",
         11900 => x"6d646966",
         11901 => x"66000000",
         11902 => x"6d64756d",
         11903 => x"70000000",
         11904 => x"6d656200",
         11905 => x"6d656800",
         11906 => x"6d657700",
         11907 => x"68696400",
         11908 => x"68696500",
         11909 => x"68666400",
         11910 => x"68666500",
         11911 => x"63616c6c",
         11912 => x"00000000",
         11913 => x"6a6d7000",
         11914 => x"72657374",
         11915 => x"61727400",
         11916 => x"72657365",
         11917 => x"74000000",
         11918 => x"696e666f",
         11919 => x"00000000",
         11920 => x"74657374",
         11921 => x"00000000",
         11922 => x"74626173",
         11923 => x"69630000",
         11924 => x"6d626173",
         11925 => x"69630000",
         11926 => x"6b696c6f",
         11927 => x"00000000",
         11928 => x"65640000",
         11929 => x"4469736b",
         11930 => x"20457272",
         11931 => x"6f720000",
         11932 => x"496e7465",
         11933 => x"726e616c",
         11934 => x"20657272",
         11935 => x"6f722e00",
         11936 => x"4469736b",
         11937 => x"206e6f74",
         11938 => x"20726561",
         11939 => x"64792e00",
         11940 => x"4e6f2066",
         11941 => x"696c6520",
         11942 => x"666f756e",
         11943 => x"642e0000",
         11944 => x"4e6f2070",
         11945 => x"61746820",
         11946 => x"666f756e",
         11947 => x"642e0000",
         11948 => x"496e7661",
         11949 => x"6c696420",
         11950 => x"66696c65",
         11951 => x"6e616d65",
         11952 => x"2e000000",
         11953 => x"41636365",
         11954 => x"73732064",
         11955 => x"656e6965",
         11956 => x"642e0000",
         11957 => x"46696c65",
         11958 => x"20616c72",
         11959 => x"65616479",
         11960 => x"20657869",
         11961 => x"7374732e",
         11962 => x"00000000",
         11963 => x"46696c65",
         11964 => x"2068616e",
         11965 => x"646c6520",
         11966 => x"696e7661",
         11967 => x"6c69642e",
         11968 => x"00000000",
         11969 => x"53442069",
         11970 => x"73207772",
         11971 => x"69746520",
         11972 => x"70726f74",
         11973 => x"65637465",
         11974 => x"642e0000",
         11975 => x"44726976",
         11976 => x"65206e75",
         11977 => x"6d626572",
         11978 => x"20697320",
         11979 => x"696e7661",
         11980 => x"6c69642e",
         11981 => x"00000000",
         11982 => x"4469736b",
         11983 => x"206e6f74",
         11984 => x"20656e61",
         11985 => x"626c6564",
         11986 => x"2e000000",
         11987 => x"4e6f2063",
         11988 => x"6f6d7061",
         11989 => x"7469626c",
         11990 => x"65206669",
         11991 => x"6c657379",
         11992 => x"7374656d",
         11993 => x"20666f75",
         11994 => x"6e64206f",
         11995 => x"6e206469",
         11996 => x"736b2e00",
         11997 => x"466f726d",
         11998 => x"61742061",
         11999 => x"626f7274",
         12000 => x"65642e00",
         12001 => x"54696d65",
         12002 => x"6f75742c",
         12003 => x"206f7065",
         12004 => x"72617469",
         12005 => x"6f6e2063",
         12006 => x"616e6365",
         12007 => x"6c6c6564",
         12008 => x"2e000000",
         12009 => x"46696c65",
         12010 => x"20697320",
         12011 => x"6c6f636b",
         12012 => x"65642e00",
         12013 => x"496e7375",
         12014 => x"66666963",
         12015 => x"69656e74",
         12016 => x"206d656d",
         12017 => x"6f72792e",
         12018 => x"00000000",
         12019 => x"546f6f20",
         12020 => x"6d616e79",
         12021 => x"206f7065",
         12022 => x"6e206669",
         12023 => x"6c65732e",
         12024 => x"00000000",
         12025 => x"50617261",
         12026 => x"6d657465",
         12027 => x"72732069",
         12028 => x"6e636f72",
         12029 => x"72656374",
         12030 => x"2e000000",
         12031 => x"53756363",
         12032 => x"6573732e",
         12033 => x"00000000",
         12034 => x"556e6b6e",
         12035 => x"6f776e20",
         12036 => x"6572726f",
         12037 => x"722e0000",
         12038 => x"0a256c75",
         12039 => x"20627974",
         12040 => x"65732025",
         12041 => x"73206174",
         12042 => x"20256c75",
         12043 => x"20627974",
         12044 => x"65732f73",
         12045 => x"65632e0a",
         12046 => x"00000000",
         12047 => x"72656164",
         12048 => x"00000000",
         12049 => x"303d2530",
         12050 => x"386c782c",
         12051 => x"20313d25",
         12052 => x"30386c78",
         12053 => x"2c20323d",
         12054 => x"2530386c",
         12055 => x"782c205f",
         12056 => x"494f423d",
         12057 => x"2530386c",
         12058 => x"78202530",
         12059 => x"386c7820",
         12060 => x"2530386c",
         12061 => x"780a0000",
         12062 => x"2530386c",
         12063 => x"58000000",
         12064 => x"3a202000",
         12065 => x"25303458",
         12066 => x"00000000",
         12067 => x"20202020",
         12068 => x"20202020",
         12069 => x"00000000",
         12070 => x"25303258",
         12071 => x"00000000",
         12072 => x"20200000",
         12073 => x"207c0000",
         12074 => x"7c000000",
         12075 => x"5a505554",
         12076 => x"41000000",
         12077 => x"0a2a2a20",
         12078 => x"25732028",
         12079 => x"00000000",
         12080 => x"30322f30",
         12081 => x"352f3230",
         12082 => x"32300000",
         12083 => x"76312e35",
         12084 => x"32000000",
         12085 => x"205a5055",
         12086 => x"2c207265",
         12087 => x"76202530",
         12088 => x"32782920",
         12089 => x"25732025",
         12090 => x"73202a2a",
         12091 => x"0a0a0000",
         12092 => x"5a505554",
         12093 => x"4120496e",
         12094 => x"74657272",
         12095 => x"75707420",
         12096 => x"48616e64",
         12097 => x"6c657200",
         12098 => x"54696d65",
         12099 => x"7220696e",
         12100 => x"74657272",
         12101 => x"75707400",
         12102 => x"50533220",
         12103 => x"696e7465",
         12104 => x"72727570",
         12105 => x"74000000",
         12106 => x"494f4354",
         12107 => x"4c205244",
         12108 => x"20696e74",
         12109 => x"65727275",
         12110 => x"70740000",
         12111 => x"494f4354",
         12112 => x"4c205752",
         12113 => x"20696e74",
         12114 => x"65727275",
         12115 => x"70740000",
         12116 => x"55415254",
         12117 => x"30205258",
         12118 => x"20696e74",
         12119 => x"65727275",
         12120 => x"70740000",
         12121 => x"55415254",
         12122 => x"30205458",
         12123 => x"20696e74",
         12124 => x"65727275",
         12125 => x"70740000",
         12126 => x"55415254",
         12127 => x"31205258",
         12128 => x"20696e74",
         12129 => x"65727275",
         12130 => x"70740000",
         12131 => x"55415254",
         12132 => x"31205458",
         12133 => x"20696e74",
         12134 => x"65727275",
         12135 => x"70740000",
         12136 => x"53657474",
         12137 => x"696e6720",
         12138 => x"75702074",
         12139 => x"696d6572",
         12140 => x"2e2e2e00",
         12141 => x"456e6162",
         12142 => x"6c696e67",
         12143 => x"2074696d",
         12144 => x"65722e2e",
         12145 => x"2e000000",
         12146 => x"6175746f",
         12147 => x"65786563",
         12148 => x"2e626174",
         12149 => x"00000000",
         12150 => x"7a707574",
         12151 => x"612e6873",
         12152 => x"74000000",
         12153 => x"303a0000",
         12154 => x"4661696c",
         12155 => x"65642074",
         12156 => x"6f20696e",
         12157 => x"69746961",
         12158 => x"6c697365",
         12159 => x"20736420",
         12160 => x"63617264",
         12161 => x"20302c20",
         12162 => x"706c6561",
         12163 => x"73652069",
         12164 => x"6e697420",
         12165 => x"6d616e75",
         12166 => x"616c6c79",
         12167 => x"2e000000",
         12168 => x"2a200000",
         12169 => x"42616420",
         12170 => x"6469736b",
         12171 => x"20696421",
         12172 => x"00000000",
         12173 => x"496e6974",
         12174 => x"69616c69",
         12175 => x"7365642e",
         12176 => x"00000000",
         12177 => x"4661696c",
         12178 => x"65642074",
         12179 => x"6f20696e",
         12180 => x"69746961",
         12181 => x"6c697365",
         12182 => x"2e000000",
         12183 => x"72633d25",
         12184 => x"640a0000",
         12185 => x"25753a00",
         12186 => x"436c6561",
         12187 => x"72696e67",
         12188 => x"2e2e2e2e",
         12189 => x"00000000",
         12190 => x"436f7079",
         12191 => x"696e672e",
         12192 => x"2e2e0000",
         12193 => x"436f6d70",
         12194 => x"6172696e",
         12195 => x"672e2e2e",
         12196 => x"00000000",
         12197 => x"2530386c",
         12198 => x"78282530",
         12199 => x"3878292d",
         12200 => x"3e253038",
         12201 => x"6c782825",
         12202 => x"30387829",
         12203 => x"0a000000",
         12204 => x"44756d70",
         12205 => x"204d656d",
         12206 => x"6f727900",
         12207 => x"0a436f6d",
         12208 => x"706c6574",
         12209 => x"652e0000",
         12210 => x"2530386c",
         12211 => x"58202530",
         12212 => x"32582d00",
         12213 => x"3f3f3f00",
         12214 => x"2530386c",
         12215 => x"58202530",
         12216 => x"34582d00",
         12217 => x"2530386c",
         12218 => x"58202530",
         12219 => x"386c582d",
         12220 => x"00000000",
         12221 => x"44697361",
         12222 => x"626c696e",
         12223 => x"6720696e",
         12224 => x"74657272",
         12225 => x"75707473",
         12226 => x"00000000",
         12227 => x"456e6162",
         12228 => x"6c696e67",
         12229 => x"20696e74",
         12230 => x"65727275",
         12231 => x"70747300",
         12232 => x"44697361",
         12233 => x"626c6564",
         12234 => x"20756172",
         12235 => x"74206669",
         12236 => x"666f0000",
         12237 => x"456e6162",
         12238 => x"6c696e67",
         12239 => x"20756172",
         12240 => x"74206669",
         12241 => x"666f0000",
         12242 => x"45786563",
         12243 => x"7574696e",
         12244 => x"6720636f",
         12245 => x"64652040",
         12246 => x"20253038",
         12247 => x"6c78202e",
         12248 => x"2e2e0a00",
         12249 => x"43616c6c",
         12250 => x"696e6720",
         12251 => x"636f6465",
         12252 => x"20402025",
         12253 => x"30386c78",
         12254 => x"202e2e2e",
         12255 => x"0a000000",
         12256 => x"43616c6c",
         12257 => x"20726574",
         12258 => x"75726e65",
         12259 => x"6420636f",
         12260 => x"64652028",
         12261 => x"2564292e",
         12262 => x"0a000000",
         12263 => x"52657374",
         12264 => x"61727469",
         12265 => x"6e672061",
         12266 => x"70706c69",
         12267 => x"63617469",
         12268 => x"6f6e2e2e",
         12269 => x"2e000000",
         12270 => x"436f6c64",
         12271 => x"20726562",
         12272 => x"6f6f7469",
         12273 => x"6e672e2e",
         12274 => x"2e000000",
         12275 => x"5a505500",
         12276 => x"62696e00",
         12277 => x"25643a5c",
         12278 => x"25735c25",
         12279 => x"732e2573",
         12280 => x"00000000",
         12281 => x"25643a5c",
         12282 => x"25735c25",
         12283 => x"73000000",
         12284 => x"25643a5c",
         12285 => x"25730000",
         12286 => x"42616420",
         12287 => x"636f6d6d",
         12288 => x"616e642e",
         12289 => x"00000000",
         12290 => x"52756e6e",
         12291 => x"696e672e",
         12292 => x"2e2e0000",
         12293 => x"456e6162",
         12294 => x"6c696e67",
         12295 => x"20696e74",
         12296 => x"65727275",
         12297 => x"7074732e",
         12298 => x"2e2e0000",
         12299 => x"25642f25",
         12300 => x"642f2564",
         12301 => x"2025643a",
         12302 => x"25643a25",
         12303 => x"642e2564",
         12304 => x"25640a00",
         12305 => x"536f4320",
         12306 => x"436f6e66",
         12307 => x"69677572",
         12308 => x"6174696f",
         12309 => x"6e000000",
         12310 => x"20286672",
         12311 => x"6f6d2053",
         12312 => x"6f432063",
         12313 => x"6f6e6669",
         12314 => x"67290000",
         12315 => x"3a0a4465",
         12316 => x"76696365",
         12317 => x"7320696d",
         12318 => x"706c656d",
         12319 => x"656e7465",
         12320 => x"643a0000",
         12321 => x"20202020",
         12322 => x"57422053",
         12323 => x"4452414d",
         12324 => x"20202825",
         12325 => x"3038583a",
         12326 => x"25303858",
         12327 => x"292e0a00",
         12328 => x"20202020",
         12329 => x"53445241",
         12330 => x"4d202020",
         12331 => x"20202825",
         12332 => x"3038583a",
         12333 => x"25303858",
         12334 => x"292e0a00",
         12335 => x"20202020",
         12336 => x"494e534e",
         12337 => x"20425241",
         12338 => x"4d202825",
         12339 => x"3038583a",
         12340 => x"25303858",
         12341 => x"292e0a00",
         12342 => x"20202020",
         12343 => x"4252414d",
         12344 => x"20202020",
         12345 => x"20202825",
         12346 => x"3038583a",
         12347 => x"25303858",
         12348 => x"292e0a00",
         12349 => x"20202020",
         12350 => x"52414d20",
         12351 => x"20202020",
         12352 => x"20202825",
         12353 => x"3038583a",
         12354 => x"25303858",
         12355 => x"292e0a00",
         12356 => x"20202020",
         12357 => x"53442043",
         12358 => x"41524420",
         12359 => x"20202844",
         12360 => x"65766963",
         12361 => x"6573203d",
         12362 => x"25303264",
         12363 => x"292e0a00",
         12364 => x"20202020",
         12365 => x"54494d45",
         12366 => x"52312020",
         12367 => x"20202854",
         12368 => x"696d6572",
         12369 => x"7320203d",
         12370 => x"25303264",
         12371 => x"292e0a00",
         12372 => x"20202020",
         12373 => x"494e5452",
         12374 => x"20435452",
         12375 => x"4c202843",
         12376 => x"68616e6e",
         12377 => x"656c733d",
         12378 => x"25303264",
         12379 => x"292e0a00",
         12380 => x"20202020",
         12381 => x"57495348",
         12382 => x"424f4e45",
         12383 => x"20425553",
         12384 => x"00000000",
         12385 => x"20202020",
         12386 => x"57422049",
         12387 => x"32430000",
         12388 => x"20202020",
         12389 => x"494f4354",
         12390 => x"4c000000",
         12391 => x"20202020",
         12392 => x"50533200",
         12393 => x"20202020",
         12394 => x"53504900",
         12395 => x"41646472",
         12396 => x"65737365",
         12397 => x"733a0000",
         12398 => x"20202020",
         12399 => x"43505520",
         12400 => x"52657365",
         12401 => x"74205665",
         12402 => x"63746f72",
         12403 => x"20416464",
         12404 => x"72657373",
         12405 => x"203d2025",
         12406 => x"3038580a",
         12407 => x"00000000",
         12408 => x"20202020",
         12409 => x"43505520",
         12410 => x"4d656d6f",
         12411 => x"72792053",
         12412 => x"74617274",
         12413 => x"20416464",
         12414 => x"72657373",
         12415 => x"203d2025",
         12416 => x"3038580a",
         12417 => x"00000000",
         12418 => x"20202020",
         12419 => x"53746163",
         12420 => x"6b205374",
         12421 => x"61727420",
         12422 => x"41646472",
         12423 => x"65737320",
         12424 => x"20202020",
         12425 => x"203d2025",
         12426 => x"3038580a",
         12427 => x"00000000",
         12428 => x"4d697363",
         12429 => x"3a000000",
         12430 => x"20202020",
         12431 => x"5a505520",
         12432 => x"49642020",
         12433 => x"20202020",
         12434 => x"20202020",
         12435 => x"20202020",
         12436 => x"20202020",
         12437 => x"203d2025",
         12438 => x"3034580a",
         12439 => x"00000000",
         12440 => x"20202020",
         12441 => x"53797374",
         12442 => x"656d2043",
         12443 => x"6c6f636b",
         12444 => x"20467265",
         12445 => x"71202020",
         12446 => x"20202020",
         12447 => x"203d2025",
         12448 => x"642e2530",
         12449 => x"34644d48",
         12450 => x"7a0a0000",
         12451 => x"20202020",
         12452 => x"53445241",
         12453 => x"4d20436c",
         12454 => x"6f636b20",
         12455 => x"46726571",
         12456 => x"20202020",
         12457 => x"20202020",
         12458 => x"203d2025",
         12459 => x"642e2530",
         12460 => x"34644d48",
         12461 => x"7a0a0000",
         12462 => x"20202020",
         12463 => x"57697368",
         12464 => x"626f6e65",
         12465 => x"20534452",
         12466 => x"414d2043",
         12467 => x"6c6f636b",
         12468 => x"20467265",
         12469 => x"713d2025",
         12470 => x"642e2530",
         12471 => x"34644d48",
         12472 => x"7a0a0000",
         12473 => x"536d616c",
         12474 => x"6c000000",
         12475 => x"4d656469",
         12476 => x"756d0000",
         12477 => x"466c6578",
         12478 => x"00000000",
         12479 => x"45564f00",
         12480 => x"45564f6d",
         12481 => x"00000000",
         12482 => x"556e6b6e",
         12483 => x"6f776e00",
         12484 => x"0000a46c",
         12485 => x"01000000",
         12486 => x"00000002",
         12487 => x"0000a468",
         12488 => x"01000000",
         12489 => x"00000003",
         12490 => x"0000a464",
         12491 => x"01000000",
         12492 => x"00000004",
         12493 => x"0000a460",
         12494 => x"01000000",
         12495 => x"00000005",
         12496 => x"0000a45c",
         12497 => x"01000000",
         12498 => x"00000006",
         12499 => x"0000a458",
         12500 => x"01000000",
         12501 => x"00000007",
         12502 => x"0000a454",
         12503 => x"01000000",
         12504 => x"00000001",
         12505 => x"0000a450",
         12506 => x"01000000",
         12507 => x"00000008",
         12508 => x"0000a44c",
         12509 => x"01000000",
         12510 => x"0000000b",
         12511 => x"0000a448",
         12512 => x"01000000",
         12513 => x"00000009",
         12514 => x"0000a444",
         12515 => x"01000000",
         12516 => x"0000000a",
         12517 => x"0000a440",
         12518 => x"04000000",
         12519 => x"0000000d",
         12520 => x"0000a43c",
         12521 => x"04000000",
         12522 => x"0000000c",
         12523 => x"0000a438",
         12524 => x"04000000",
         12525 => x"0000000e",
         12526 => x"0000a434",
         12527 => x"03000000",
         12528 => x"0000000f",
         12529 => x"0000a430",
         12530 => x"04000000",
         12531 => x"0000000f",
         12532 => x"0000a42c",
         12533 => x"04000000",
         12534 => x"00000010",
         12535 => x"0000a428",
         12536 => x"04000000",
         12537 => x"00000011",
         12538 => x"0000a424",
         12539 => x"03000000",
         12540 => x"00000012",
         12541 => x"0000a420",
         12542 => x"03000000",
         12543 => x"00000013",
         12544 => x"0000a41c",
         12545 => x"03000000",
         12546 => x"00000014",
         12547 => x"0000a418",
         12548 => x"03000000",
         12549 => x"00000015",
         12550 => x"1b5b4400",
         12551 => x"1b5b4300",
         12552 => x"1b5b4200",
         12553 => x"1b5b4100",
         12554 => x"1b5b367e",
         12555 => x"1b5b357e",
         12556 => x"1b5b347e",
         12557 => x"1b304600",
         12558 => x"1b5b337e",
         12559 => x"1b5b327e",
         12560 => x"1b5b317e",
         12561 => x"10000000",
         12562 => x"0e000000",
         12563 => x"0d000000",
         12564 => x"0b000000",
         12565 => x"08000000",
         12566 => x"06000000",
         12567 => x"05000000",
         12568 => x"04000000",
         12569 => x"03000000",
         12570 => x"02000000",
         12571 => x"01000000",
         12572 => x"68697374",
         12573 => x"6f727900",
         12574 => x"68697374",
         12575 => x"00000000",
         12576 => x"21000000",
         12577 => x"2530346c",
         12578 => x"75202025",
         12579 => x"730a0000",
         12580 => x"4661696c",
         12581 => x"65642074",
         12582 => x"6f207265",
         12583 => x"73657420",
         12584 => x"74686520",
         12585 => x"68697374",
         12586 => x"6f727920",
         12587 => x"66696c65",
         12588 => x"20746f20",
         12589 => x"454f462e",
         12590 => x"00000000",
         12591 => x"43616e6e",
         12592 => x"6f74206f",
         12593 => x"70656e2f",
         12594 => x"63726561",
         12595 => x"74652068",
         12596 => x"6973746f",
         12597 => x"72792066",
         12598 => x"696c652c",
         12599 => x"20646973",
         12600 => x"61626c69",
         12601 => x"6e672e00",
         12602 => x"53440000",
         12603 => x"222a3a3c",
         12604 => x"3e3f7c7f",
         12605 => x"00000000",
         12606 => x"2b2c3b3d",
         12607 => x"5b5d0000",
         12608 => x"46415400",
         12609 => x"46415433",
         12610 => x"32000000",
         12611 => x"ebfe904d",
         12612 => x"53444f53",
         12613 => x"352e3000",
         12614 => x"4e4f204e",
         12615 => x"414d4520",
         12616 => x"20202046",
         12617 => x"41543332",
         12618 => x"20202000",
         12619 => x"4e4f204e",
         12620 => x"414d4520",
         12621 => x"20202046",
         12622 => x"41542020",
         12623 => x"20202000",
         12624 => x"0000a4e8",
         12625 => x"00000000",
         12626 => x"00000000",
         12627 => x"00000000",
         12628 => x"01030507",
         12629 => x"090e1012",
         12630 => x"1416181c",
         12631 => x"1e000000",
         12632 => x"809a4541",
         12633 => x"8e418f80",
         12634 => x"45454549",
         12635 => x"49498e8f",
         12636 => x"9092924f",
         12637 => x"994f5555",
         12638 => x"59999a9b",
         12639 => x"9c9d9e9f",
         12640 => x"41494f55",
         12641 => x"a5a5a6a7",
         12642 => x"a8a9aaab",
         12643 => x"acadaeaf",
         12644 => x"b0b1b2b3",
         12645 => x"b4b5b6b7",
         12646 => x"b8b9babb",
         12647 => x"bcbdbebf",
         12648 => x"c0c1c2c3",
         12649 => x"c4c5c6c7",
         12650 => x"c8c9cacb",
         12651 => x"cccdcecf",
         12652 => x"d0d1d2d3",
         12653 => x"d4d5d6d7",
         12654 => x"d8d9dadb",
         12655 => x"dcdddedf",
         12656 => x"e0e1e2e3",
         12657 => x"e4e5e6e7",
         12658 => x"e8e9eaeb",
         12659 => x"ecedeeef",
         12660 => x"f0f1f2f3",
         12661 => x"f4f5f6f7",
         12662 => x"f8f9fafb",
         12663 => x"fcfdfeff",
         12664 => x"2b2e2c3b",
         12665 => x"3d5b5d2f",
         12666 => x"5c222a3a",
         12667 => x"3c3e3f7c",
         12668 => x"7f000000",
         12669 => x"00010004",
         12670 => x"00100040",
         12671 => x"01000200",
         12672 => x"00000000",
         12673 => x"00010002",
         12674 => x"00040008",
         12675 => x"00100020",
         12676 => x"00000000",
         12677 => x"00c700fc",
         12678 => x"00e900e2",
         12679 => x"00e400e0",
         12680 => x"00e500e7",
         12681 => x"00ea00eb",
         12682 => x"00e800ef",
         12683 => x"00ee00ec",
         12684 => x"00c400c5",
         12685 => x"00c900e6",
         12686 => x"00c600f4",
         12687 => x"00f600f2",
         12688 => x"00fb00f9",
         12689 => x"00ff00d6",
         12690 => x"00dc00a2",
         12691 => x"00a300a5",
         12692 => x"20a70192",
         12693 => x"00e100ed",
         12694 => x"00f300fa",
         12695 => x"00f100d1",
         12696 => x"00aa00ba",
         12697 => x"00bf2310",
         12698 => x"00ac00bd",
         12699 => x"00bc00a1",
         12700 => x"00ab00bb",
         12701 => x"25912592",
         12702 => x"25932502",
         12703 => x"25242561",
         12704 => x"25622556",
         12705 => x"25552563",
         12706 => x"25512557",
         12707 => x"255d255c",
         12708 => x"255b2510",
         12709 => x"25142534",
         12710 => x"252c251c",
         12711 => x"2500253c",
         12712 => x"255e255f",
         12713 => x"255a2554",
         12714 => x"25692566",
         12715 => x"25602550",
         12716 => x"256c2567",
         12717 => x"25682564",
         12718 => x"25652559",
         12719 => x"25582552",
         12720 => x"2553256b",
         12721 => x"256a2518",
         12722 => x"250c2588",
         12723 => x"2584258c",
         12724 => x"25902580",
         12725 => x"03b100df",
         12726 => x"039303c0",
         12727 => x"03a303c3",
         12728 => x"00b503c4",
         12729 => x"03a60398",
         12730 => x"03a903b4",
         12731 => x"221e03c6",
         12732 => x"03b52229",
         12733 => x"226100b1",
         12734 => x"22652264",
         12735 => x"23202321",
         12736 => x"00f72248",
         12737 => x"00b02219",
         12738 => x"00b7221a",
         12739 => x"207f00b2",
         12740 => x"25a000a0",
         12741 => x"0061031a",
         12742 => x"00e00317",
         12743 => x"00f80307",
         12744 => x"00ff0001",
         12745 => x"01780100",
         12746 => x"01300132",
         12747 => x"01060139",
         12748 => x"0110014a",
         12749 => x"012e0179",
         12750 => x"01060180",
         12751 => x"004d0243",
         12752 => x"01810182",
         12753 => x"01820184",
         12754 => x"01840186",
         12755 => x"01870187",
         12756 => x"0189018a",
         12757 => x"018b018b",
         12758 => x"018d018e",
         12759 => x"018f0190",
         12760 => x"01910191",
         12761 => x"01930194",
         12762 => x"01f60196",
         12763 => x"01970198",
         12764 => x"0198023d",
         12765 => x"019b019c",
         12766 => x"019d0220",
         12767 => x"019f01a0",
         12768 => x"01a001a2",
         12769 => x"01a201a4",
         12770 => x"01a401a6",
         12771 => x"01a701a7",
         12772 => x"01a901aa",
         12773 => x"01ab01ac",
         12774 => x"01ac01ae",
         12775 => x"01af01af",
         12776 => x"01b101b2",
         12777 => x"01b301b3",
         12778 => x"01b501b5",
         12779 => x"01b701b8",
         12780 => x"01b801ba",
         12781 => x"01bb01bc",
         12782 => x"01bc01be",
         12783 => x"01f701c0",
         12784 => x"01c101c2",
         12785 => x"01c301c4",
         12786 => x"01c501c4",
         12787 => x"01c701c8",
         12788 => x"01c701ca",
         12789 => x"01cb01ca",
         12790 => x"01cd0110",
         12791 => x"01dd0001",
         12792 => x"018e01de",
         12793 => x"011201f3",
         12794 => x"000301f1",
         12795 => x"01f401f4",
         12796 => x"01f80128",
         12797 => x"02220112",
         12798 => x"023a0009",
         12799 => x"2c65023b",
         12800 => x"023b023d",
         12801 => x"2c66023f",
         12802 => x"02400241",
         12803 => x"02410246",
         12804 => x"010a0253",
         12805 => x"00400181",
         12806 => x"01860255",
         12807 => x"0189018a",
         12808 => x"0258018f",
         12809 => x"025a0190",
         12810 => x"025c025d",
         12811 => x"025e025f",
         12812 => x"01930261",
         12813 => x"02620194",
         12814 => x"02640265",
         12815 => x"02660267",
         12816 => x"01970196",
         12817 => x"026a2c62",
         12818 => x"026c026d",
         12819 => x"026e019c",
         12820 => x"02700271",
         12821 => x"019d0273",
         12822 => x"0274019f",
         12823 => x"02760277",
         12824 => x"02780279",
         12825 => x"027a027b",
         12826 => x"027c2c64",
         12827 => x"027e027f",
         12828 => x"01a60281",
         12829 => x"028201a9",
         12830 => x"02840285",
         12831 => x"02860287",
         12832 => x"01ae0244",
         12833 => x"01b101b2",
         12834 => x"0245028d",
         12835 => x"028e028f",
         12836 => x"02900291",
         12837 => x"01b7037b",
         12838 => x"000303fd",
         12839 => x"03fe03ff",
         12840 => x"03ac0004",
         12841 => x"03860388",
         12842 => x"0389038a",
         12843 => x"03b10311",
         12844 => x"03c20002",
         12845 => x"03a303a3",
         12846 => x"03c40308",
         12847 => x"03cc0003",
         12848 => x"038c038e",
         12849 => x"038f03d8",
         12850 => x"011803f2",
         12851 => x"000a03f9",
         12852 => x"03f303f4",
         12853 => x"03f503f6",
         12854 => x"03f703f7",
         12855 => x"03f903fa",
         12856 => x"03fa0430",
         12857 => x"03200450",
         12858 => x"07100460",
         12859 => x"0122048a",
         12860 => x"013604c1",
         12861 => x"010e04cf",
         12862 => x"000104c0",
         12863 => x"04d00144",
         12864 => x"05610426",
         12865 => x"00000000",
         12866 => x"1d7d0001",
         12867 => x"2c631e00",
         12868 => x"01961ea0",
         12869 => x"015a1f00",
         12870 => x"06081f10",
         12871 => x"06061f20",
         12872 => x"06081f30",
         12873 => x"06081f40",
         12874 => x"06061f51",
         12875 => x"00071f59",
         12876 => x"1f521f5b",
         12877 => x"1f541f5d",
         12878 => x"1f561f5f",
         12879 => x"1f600608",
         12880 => x"1f70000e",
         12881 => x"1fba1fbb",
         12882 => x"1fc81fc9",
         12883 => x"1fca1fcb",
         12884 => x"1fda1fdb",
         12885 => x"1ff81ff9",
         12886 => x"1fea1feb",
         12887 => x"1ffa1ffb",
         12888 => x"1f800608",
         12889 => x"1f900608",
         12890 => x"1fa00608",
         12891 => x"1fb00004",
         12892 => x"1fb81fb9",
         12893 => x"1fb21fbc",
         12894 => x"1fcc0001",
         12895 => x"1fc31fd0",
         12896 => x"06021fe0",
         12897 => x"06021fe5",
         12898 => x"00011fec",
         12899 => x"1ff30001",
         12900 => x"1ffc214e",
         12901 => x"00012132",
         12902 => x"21700210",
         12903 => x"21840001",
         12904 => x"218324d0",
         12905 => x"051a2c30",
         12906 => x"042f2c60",
         12907 => x"01022c67",
         12908 => x"01062c75",
         12909 => x"01022c80",
         12910 => x"01642d00",
         12911 => x"0826ff41",
         12912 => x"031a0000",
         12913 => x"00000000",
         12914 => x"000099b8",
         12915 => x"01020100",
         12916 => x"00000000",
         12917 => x"00000000",
         12918 => x"000099c0",
         12919 => x"01040100",
         12920 => x"00000000",
         12921 => x"00000000",
         12922 => x"000099c8",
         12923 => x"01140300",
         12924 => x"00000000",
         12925 => x"00000000",
         12926 => x"000099d0",
         12927 => x"012b0300",
         12928 => x"00000000",
         12929 => x"00000000",
         12930 => x"000099d8",
         12931 => x"01300300",
         12932 => x"00000000",
         12933 => x"00000000",
         12934 => x"000099e0",
         12935 => x"013c0400",
         12936 => x"00000000",
         12937 => x"00000000",
         12938 => x"000099e8",
         12939 => x"013d0400",
         12940 => x"00000000",
         12941 => x"00000000",
         12942 => x"000099f0",
         12943 => x"013f0400",
         12944 => x"00000000",
         12945 => x"00000000",
         12946 => x"000099f8",
         12947 => x"01400400",
         12948 => x"00000000",
         12949 => x"00000000",
         12950 => x"00009a00",
         12951 => x"01410400",
         12952 => x"00000000",
         12953 => x"00000000",
         12954 => x"00009a04",
         12955 => x"01420400",
         12956 => x"00000000",
         12957 => x"00000000",
         12958 => x"00009a08",
         12959 => x"01430400",
         12960 => x"00000000",
         12961 => x"00000000",
         12962 => x"00009a0c",
         12963 => x"01500500",
         12964 => x"00000000",
         12965 => x"00000000",
         12966 => x"00009a10",
         12967 => x"01510500",
         12968 => x"00000000",
         12969 => x"00000000",
         12970 => x"00009a14",
         12971 => x"01540500",
         12972 => x"00000000",
         12973 => x"00000000",
         12974 => x"00009a18",
         12975 => x"01550500",
         12976 => x"00000000",
         12977 => x"00000000",
         12978 => x"00009a1c",
         12979 => x"01790700",
         12980 => x"00000000",
         12981 => x"00000000",
         12982 => x"00009a24",
         12983 => x"01780700",
         12984 => x"00000000",
         12985 => x"00000000",
         12986 => x"00009a28",
         12987 => x"01820800",
         12988 => x"00000000",
         12989 => x"00000000",
         12990 => x"00009a30",
         12991 => x"01830800",
         12992 => x"00000000",
         12993 => x"00000000",
         12994 => x"00009a38",
         12995 => x"01850800",
         12996 => x"00000000",
         12997 => x"00000000",
         12998 => x"00009a40",
         12999 => x"01870800",
         13000 => x"00000000",
         13001 => x"00000000",
         13002 => x"00009a48",
         13003 => x"018c0900",
         13004 => x"00000000",
         13005 => x"00000000",
         13006 => x"00009a50",
         13007 => x"018d0900",
         13008 => x"00000000",
         13009 => x"00000000",
         13010 => x"00009a58",
         13011 => x"018e0900",
         13012 => x"00000000",
         13013 => x"00000000",
         13014 => x"00009a60",
         13015 => x"018f0900",
         13016 => x"00000000",
         13017 => x"00000000",
         13018 => x"00000000",
         13019 => x"00000000",
         13020 => x"00007fff",
         13021 => x"00000000",
         13022 => x"00007fff",
         13023 => x"00010000",
         13024 => x"00007fff",
         13025 => x"00010000",
         13026 => x"00810000",
         13027 => x"01000000",
         13028 => x"017fffff",
         13029 => x"00000000",
         13030 => x"00000000",
         13031 => x"00007800",
         13032 => x"00000000",
         13033 => x"05f5e100",
         13034 => x"05f5e100",
         13035 => x"05f5e100",
         13036 => x"00000000",
         13037 => x"01010101",
         13038 => x"01010101",
         13039 => x"01011001",
         13040 => x"01000000",
         13041 => x"00000000",
         13042 => x"00000000",
         13043 => x"00000000",
         13044 => x"00000000",
         13045 => x"00000000",
         13046 => x"00000000",
         13047 => x"00000000",
         13048 => x"00000000",
         13049 => x"00000000",
         13050 => x"00000000",
         13051 => x"00000000",
         13052 => x"00000000",
         13053 => x"00000000",
         13054 => x"00000000",
         13055 => x"00000000",
         13056 => x"00000000",
         13057 => x"00000000",
         13058 => x"00000000",
         13059 => x"00000000",
         13060 => x"00000000",
         13061 => x"00000000",
         13062 => x"00000000",
         13063 => x"00000000",
         13064 => x"00000000",
         13065 => x"0000a470",
         13066 => x"01000000",
         13067 => x"0000a478",
         13068 => x"01000000",
         13069 => x"0000a480",
         13070 => x"02000000",
         13071 => x"00000000",
         13072 => x"00000000",
         13073 => x"01000000",
        others => x"00000000"
    );

begin

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
            report "write collision" severity failure;
        end if;
    
        if (memAWriteEnable = '1') then
            ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE)))) := memAWrite;
            memARead <= memAWrite;
        else
            memARead <= ram(to_integer(unsigned(memAAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;

process (clk)
begin
    if (clk'event and clk = '1') then
        if (memBWriteEnable = '1') then
            ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE)))) := memBWrite;
            memBRead <= memBWrite;
        else
            memBRead <= ram(to_integer(unsigned(memBAddr(ADDR_32BIT_BRAM_RANGE))));
        end if;
    end if;
end process;


end arch;

