-- Byte Addressed 32bit BRAM module for the ZPU Evo implementation.
--
-- Copyright 2018-2019 - Philip Smart for the ZPU Evo implementation.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
library pkgs;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use pkgs.config_pkg.all;
use work.zpu_pkg.all;
use work.zpu_soc_pkg.all;

entity SinglePortBRAM is
    generic
    (
        addrbits             : integer := 16
    );
    port
    (
        clk                  : in  std_logic;
        memAAddr             : in  std_logic_vector(addrbits-1 downto 0);
        memAWriteEnable      : in  std_logic;
        memAWriteByte        : in  std_logic;
        memAWriteHalfWord    : in  std_logic;
        memAWrite            : in  std_logic_vector(WORD_32BIT_RANGE);
        memARead             : out std_logic_vector(WORD_32BIT_RANGE)
    );
end SinglePortBRAM;

architecture arch of SinglePortBRAM is

    type ramArray is array(natural range 0 to (2**(addrbits-2))-1) of std_logic_vector(7 downto 0);

    shared variable RAM0 : ramArray :=
    (
             0 => x"84",
             1 => x"0b",
             2 => x"04",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"84",
             9 => x"0b",
            10 => x"04",
            11 => x"84",
            12 => x"0b",
            13 => x"04",
            14 => x"84",
            15 => x"0b",
            16 => x"04",
            17 => x"84",
            18 => x"0b",
            19 => x"04",
            20 => x"84",
            21 => x"0b",
            22 => x"04",
            23 => x"85",
            24 => x"0b",
            25 => x"04",
            26 => x"85",
            27 => x"0b",
            28 => x"04",
            29 => x"85",
            30 => x"0b",
            31 => x"04",
            32 => x"85",
            33 => x"0b",
            34 => x"04",
            35 => x"86",
            36 => x"0b",
            37 => x"04",
            38 => x"86",
            39 => x"0b",
            40 => x"04",
            41 => x"86",
            42 => x"0b",
            43 => x"04",
            44 => x"86",
            45 => x"0b",
            46 => x"04",
            47 => x"87",
            48 => x"0b",
            49 => x"04",
            50 => x"87",
            51 => x"0b",
            52 => x"04",
            53 => x"87",
            54 => x"0b",
            55 => x"04",
            56 => x"87",
            57 => x"0b",
            58 => x"04",
            59 => x"88",
            60 => x"0b",
            61 => x"04",
            62 => x"88",
            63 => x"0b",
            64 => x"04",
            65 => x"88",
            66 => x"0b",
            67 => x"04",
            68 => x"88",
            69 => x"0b",
            70 => x"04",
            71 => x"89",
            72 => x"0b",
            73 => x"04",
            74 => x"89",
            75 => x"0b",
            76 => x"04",
            77 => x"89",
            78 => x"0b",
            79 => x"04",
            80 => x"89",
            81 => x"0b",
            82 => x"04",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"80",
           129 => x"d4",
           130 => x"80",
           131 => x"d4",
           132 => x"90",
           133 => x"d4",
           134 => x"c0",
           135 => x"d4",
           136 => x"90",
           137 => x"d4",
           138 => x"85",
           139 => x"d4",
           140 => x"90",
           141 => x"d4",
           142 => x"a3",
           143 => x"d4",
           144 => x"90",
           145 => x"d4",
           146 => x"f7",
           147 => x"d4",
           148 => x"90",
           149 => x"d4",
           150 => x"8b",
           151 => x"d4",
           152 => x"90",
           153 => x"d4",
           154 => x"c4",
           155 => x"d4",
           156 => x"90",
           157 => x"d4",
           158 => x"a8",
           159 => x"d4",
           160 => x"90",
           161 => x"d4",
           162 => x"be",
           163 => x"d4",
           164 => x"90",
           165 => x"d4",
           166 => x"9d",
           167 => x"d4",
           168 => x"90",
           169 => x"d4",
           170 => x"b3",
           171 => x"d4",
           172 => x"90",
           173 => x"d4",
           174 => x"d7",
           175 => x"d4",
           176 => x"90",
           177 => x"d4",
           178 => x"80",
           179 => x"d4",
           180 => x"90",
           181 => x"d4",
           182 => x"ce",
           183 => x"d4",
           184 => x"90",
           185 => x"d4",
           186 => x"d8",
           187 => x"d4",
           188 => x"90",
           189 => x"d4",
           190 => x"90",
           191 => x"d4",
           192 => x"90",
           193 => x"d4",
           194 => x"ea",
           195 => x"d4",
           196 => x"90",
           197 => x"d4",
           198 => x"f2",
           199 => x"d4",
           200 => x"90",
           201 => x"d4",
           202 => x"e9",
           203 => x"d4",
           204 => x"90",
           205 => x"d4",
           206 => x"f8",
           207 => x"d4",
           208 => x"90",
           209 => x"d4",
           210 => x"df",
           211 => x"d4",
           212 => x"90",
           213 => x"d4",
           214 => x"92",
           215 => x"d4",
           216 => x"90",
           217 => x"d4",
           218 => x"86",
           219 => x"d4",
           220 => x"90",
           221 => x"d4",
           222 => x"9a",
           223 => x"d4",
           224 => x"90",
           225 => x"d4",
           226 => x"bd",
           227 => x"d4",
           228 => x"90",
           229 => x"d4",
           230 => x"e1",
           231 => x"d4",
           232 => x"90",
           233 => x"d4",
           234 => x"8a",
           235 => x"d4",
           236 => x"90",
           237 => x"d4",
           238 => x"9a",
           239 => x"d4",
           240 => x"90",
           241 => x"d4",
           242 => x"92",
           243 => x"d4",
           244 => x"90",
           245 => x"d4",
           246 => x"f3",
           247 => x"d4",
           248 => x"90",
           249 => x"d4",
           250 => x"80",
           251 => x"d4",
           252 => x"90",
           253 => x"d4",
           254 => x"f7",
           255 => x"d4",
           256 => x"90",
           257 => x"d4",
           258 => x"fd",
           259 => x"d4",
           260 => x"90",
           261 => x"d4",
           262 => x"c9",
           263 => x"d4",
           264 => x"90",
           265 => x"d4",
           266 => x"a2",
           267 => x"d4",
           268 => x"90",
           269 => x"d4",
           270 => x"cc",
           271 => x"d4",
           272 => x"90",
           273 => x"d4",
           274 => x"da",
           275 => x"d4",
           276 => x"90",
           277 => x"d4",
           278 => x"f6",
           279 => x"d4",
           280 => x"90",
           281 => x"d4",
           282 => x"81",
           283 => x"d4",
           284 => x"90",
           285 => x"d4",
           286 => x"ee",
           287 => x"d4",
           288 => x"90",
           289 => x"d4",
           290 => x"83",
           291 => x"d4",
           292 => x"90",
           293 => x"d4",
           294 => x"df",
           295 => x"d4",
           296 => x"90",
           297 => x"d4",
           298 => x"fe",
           299 => x"d4",
           300 => x"90",
           301 => x"d4",
           302 => x"d7",
           303 => x"d4",
           304 => x"90",
           305 => x"d4",
           306 => x"b1",
           307 => x"d4",
           308 => x"90",
           309 => x"d4",
           310 => x"81",
           311 => x"d4",
           312 => x"90",
           313 => x"d4",
           314 => x"e6",
           315 => x"d4",
           316 => x"90",
           317 => x"d4",
           318 => x"f3",
           319 => x"d4",
           320 => x"90",
           321 => x"d4",
           322 => x"dd",
           323 => x"d4",
           324 => x"90",
           325 => x"c8",
           326 => x"cc",
           327 => x"80",
           328 => x"05",
           329 => x"0b",
           330 => x"04",
           331 => x"51",
           332 => x"04",
           333 => x"d3",
           334 => x"91",
           335 => x"fd",
           336 => x"53",
           337 => x"08",
           338 => x"52",
           339 => x"08",
           340 => x"51",
           341 => x"91",
           342 => x"70",
           343 => x"0c",
           344 => x"0d",
           345 => x"0c",
           346 => x"d4",
           347 => x"d3",
           348 => x"3d",
           349 => x"91",
           350 => x"8c",
           351 => x"91",
           352 => x"88",
           353 => x"93",
           354 => x"c8",
           355 => x"d3",
           356 => x"85",
           357 => x"d3",
           358 => x"91",
           359 => x"02",
           360 => x"0c",
           361 => x"81",
           362 => x"d4",
           363 => x"0c",
           364 => x"d3",
           365 => x"05",
           366 => x"d4",
           367 => x"08",
           368 => x"08",
           369 => x"27",
           370 => x"d3",
           371 => x"05",
           372 => x"ae",
           373 => x"91",
           374 => x"8c",
           375 => x"a2",
           376 => x"d4",
           377 => x"08",
           378 => x"d4",
           379 => x"0c",
           380 => x"08",
           381 => x"10",
           382 => x"08",
           383 => x"ff",
           384 => x"d3",
           385 => x"05",
           386 => x"80",
           387 => x"d3",
           388 => x"05",
           389 => x"d4",
           390 => x"08",
           391 => x"91",
           392 => x"88",
           393 => x"d3",
           394 => x"05",
           395 => x"d3",
           396 => x"05",
           397 => x"d4",
           398 => x"08",
           399 => x"08",
           400 => x"07",
           401 => x"08",
           402 => x"91",
           403 => x"fc",
           404 => x"2a",
           405 => x"08",
           406 => x"91",
           407 => x"8c",
           408 => x"2a",
           409 => x"08",
           410 => x"ff",
           411 => x"d3",
           412 => x"05",
           413 => x"93",
           414 => x"d4",
           415 => x"08",
           416 => x"d4",
           417 => x"0c",
           418 => x"91",
           419 => x"f8",
           420 => x"91",
           421 => x"f4",
           422 => x"91",
           423 => x"f4",
           424 => x"d3",
           425 => x"3d",
           426 => x"d4",
           427 => x"3d",
           428 => x"71",
           429 => x"9f",
           430 => x"55",
           431 => x"72",
           432 => x"74",
           433 => x"70",
           434 => x"38",
           435 => x"71",
           436 => x"38",
           437 => x"81",
           438 => x"ff",
           439 => x"ff",
           440 => x"06",
           441 => x"91",
           442 => x"86",
           443 => x"74",
           444 => x"75",
           445 => x"90",
           446 => x"54",
           447 => x"27",
           448 => x"71",
           449 => x"53",
           450 => x"70",
           451 => x"0c",
           452 => x"84",
           453 => x"72",
           454 => x"05",
           455 => x"12",
           456 => x"26",
           457 => x"72",
           458 => x"72",
           459 => x"05",
           460 => x"12",
           461 => x"26",
           462 => x"53",
           463 => x"fb",
           464 => x"79",
           465 => x"83",
           466 => x"52",
           467 => x"71",
           468 => x"54",
           469 => x"73",
           470 => x"c6",
           471 => x"54",
           472 => x"70",
           473 => x"52",
           474 => x"2e",
           475 => x"33",
           476 => x"2e",
           477 => x"95",
           478 => x"81",
           479 => x"70",
           480 => x"54",
           481 => x"70",
           482 => x"33",
           483 => x"ff",
           484 => x"ff",
           485 => x"31",
           486 => x"0c",
           487 => x"3d",
           488 => x"09",
           489 => x"fd",
           490 => x"70",
           491 => x"81",
           492 => x"51",
           493 => x"38",
           494 => x"16",
           495 => x"56",
           496 => x"08",
           497 => x"73",
           498 => x"ff",
           499 => x"0b",
           500 => x"0c",
           501 => x"04",
           502 => x"80",
           503 => x"71",
           504 => x"87",
           505 => x"d3",
           506 => x"ff",
           507 => x"81",
           508 => x"83",
           509 => x"38",
           510 => x"c8",
           511 => x"0d",
           512 => x"0d",
           513 => x"70",
           514 => x"73",
           515 => x"cd",
           516 => x"51",
           517 => x"09",
           518 => x"38",
           519 => x"33",
           520 => x"a0",
           521 => x"73",
           522 => x"81",
           523 => x"72",
           524 => x"70",
           525 => x"38",
           526 => x"30",
           527 => x"74",
           528 => x"70",
           529 => x"33",
           530 => x"2e",
           531 => x"88",
           532 => x"70",
           533 => x"34",
           534 => x"73",
           535 => x"d3",
           536 => x"3d",
           537 => x"3d",
           538 => x"72",
           539 => x"91",
           540 => x"fc",
           541 => x"51",
           542 => x"91",
           543 => x"85",
           544 => x"83",
           545 => x"72",
           546 => x"0c",
           547 => x"04",
           548 => x"7d",
           549 => x"ff",
           550 => x"81",
           551 => x"26",
           552 => x"83",
           553 => x"05",
           554 => x"79",
           555 => x"b1",
           556 => x"33",
           557 => x"79",
           558 => x"a5",
           559 => x"33",
           560 => x"79",
           561 => x"99",
           562 => x"33",
           563 => x"79",
           564 => x"8d",
           565 => x"22",
           566 => x"79",
           567 => x"81",
           568 => x"1c",
           569 => x"5b",
           570 => x"26",
           571 => x"8a",
           572 => x"88",
           573 => x"86",
           574 => x"85",
           575 => x"84",
           576 => x"83",
           577 => x"82",
           578 => x"7b",
           579 => x"b6",
           580 => x"89",
           581 => x"98",
           582 => x"7b",
           583 => x"87",
           584 => x"0c",
           585 => x"87",
           586 => x"0c",
           587 => x"87",
           588 => x"0c",
           589 => x"87",
           590 => x"0c",
           591 => x"87",
           592 => x"0c",
           593 => x"87",
           594 => x"0c",
           595 => x"87",
           596 => x"0c",
           597 => x"87",
           598 => x"0c",
           599 => x"80",
           600 => x"d3",
           601 => x"3d",
           602 => x"3d",
           603 => x"87",
           604 => x"5c",
           605 => x"87",
           606 => x"08",
           607 => x"23",
           608 => x"b8",
           609 => x"82",
           610 => x"c0",
           611 => x"5b",
           612 => x"34",
           613 => x"b0",
           614 => x"84",
           615 => x"c0",
           616 => x"5b",
           617 => x"34",
           618 => x"a8",
           619 => x"86",
           620 => x"c0",
           621 => x"5b",
           622 => x"23",
           623 => x"a0",
           624 => x"8a",
           625 => x"7c",
           626 => x"22",
           627 => x"22",
           628 => x"33",
           629 => x"33",
           630 => x"33",
           631 => x"33",
           632 => x"33",
           633 => x"52",
           634 => x"51",
           635 => x"8d",
           636 => x"80",
           637 => x"8b",
           638 => x"30",
           639 => x"51",
           640 => x"0b",
           641 => x"c0",
           642 => x"0d",
           643 => x"0d",
           644 => x"91",
           645 => x"54",
           646 => x"94",
           647 => x"80",
           648 => x"87",
           649 => x"51",
           650 => x"96",
           651 => x"06",
           652 => x"70",
           653 => x"38",
           654 => x"70",
           655 => x"51",
           656 => x"71",
           657 => x"32",
           658 => x"51",
           659 => x"2e",
           660 => x"93",
           661 => x"06",
           662 => x"ff",
           663 => x"0b",
           664 => x"33",
           665 => x"94",
           666 => x"80",
           667 => x"87",
           668 => x"52",
           669 => x"73",
           670 => x"0c",
           671 => x"04",
           672 => x"02",
           673 => x"0b",
           674 => x"c0",
           675 => x"87",
           676 => x"51",
           677 => x"86",
           678 => x"94",
           679 => x"08",
           680 => x"70",
           681 => x"52",
           682 => x"2e",
           683 => x"91",
           684 => x"06",
           685 => x"d7",
           686 => x"2a",
           687 => x"81",
           688 => x"70",
           689 => x"38",
           690 => x"70",
           691 => x"51",
           692 => x"38",
           693 => x"cb",
           694 => x"87",
           695 => x"52",
           696 => x"86",
           697 => x"94",
           698 => x"72",
           699 => x"0d",
           700 => x"0d",
           701 => x"74",
           702 => x"70",
           703 => x"f7",
           704 => x"81",
           705 => x"0b",
           706 => x"c0",
           707 => x"87",
           708 => x"51",
           709 => x"86",
           710 => x"94",
           711 => x"08",
           712 => x"70",
           713 => x"52",
           714 => x"2e",
           715 => x"91",
           716 => x"06",
           717 => x"d7",
           718 => x"2a",
           719 => x"81",
           720 => x"70",
           721 => x"38",
           722 => x"70",
           723 => x"51",
           724 => x"38",
           725 => x"cb",
           726 => x"87",
           727 => x"52",
           728 => x"86",
           729 => x"94",
           730 => x"72",
           731 => x"74",
           732 => x"70",
           733 => x"75",
           734 => x"0c",
           735 => x"04",
           736 => x"0b",
           737 => x"c0",
           738 => x"c0",
           739 => x"71",
           740 => x"38",
           741 => x"94",
           742 => x"70",
           743 => x"81",
           744 => x"51",
           745 => x"e2",
           746 => x"91",
           747 => x"51",
           748 => x"80",
           749 => x"2e",
           750 => x"c0",
           751 => x"71",
           752 => x"ff",
           753 => x"c8",
           754 => x"3d",
           755 => x"3d",
           756 => x"91",
           757 => x"51",
           758 => x"84",
           759 => x"2e",
           760 => x"c0",
           761 => x"71",
           762 => x"2a",
           763 => x"51",
           764 => x"52",
           765 => x"a2",
           766 => x"91",
           767 => x"51",
           768 => x"80",
           769 => x"2e",
           770 => x"c0",
           771 => x"71",
           772 => x"2b",
           773 => x"51",
           774 => x"91",
           775 => x"83",
           776 => x"fd",
           777 => x"c0",
           778 => x"08",
           779 => x"8a",
           780 => x"53",
           781 => x"83",
           782 => x"cb",
           783 => x"c0",
           784 => x"71",
           785 => x"87",
           786 => x"08",
           787 => x"88",
           788 => x"9e",
           789 => x"0c",
           790 => x"87",
           791 => x"08",
           792 => x"90",
           793 => x"9e",
           794 => x"0c",
           795 => x"87",
           796 => x"08",
           797 => x"98",
           798 => x"9e",
           799 => x"0c",
           800 => x"87",
           801 => x"08",
           802 => x"a0",
           803 => x"9e",
           804 => x"0c",
           805 => x"52",
           806 => x"13",
           807 => x"87",
           808 => x"08",
           809 => x"81",
           810 => x"34",
           811 => x"80",
           812 => x"9e",
           813 => x"a0",
           814 => x"52",
           815 => x"2e",
           816 => x"53",
           817 => x"80",
           818 => x"9e",
           819 => x"81",
           820 => x"51",
           821 => x"80",
           822 => x"81",
           823 => x"cb",
           824 => x"0b",
           825 => x"88",
           826 => x"c0",
           827 => x"52",
           828 => x"2e",
           829 => x"52",
           830 => x"f3",
           831 => x"87",
           832 => x"08",
           833 => x"06",
           834 => x"70",
           835 => x"38",
           836 => x"91",
           837 => x"80",
           838 => x"9e",
           839 => x"88",
           840 => x"52",
           841 => x"2e",
           842 => x"52",
           843 => x"f5",
           844 => x"87",
           845 => x"08",
           846 => x"06",
           847 => x"70",
           848 => x"38",
           849 => x"91",
           850 => x"80",
           851 => x"9e",
           852 => x"82",
           853 => x"52",
           854 => x"2e",
           855 => x"52",
           856 => x"f7",
           857 => x"87",
           858 => x"08",
           859 => x"06",
           860 => x"70",
           861 => x"38",
           862 => x"91",
           863 => x"91",
           864 => x"87",
           865 => x"70",
           866 => x"e0",
           867 => x"2c",
           868 => x"53",
           869 => x"81",
           870 => x"71",
           871 => x"08",
           872 => x"51",
           873 => x"80",
           874 => x"81",
           875 => x"34",
           876 => x"c0",
           877 => x"70",
           878 => x"52",
           879 => x"2e",
           880 => x"52",
           881 => x"fb",
           882 => x"9e",
           883 => x"87",
           884 => x"70",
           885 => x"34",
           886 => x"04",
           887 => x"91",
           888 => x"84",
           889 => x"cb",
           890 => x"73",
           891 => x"38",
           892 => x"51",
           893 => x"91",
           894 => x"84",
           895 => x"cb",
           896 => x"55",
           897 => x"2e",
           898 => x"15",
           899 => x"cb",
           900 => x"91",
           901 => x"8a",
           902 => x"cb",
           903 => x"55",
           904 => x"2e",
           905 => x"15",
           906 => x"15",
           907 => x"b7",
           908 => x"e9",
           909 => x"f3",
           910 => x"55",
           911 => x"81",
           912 => x"73",
           913 => x"38",
           914 => x"70",
           915 => x"11",
           916 => x"91",
           917 => x"89",
           918 => x"cb",
           919 => x"73",
           920 => x"38",
           921 => x"51",
           922 => x"91",
           923 => x"54",
           924 => x"88",
           925 => x"fc",
           926 => x"3f",
           927 => x"33",
           928 => x"2e",
           929 => x"b8",
           930 => x"97",
           931 => x"f8",
           932 => x"55",
           933 => x"8c",
           934 => x"33",
           935 => x"94",
           936 => x"3f",
           937 => x"33",
           938 => x"2e",
           939 => x"b8",
           940 => x"ef",
           941 => x"fb",
           942 => x"55",
           943 => x"8c",
           944 => x"33",
           945 => x"d0",
           946 => x"3f",
           947 => x"51",
           948 => x"91",
           949 => x"70",
           950 => x"52",
           951 => x"b8",
           952 => x"55",
           953 => x"73",
           954 => x"b9",
           955 => x"ad",
           956 => x"08",
           957 => x"c8",
           958 => x"3f",
           959 => x"52",
           960 => x"51",
           961 => x"90",
           962 => x"91",
           963 => x"88",
           964 => x"3d",
           965 => x"3d",
           966 => x"05",
           967 => x"85",
           968 => x"71",
           969 => x"0b",
           970 => x"05",
           971 => x"04",
           972 => x"51",
           973 => x"ac",
           974 => x"c8",
           975 => x"3f",
           976 => x"ba",
           977 => x"a9",
           978 => x"91",
           979 => x"f7",
           980 => x"39",
           981 => x"51",
           982 => x"88",
           983 => x"e4",
           984 => x"3f",
           985 => x"04",
           986 => x"0c",
           987 => x"87",
           988 => x"0c",
           989 => x"0d",
           990 => x"84",
           991 => x"52",
           992 => x"70",
           993 => x"91",
           994 => x"72",
           995 => x"0d",
           996 => x"0d",
           997 => x"84",
           998 => x"cc",
           999 => x"80",
          1000 => x"09",
          1001 => x"80",
          1002 => x"91",
          1003 => x"73",
          1004 => x"3d",
          1005 => x"cc",
          1006 => x"c0",
          1007 => x"04",
          1008 => x"02",
          1009 => x"53",
          1010 => x"09",
          1011 => x"38",
          1012 => x"3f",
          1013 => x"08",
          1014 => x"38",
          1015 => x"08",
          1016 => x"34",
          1017 => x"08",
          1018 => x"d3",
          1019 => x"39",
          1020 => x"08",
          1021 => x"38",
          1022 => x"d3",
          1023 => x"71",
          1024 => x"0d",
          1025 => x"0d",
          1026 => x"33",
          1027 => x"08",
          1028 => x"d8",
          1029 => x"ff",
          1030 => x"91",
          1031 => x"84",
          1032 => x"fe",
          1033 => x"70",
          1034 => x"71",
          1035 => x"38",
          1036 => x"05",
          1037 => x"ff",
          1038 => x"33",
          1039 => x"38",
          1040 => x"04",
          1041 => x"76",
          1042 => x"08",
          1043 => x"d8",
          1044 => x"54",
          1045 => x"80",
          1046 => x"72",
          1047 => x"54",
          1048 => x"dc",
          1049 => x"52",
          1050 => x"73",
          1051 => x"0c",
          1052 => x"04",
          1053 => x"66",
          1054 => x"78",
          1055 => x"5a",
          1056 => x"80",
          1057 => x"38",
          1058 => x"88",
          1059 => x"fe",
          1060 => x"39",
          1061 => x"70",
          1062 => x"33",
          1063 => x"75",
          1064 => x"81",
          1065 => x"81",
          1066 => x"05",
          1067 => x"5d",
          1068 => x"ad",
          1069 => x"06",
          1070 => x"79",
          1071 => x"5b",
          1072 => x"75",
          1073 => x"81",
          1074 => x"7b",
          1075 => x"08",
          1076 => x"05",
          1077 => x"5c",
          1078 => x"39",
          1079 => x"72",
          1080 => x"38",
          1081 => x"16",
          1082 => x"70",
          1083 => x"33",
          1084 => x"57",
          1085 => x"27",
          1086 => x"80",
          1087 => x"30",
          1088 => x"80",
          1089 => x"cc",
          1090 => x"70",
          1091 => x"25",
          1092 => x"59",
          1093 => x"54",
          1094 => x"8c",
          1095 => x"07",
          1096 => x"05",
          1097 => x"5d",
          1098 => x"83",
          1099 => x"55",
          1100 => x"27",
          1101 => x"16",
          1102 => x"06",
          1103 => x"be",
          1104 => x"96",
          1105 => x"38",
          1106 => x"91",
          1107 => x"53",
          1108 => x"7b",
          1109 => x"08",
          1110 => x"80",
          1111 => x"54",
          1112 => x"8d",
          1113 => x"70",
          1114 => x"51",
          1115 => x"f5",
          1116 => x"2a",
          1117 => x"51",
          1118 => x"38",
          1119 => x"55",
          1120 => x"27",
          1121 => x"81",
          1122 => x"56",
          1123 => x"b0",
          1124 => x"38",
          1125 => x"55",
          1126 => x"26",
          1127 => x"51",
          1128 => x"73",
          1129 => x"53",
          1130 => x"fd",
          1131 => x"51",
          1132 => x"73",
          1133 => x"53",
          1134 => x"f2",
          1135 => x"39",
          1136 => x"83",
          1137 => x"5d",
          1138 => x"3f",
          1139 => x"82",
          1140 => x"88",
          1141 => x"8a",
          1142 => x"90",
          1143 => x"75",
          1144 => x"3f",
          1145 => x"7c",
          1146 => x"81",
          1147 => x"72",
          1148 => x"38",
          1149 => x"71",
          1150 => x"53",
          1151 => x"80",
          1152 => x"81",
          1153 => x"7b",
          1154 => x"08",
          1155 => x"89",
          1156 => x"1d",
          1157 => x"5d",
          1158 => x"c4",
          1159 => x"70",
          1160 => x"25",
          1161 => x"24",
          1162 => x"55",
          1163 => x"2e",
          1164 => x"30",
          1165 => x"5e",
          1166 => x"7a",
          1167 => x"e6",
          1168 => x"d3",
          1169 => x"ff",
          1170 => x"77",
          1171 => x"e6",
          1172 => x"c8",
          1173 => x"75",
          1174 => x"74",
          1175 => x"81",
          1176 => x"54",
          1177 => x"f8",
          1178 => x"87",
          1179 => x"ff",
          1180 => x"96",
          1181 => x"e0",
          1182 => x"54",
          1183 => x"34",
          1184 => x"30",
          1185 => x"9f",
          1186 => x"74",
          1187 => x"51",
          1188 => x"ff",
          1189 => x"84",
          1190 => x"06",
          1191 => x"80",
          1192 => x"96",
          1193 => x"e0",
          1194 => x"73",
          1195 => x"58",
          1196 => x"06",
          1197 => x"55",
          1198 => x"a0",
          1199 => x"2a",
          1200 => x"51",
          1201 => x"38",
          1202 => x"55",
          1203 => x"27",
          1204 => x"81",
          1205 => x"56",
          1206 => x"e4",
          1207 => x"38",
          1208 => x"55",
          1209 => x"26",
          1210 => x"18",
          1211 => x"05",
          1212 => x"53",
          1213 => x"c8",
          1214 => x"38",
          1215 => x"55",
          1216 => x"27",
          1217 => x"a0",
          1218 => x"3f",
          1219 => x"55",
          1220 => x"26",
          1221 => x"e3",
          1222 => x"0d",
          1223 => x"0d",
          1224 => x"70",
          1225 => x"08",
          1226 => x"51",
          1227 => x"85",
          1228 => x"fe",
          1229 => x"91",
          1230 => x"85",
          1231 => x"52",
          1232 => x"b0",
          1233 => x"e0",
          1234 => x"73",
          1235 => x"91",
          1236 => x"84",
          1237 => x"fd",
          1238 => x"d3",
          1239 => x"91",
          1240 => x"87",
          1241 => x"53",
          1242 => x"fa",
          1243 => x"91",
          1244 => x"85",
          1245 => x"fa",
          1246 => x"7a",
          1247 => x"53",
          1248 => x"08",
          1249 => x"fa",
          1250 => x"73",
          1251 => x"39",
          1252 => x"d3",
          1253 => x"71",
          1254 => x"c8",
          1255 => x"06",
          1256 => x"2e",
          1257 => x"8d",
          1258 => x"38",
          1259 => x"70",
          1260 => x"70",
          1261 => x"2a",
          1262 => x"06",
          1263 => x"53",
          1264 => x"8e",
          1265 => x"74",
          1266 => x"52",
          1267 => x"3f",
          1268 => x"74",
          1269 => x"38",
          1270 => x"74",
          1271 => x"b2",
          1272 => x"52",
          1273 => x"81",
          1274 => x"ff",
          1275 => x"f7",
          1276 => x"9e",
          1277 => x"52",
          1278 => x"8a",
          1279 => x"3f",
          1280 => x"91",
          1281 => x"88",
          1282 => x"fe",
          1283 => x"d3",
          1284 => x"91",
          1285 => x"77",
          1286 => x"53",
          1287 => x"72",
          1288 => x"0c",
          1289 => x"04",
          1290 => x"7a",
          1291 => x"80",
          1292 => x"75",
          1293 => x"56",
          1294 => x"a0",
          1295 => x"06",
          1296 => x"08",
          1297 => x"0c",
          1298 => x"33",
          1299 => x"a0",
          1300 => x"73",
          1301 => x"81",
          1302 => x"81",
          1303 => x"76",
          1304 => x"70",
          1305 => x"58",
          1306 => x"09",
          1307 => x"d3",
          1308 => x"81",
          1309 => x"74",
          1310 => x"55",
          1311 => x"e2",
          1312 => x"73",
          1313 => x"09",
          1314 => x"38",
          1315 => x"14",
          1316 => x"08",
          1317 => x"54",
          1318 => x"39",
          1319 => x"81",
          1320 => x"75",
          1321 => x"56",
          1322 => x"39",
          1323 => x"74",
          1324 => x"38",
          1325 => x"80",
          1326 => x"89",
          1327 => x"38",
          1328 => x"d0",
          1329 => x"56",
          1330 => x"80",
          1331 => x"39",
          1332 => x"e1",
          1333 => x"80",
          1334 => x"57",
          1335 => x"74",
          1336 => x"38",
          1337 => x"27",
          1338 => x"14",
          1339 => x"06",
          1340 => x"14",
          1341 => x"06",
          1342 => x"74",
          1343 => x"f9",
          1344 => x"ff",
          1345 => x"89",
          1346 => x"38",
          1347 => x"c5",
          1348 => x"29",
          1349 => x"81",
          1350 => x"75",
          1351 => x"56",
          1352 => x"a0",
          1353 => x"38",
          1354 => x"84",
          1355 => x"56",
          1356 => x"81",
          1357 => x"d3",
          1358 => x"3d",
          1359 => x"3d",
          1360 => x"5a",
          1361 => x"7a",
          1362 => x"70",
          1363 => x"58",
          1364 => x"09",
          1365 => x"38",
          1366 => x"05",
          1367 => x"08",
          1368 => x"53",
          1369 => x"f0",
          1370 => x"2e",
          1371 => x"8e",
          1372 => x"08",
          1373 => x"75",
          1374 => x"56",
          1375 => x"b0",
          1376 => x"06",
          1377 => x"74",
          1378 => x"75",
          1379 => x"70",
          1380 => x"73",
          1381 => x"9a",
          1382 => x"f8",
          1383 => x"06",
          1384 => x"0b",
          1385 => x"0c",
          1386 => x"33",
          1387 => x"80",
          1388 => x"75",
          1389 => x"76",
          1390 => x"70",
          1391 => x"57",
          1392 => x"56",
          1393 => x"81",
          1394 => x"14",
          1395 => x"88",
          1396 => x"27",
          1397 => x"f3",
          1398 => x"53",
          1399 => x"89",
          1400 => x"38",
          1401 => x"56",
          1402 => x"80",
          1403 => x"39",
          1404 => x"56",
          1405 => x"80",
          1406 => x"e0",
          1407 => x"38",
          1408 => x"81",
          1409 => x"53",
          1410 => x"81",
          1411 => x"53",
          1412 => x"8e",
          1413 => x"70",
          1414 => x"55",
          1415 => x"27",
          1416 => x"77",
          1417 => x"76",
          1418 => x"75",
          1419 => x"76",
          1420 => x"70",
          1421 => x"56",
          1422 => x"ff",
          1423 => x"80",
          1424 => x"75",
          1425 => x"79",
          1426 => x"75",
          1427 => x"0c",
          1428 => x"04",
          1429 => x"02",
          1430 => x"51",
          1431 => x"72",
          1432 => x"91",
          1433 => x"33",
          1434 => x"d3",
          1435 => x"3d",
          1436 => x"3d",
          1437 => x"05",
          1438 => x"05",
          1439 => x"55",
          1440 => x"72",
          1441 => x"ed",
          1442 => x"29",
          1443 => x"8c",
          1444 => x"52",
          1445 => x"84",
          1446 => x"52",
          1447 => x"72",
          1448 => x"c0",
          1449 => x"51",
          1450 => x"85",
          1451 => x"98",
          1452 => x"52",
          1453 => x"8c",
          1454 => x"70",
          1455 => x"51",
          1456 => x"87",
          1457 => x"51",
          1458 => x"72",
          1459 => x"c0",
          1460 => x"70",
          1461 => x"80",
          1462 => x"71",
          1463 => x"c0",
          1464 => x"51",
          1465 => x"87",
          1466 => x"cc",
          1467 => x"91",
          1468 => x"33",
          1469 => x"d3",
          1470 => x"3d",
          1471 => x"3d",
          1472 => x"65",
          1473 => x"80",
          1474 => x"56",
          1475 => x"83",
          1476 => x"fe",
          1477 => x"d3",
          1478 => x"06",
          1479 => x"71",
          1480 => x"80",
          1481 => x"87",
          1482 => x"73",
          1483 => x"c0",
          1484 => x"87",
          1485 => x"12",
          1486 => x"57",
          1487 => x"76",
          1488 => x"92",
          1489 => x"71",
          1490 => x"75",
          1491 => x"70",
          1492 => x"81",
          1493 => x"54",
          1494 => x"8e",
          1495 => x"52",
          1496 => x"81",
          1497 => x"81",
          1498 => x"a2",
          1499 => x"80",
          1500 => x"75",
          1501 => x"d5",
          1502 => x"52",
          1503 => x"87",
          1504 => x"80",
          1505 => x"81",
          1506 => x"c0",
          1507 => x"53",
          1508 => x"82",
          1509 => x"71",
          1510 => x"1b",
          1511 => x"84",
          1512 => x"1e",
          1513 => x"06",
          1514 => x"7a",
          1515 => x"38",
          1516 => x"80",
          1517 => x"87",
          1518 => x"26",
          1519 => x"73",
          1520 => x"06",
          1521 => x"2e",
          1522 => x"52",
          1523 => x"91",
          1524 => x"90",
          1525 => x"f3",
          1526 => x"62",
          1527 => x"05",
          1528 => x"56",
          1529 => x"83",
          1530 => x"fc",
          1531 => x"d3",
          1532 => x"06",
          1533 => x"71",
          1534 => x"80",
          1535 => x"98",
          1536 => x"2b",
          1537 => x"8c",
          1538 => x"92",
          1539 => x"41",
          1540 => x"56",
          1541 => x"87",
          1542 => x"19",
          1543 => x"52",
          1544 => x"80",
          1545 => x"70",
          1546 => x"81",
          1547 => x"54",
          1548 => x"8c",
          1549 => x"81",
          1550 => x"78",
          1551 => x"53",
          1552 => x"70",
          1553 => x"52",
          1554 => x"87",
          1555 => x"52",
          1556 => x"75",
          1557 => x"80",
          1558 => x"72",
          1559 => x"99",
          1560 => x"0c",
          1561 => x"8c",
          1562 => x"08",
          1563 => x"51",
          1564 => x"38",
          1565 => x"8d",
          1566 => x"70",
          1567 => x"84",
          1568 => x"5d",
          1569 => x"2e",
          1570 => x"fc",
          1571 => x"52",
          1572 => x"7d",
          1573 => x"fc",
          1574 => x"80",
          1575 => x"71",
          1576 => x"38",
          1577 => x"54",
          1578 => x"c8",
          1579 => x"0d",
          1580 => x"0d",
          1581 => x"05",
          1582 => x"02",
          1583 => x"05",
          1584 => x"55",
          1585 => x"8c",
          1586 => x"c8",
          1587 => x"52",
          1588 => x"bc",
          1589 => x"72",
          1590 => x"38",
          1591 => x"88",
          1592 => x"2e",
          1593 => x"39",
          1594 => x"9a",
          1595 => x"74",
          1596 => x"c0",
          1597 => x"70",
          1598 => x"94",
          1599 => x"0a",
          1600 => x"54",
          1601 => x"80",
          1602 => x"54",
          1603 => x"54",
          1604 => x"c8",
          1605 => x"0d",
          1606 => x"0d",
          1607 => x"81",
          1608 => x"88",
          1609 => x"91",
          1610 => x"52",
          1611 => x"3d",
          1612 => x"3d",
          1613 => x"11",
          1614 => x"33",
          1615 => x"71",
          1616 => x"81",
          1617 => x"07",
          1618 => x"88",
          1619 => x"d3",
          1620 => x"54",
          1621 => x"85",
          1622 => x"ff",
          1623 => x"02",
          1624 => x"05",
          1625 => x"70",
          1626 => x"05",
          1627 => x"88",
          1628 => x"72",
          1629 => x"0d",
          1630 => x"0d",
          1631 => x"52",
          1632 => x"81",
          1633 => x"70",
          1634 => x"70",
          1635 => x"05",
          1636 => x"88",
          1637 => x"72",
          1638 => x"54",
          1639 => x"2a",
          1640 => x"34",
          1641 => x"04",
          1642 => x"76",
          1643 => x"54",
          1644 => x"2e",
          1645 => x"70",
          1646 => x"33",
          1647 => x"05",
          1648 => x"11",
          1649 => x"38",
          1650 => x"04",
          1651 => x"75",
          1652 => x"52",
          1653 => x"70",
          1654 => x"34",
          1655 => x"70",
          1656 => x"3d",
          1657 => x"3d",
          1658 => x"79",
          1659 => x"74",
          1660 => x"56",
          1661 => x"81",
          1662 => x"71",
          1663 => x"16",
          1664 => x"52",
          1665 => x"86",
          1666 => x"2e",
          1667 => x"91",
          1668 => x"86",
          1669 => x"fe",
          1670 => x"76",
          1671 => x"54",
          1672 => x"2e",
          1673 => x"73",
          1674 => x"81",
          1675 => x"52",
          1676 => x"2e",
          1677 => x"73",
          1678 => x"06",
          1679 => x"33",
          1680 => x"0c",
          1681 => x"04",
          1682 => x"d3",
          1683 => x"80",
          1684 => x"c8",
          1685 => x"3d",
          1686 => x"80",
          1687 => x"33",
          1688 => x"78",
          1689 => x"38",
          1690 => x"16",
          1691 => x"16",
          1692 => x"17",
          1693 => x"fa",
          1694 => x"d3",
          1695 => x"2e",
          1696 => x"b8",
          1697 => x"c8",
          1698 => x"34",
          1699 => x"a4",
          1700 => x"55",
          1701 => x"08",
          1702 => x"82",
          1703 => x"74",
          1704 => x"81",
          1705 => x"81",
          1706 => x"08",
          1707 => x"05",
          1708 => x"81",
          1709 => x"fa",
          1710 => x"39",
          1711 => x"91",
          1712 => x"89",
          1713 => x"fa",
          1714 => x"7a",
          1715 => x"56",
          1716 => x"75",
          1717 => x"76",
          1718 => x"3f",
          1719 => x"08",
          1720 => x"c8",
          1721 => x"81",
          1722 => x"b4",
          1723 => x"17",
          1724 => x"8a",
          1725 => x"c8",
          1726 => x"85",
          1727 => x"81",
          1728 => x"18",
          1729 => x"d3",
          1730 => x"3d",
          1731 => x"3d",
          1732 => x"52",
          1733 => x"3f",
          1734 => x"08",
          1735 => x"c8",
          1736 => x"38",
          1737 => x"74",
          1738 => x"81",
          1739 => x"38",
          1740 => x"59",
          1741 => x"09",
          1742 => x"e3",
          1743 => x"53",
          1744 => x"08",
          1745 => x"70",
          1746 => x"80",
          1747 => x"d5",
          1748 => x"17",
          1749 => x"3f",
          1750 => x"a4",
          1751 => x"51",
          1752 => x"86",
          1753 => x"f2",
          1754 => x"17",
          1755 => x"3f",
          1756 => x"52",
          1757 => x"51",
          1758 => x"8c",
          1759 => x"84",
          1760 => x"fb",
          1761 => x"17",
          1762 => x"70",
          1763 => x"79",
          1764 => x"52",
          1765 => x"51",
          1766 => x"77",
          1767 => x"80",
          1768 => x"81",
          1769 => x"fa",
          1770 => x"d3",
          1771 => x"2e",
          1772 => x"58",
          1773 => x"c8",
          1774 => x"0d",
          1775 => x"0d",
          1776 => x"98",
          1777 => x"05",
          1778 => x"80",
          1779 => x"27",
          1780 => x"14",
          1781 => x"29",
          1782 => x"05",
          1783 => x"91",
          1784 => x"87",
          1785 => x"f9",
          1786 => x"7a",
          1787 => x"54",
          1788 => x"27",
          1789 => x"14",
          1790 => x"86",
          1791 => x"81",
          1792 => x"74",
          1793 => x"72",
          1794 => x"f5",
          1795 => x"24",
          1796 => x"81",
          1797 => x"81",
          1798 => x"83",
          1799 => x"38",
          1800 => x"74",
          1801 => x"70",
          1802 => x"16",
          1803 => x"74",
          1804 => x"93",
          1805 => x"c8",
          1806 => x"38",
          1807 => x"06",
          1808 => x"33",
          1809 => x"89",
          1810 => x"08",
          1811 => x"54",
          1812 => x"fc",
          1813 => x"d3",
          1814 => x"fe",
          1815 => x"ff",
          1816 => x"11",
          1817 => x"2b",
          1818 => x"81",
          1819 => x"2a",
          1820 => x"51",
          1821 => x"e2",
          1822 => x"ff",
          1823 => x"da",
          1824 => x"2a",
          1825 => x"05",
          1826 => x"fc",
          1827 => x"d3",
          1828 => x"c6",
          1829 => x"83",
          1830 => x"05",
          1831 => x"f8",
          1832 => x"d3",
          1833 => x"ff",
          1834 => x"ae",
          1835 => x"2a",
          1836 => x"05",
          1837 => x"fc",
          1838 => x"d3",
          1839 => x"38",
          1840 => x"83",
          1841 => x"05",
          1842 => x"f8",
          1843 => x"d3",
          1844 => x"0a",
          1845 => x"39",
          1846 => x"91",
          1847 => x"89",
          1848 => x"f7",
          1849 => x"7d",
          1850 => x"55",
          1851 => x"74",
          1852 => x"38",
          1853 => x"08",
          1854 => x"38",
          1855 => x"72",
          1856 => x"a8",
          1857 => x"24",
          1858 => x"81",
          1859 => x"82",
          1860 => x"83",
          1861 => x"38",
          1862 => x"73",
          1863 => x"70",
          1864 => x"17",
          1865 => x"75",
          1866 => x"9b",
          1867 => x"c8",
          1868 => x"d3",
          1869 => x"ea",
          1870 => x"ff",
          1871 => x"11",
          1872 => x"81",
          1873 => x"51",
          1874 => x"72",
          1875 => x"38",
          1876 => x"9f",
          1877 => x"33",
          1878 => x"07",
          1879 => x"78",
          1880 => x"83",
          1881 => x"89",
          1882 => x"08",
          1883 => x"51",
          1884 => x"91",
          1885 => x"57",
          1886 => x"08",
          1887 => x"78",
          1888 => x"15",
          1889 => x"81",
          1890 => x"2a",
          1891 => x"58",
          1892 => x"75",
          1893 => x"33",
          1894 => x"76",
          1895 => x"07",
          1896 => x"34",
          1897 => x"16",
          1898 => x"39",
          1899 => x"a4",
          1900 => x"52",
          1901 => x"8f",
          1902 => x"c8",
          1903 => x"d3",
          1904 => x"de",
          1905 => x"ff",
          1906 => x"73",
          1907 => x"06",
          1908 => x"05",
          1909 => x"3f",
          1910 => x"16",
          1911 => x"39",
          1912 => x"a4",
          1913 => x"52",
          1914 => x"db",
          1915 => x"c8",
          1916 => x"d3",
          1917 => x"38",
          1918 => x"06",
          1919 => x"83",
          1920 => x"11",
          1921 => x"54",
          1922 => x"f6",
          1923 => x"d3",
          1924 => x"0a",
          1925 => x"52",
          1926 => x"dd",
          1927 => x"83",
          1928 => x"91",
          1929 => x"8b",
          1930 => x"f9",
          1931 => x"7b",
          1932 => x"58",
          1933 => x"81",
          1934 => x"38",
          1935 => x"74",
          1936 => x"82",
          1937 => x"39",
          1938 => x"aa",
          1939 => x"75",
          1940 => x"fd",
          1941 => x"d3",
          1942 => x"91",
          1943 => x"80",
          1944 => x"39",
          1945 => x"ed",
          1946 => x"80",
          1947 => x"d3",
          1948 => x"80",
          1949 => x"52",
          1950 => x"eb",
          1951 => x"c8",
          1952 => x"d3",
          1953 => x"2e",
          1954 => x"91",
          1955 => x"81",
          1956 => x"91",
          1957 => x"ff",
          1958 => x"80",
          1959 => x"74",
          1960 => x"3f",
          1961 => x"08",
          1962 => x"15",
          1963 => x"54",
          1964 => x"74",
          1965 => x"90",
          1966 => x"05",
          1967 => x"84",
          1968 => x"07",
          1969 => x"16",
          1970 => x"98",
          1971 => x"26",
          1972 => x"80",
          1973 => x"d3",
          1974 => x"3d",
          1975 => x"3d",
          1976 => x"71",
          1977 => x"5c",
          1978 => x"8c",
          1979 => x"77",
          1980 => x"38",
          1981 => x"78",
          1982 => x"81",
          1983 => x"7a",
          1984 => x"f9",
          1985 => x"55",
          1986 => x"c8",
          1987 => x"e9",
          1988 => x"c8",
          1989 => x"d3",
          1990 => x"2e",
          1991 => x"91",
          1992 => x"55",
          1993 => x"91",
          1994 => x"26",
          1995 => x"7a",
          1996 => x"90",
          1997 => x"2e",
          1998 => x"80",
          1999 => x"2e",
          2000 => x"80",
          2001 => x"1b",
          2002 => x"08",
          2003 => x"38",
          2004 => x"52",
          2005 => x"8f",
          2006 => x"c8",
          2007 => x"5a",
          2008 => x"08",
          2009 => x"81",
          2010 => x"91",
          2011 => x"5a",
          2012 => x"70",
          2013 => x"07",
          2014 => x"7d",
          2015 => x"51",
          2016 => x"73",
          2017 => x"75",
          2018 => x"38",
          2019 => x"56",
          2020 => x"8a",
          2021 => x"1a",
          2022 => x"38",
          2023 => x"57",
          2024 => x"38",
          2025 => x"17",
          2026 => x"08",
          2027 => x"38",
          2028 => x"78",
          2029 => x"38",
          2030 => x"51",
          2031 => x"91",
          2032 => x"56",
          2033 => x"08",
          2034 => x"38",
          2035 => x"d3",
          2036 => x"2e",
          2037 => x"86",
          2038 => x"c8",
          2039 => x"ff",
          2040 => x"70",
          2041 => x"25",
          2042 => x"51",
          2043 => x"73",
          2044 => x"76",
          2045 => x"81",
          2046 => x"38",
          2047 => x"f9",
          2048 => x"76",
          2049 => x"f9",
          2050 => x"d3",
          2051 => x"d3",
          2052 => x"70",
          2053 => x"08",
          2054 => x"7d",
          2055 => x"07",
          2056 => x"06",
          2057 => x"56",
          2058 => x"2e",
          2059 => x"53",
          2060 => x"51",
          2061 => x"91",
          2062 => x"56",
          2063 => x"76",
          2064 => x"98",
          2065 => x"05",
          2066 => x"08",
          2067 => x"38",
          2068 => x"ff",
          2069 => x"0c",
          2070 => x"81",
          2071 => x"84",
          2072 => x"39",
          2073 => x"81",
          2074 => x"89",
          2075 => x"89",
          2076 => x"85",
          2077 => x"76",
          2078 => x"d3",
          2079 => x"3d",
          2080 => x"3d",
          2081 => x"52",
          2082 => x"3f",
          2083 => x"d3",
          2084 => x"db",
          2085 => x"76",
          2086 => x"3f",
          2087 => x"08",
          2088 => x"08",
          2089 => x"5a",
          2090 => x"80",
          2091 => x"70",
          2092 => x"98",
          2093 => x"81",
          2094 => x"84",
          2095 => x"56",
          2096 => x"55",
          2097 => x"97",
          2098 => x"75",
          2099 => x"52",
          2100 => x"51",
          2101 => x"91",
          2102 => x"80",
          2103 => x"80",
          2104 => x"22",
          2105 => x"76",
          2106 => x"81",
          2107 => x"74",
          2108 => x"0c",
          2109 => x"04",
          2110 => x"7a",
          2111 => x"58",
          2112 => x"f0",
          2113 => x"8a",
          2114 => x"06",
          2115 => x"2e",
          2116 => x"58",
          2117 => x"74",
          2118 => x"88",
          2119 => x"73",
          2120 => x"33",
          2121 => x"27",
          2122 => x"16",
          2123 => x"9b",
          2124 => x"2a",
          2125 => x"88",
          2126 => x"58",
          2127 => x"81",
          2128 => x"16",
          2129 => x"0c",
          2130 => x"8a",
          2131 => x"89",
          2132 => x"72",
          2133 => x"38",
          2134 => x"51",
          2135 => x"91",
          2136 => x"54",
          2137 => x"08",
          2138 => x"38",
          2139 => x"d3",
          2140 => x"8b",
          2141 => x"08",
          2142 => x"08",
          2143 => x"82",
          2144 => x"39",
          2145 => x"55",
          2146 => x"cc",
          2147 => x"75",
          2148 => x"3f",
          2149 => x"08",
          2150 => x"73",
          2151 => x"82",
          2152 => x"08",
          2153 => x"38",
          2154 => x"58",
          2155 => x"89",
          2156 => x"08",
          2157 => x"0c",
          2158 => x"06",
          2159 => x"9c",
          2160 => x"58",
          2161 => x"c8",
          2162 => x"0d",
          2163 => x"0d",
          2164 => x"08",
          2165 => x"a0",
          2166 => x"59",
          2167 => x"0a",
          2168 => x"38",
          2169 => x"16",
          2170 => x"98",
          2171 => x"2e",
          2172 => x"75",
          2173 => x"54",
          2174 => x"38",
          2175 => x"81",
          2176 => x"0c",
          2177 => x"98",
          2178 => x"2a",
          2179 => x"59",
          2180 => x"26",
          2181 => x"73",
          2182 => x"84",
          2183 => x"39",
          2184 => x"ff",
          2185 => x"2a",
          2186 => x"72",
          2187 => x"94",
          2188 => x"74",
          2189 => x"3f",
          2190 => x"08",
          2191 => x"81",
          2192 => x"c8",
          2193 => x"84",
          2194 => x"91",
          2195 => x"ff",
          2196 => x"38",
          2197 => x"91",
          2198 => x"26",
          2199 => x"77",
          2200 => x"98",
          2201 => x"53",
          2202 => x"94",
          2203 => x"74",
          2204 => x"3f",
          2205 => x"08",
          2206 => x"91",
          2207 => x"80",
          2208 => x"38",
          2209 => x"d3",
          2210 => x"2e",
          2211 => x"53",
          2212 => x"08",
          2213 => x"38",
          2214 => x"08",
          2215 => x"fb",
          2216 => x"53",
          2217 => x"08",
          2218 => x"94",
          2219 => x"52",
          2220 => x"89",
          2221 => x"c8",
          2222 => x"0c",
          2223 => x"0c",
          2224 => x"06",
          2225 => x"9c",
          2226 => x"53",
          2227 => x"c8",
          2228 => x"0d",
          2229 => x"0d",
          2230 => x"08",
          2231 => x"80",
          2232 => x"fc",
          2233 => x"d3",
          2234 => x"91",
          2235 => x"80",
          2236 => x"d3",
          2237 => x"98",
          2238 => x"77",
          2239 => x"3f",
          2240 => x"08",
          2241 => x"c8",
          2242 => x"38",
          2243 => x"08",
          2244 => x"70",
          2245 => x"55",
          2246 => x"2e",
          2247 => x"83",
          2248 => x"72",
          2249 => x"25",
          2250 => x"53",
          2251 => x"8b",
          2252 => x"57",
          2253 => x"9a",
          2254 => x"80",
          2255 => x"75",
          2256 => x"3f",
          2257 => x"08",
          2258 => x"c8",
          2259 => x"ff",
          2260 => x"84",
          2261 => x"06",
          2262 => x"54",
          2263 => x"c8",
          2264 => x"0d",
          2265 => x"0d",
          2266 => x"52",
          2267 => x"3f",
          2268 => x"08",
          2269 => x"06",
          2270 => x"51",
          2271 => x"83",
          2272 => x"06",
          2273 => x"14",
          2274 => x"3f",
          2275 => x"08",
          2276 => x"07",
          2277 => x"d3",
          2278 => x"3d",
          2279 => x"3d",
          2280 => x"70",
          2281 => x"06",
          2282 => x"53",
          2283 => x"ab",
          2284 => x"33",
          2285 => x"83",
          2286 => x"06",
          2287 => x"90",
          2288 => x"15",
          2289 => x"3f",
          2290 => x"04",
          2291 => x"7b",
          2292 => x"84",
          2293 => x"58",
          2294 => x"80",
          2295 => x"38",
          2296 => x"52",
          2297 => x"df",
          2298 => x"c8",
          2299 => x"d3",
          2300 => x"f1",
          2301 => x"08",
          2302 => x"53",
          2303 => x"84",
          2304 => x"39",
          2305 => x"8b",
          2306 => x"bf",
          2307 => x"ff",
          2308 => x"51",
          2309 => x"17",
          2310 => x"e5",
          2311 => x"76",
          2312 => x"30",
          2313 => x"9f",
          2314 => x"55",
          2315 => x"80",
          2316 => x"76",
          2317 => x"38",
          2318 => x"06",
          2319 => x"88",
          2320 => x"06",
          2321 => x"54",
          2322 => x"99",
          2323 => x"75",
          2324 => x"3f",
          2325 => x"08",
          2326 => x"c8",
          2327 => x"98",
          2328 => x"fc",
          2329 => x"2e",
          2330 => x"0b",
          2331 => x"77",
          2332 => x"0c",
          2333 => x"04",
          2334 => x"7a",
          2335 => x"56",
          2336 => x"51",
          2337 => x"91",
          2338 => x"54",
          2339 => x"08",
          2340 => x"86",
          2341 => x"80",
          2342 => x"16",
          2343 => x"51",
          2344 => x"91",
          2345 => x"57",
          2346 => x"08",
          2347 => x"9c",
          2348 => x"33",
          2349 => x"80",
          2350 => x"9c",
          2351 => x"11",
          2352 => x"55",
          2353 => x"17",
          2354 => x"33",
          2355 => x"70",
          2356 => x"55",
          2357 => x"38",
          2358 => x"16",
          2359 => x"ea",
          2360 => x"d3",
          2361 => x"2e",
          2362 => x"52",
          2363 => x"dd",
          2364 => x"c8",
          2365 => x"d3",
          2366 => x"2e",
          2367 => x"76",
          2368 => x"d3",
          2369 => x"3d",
          2370 => x"3d",
          2371 => x"08",
          2372 => x"52",
          2373 => x"bd",
          2374 => x"c8",
          2375 => x"d3",
          2376 => x"38",
          2377 => x"52",
          2378 => x"9b",
          2379 => x"c8",
          2380 => x"d3",
          2381 => x"38",
          2382 => x"d3",
          2383 => x"9c",
          2384 => x"e9",
          2385 => x"53",
          2386 => x"9c",
          2387 => x"e8",
          2388 => x"0b",
          2389 => x"74",
          2390 => x"0c",
          2391 => x"04",
          2392 => x"76",
          2393 => x"12",
          2394 => x"53",
          2395 => x"d7",
          2396 => x"c8",
          2397 => x"d3",
          2398 => x"38",
          2399 => x"53",
          2400 => x"81",
          2401 => x"34",
          2402 => x"c8",
          2403 => x"0d",
          2404 => x"0d",
          2405 => x"57",
          2406 => x"17",
          2407 => x"08",
          2408 => x"89",
          2409 => x"55",
          2410 => x"08",
          2411 => x"81",
          2412 => x"52",
          2413 => x"ad",
          2414 => x"2e",
          2415 => x"84",
          2416 => x"53",
          2417 => x"09",
          2418 => x"38",
          2419 => x"05",
          2420 => x"81",
          2421 => x"15",
          2422 => x"88",
          2423 => x"81",
          2424 => x"15",
          2425 => x"27",
          2426 => x"15",
          2427 => x"80",
          2428 => x"34",
          2429 => x"52",
          2430 => x"88",
          2431 => x"17",
          2432 => x"51",
          2433 => x"91",
          2434 => x"76",
          2435 => x"08",
          2436 => x"e6",
          2437 => x"d3",
          2438 => x"17",
          2439 => x"08",
          2440 => x"e5",
          2441 => x"d3",
          2442 => x"17",
          2443 => x"0d",
          2444 => x"0d",
          2445 => x"7f",
          2446 => x"5a",
          2447 => x"a0",
          2448 => x"e7",
          2449 => x"70",
          2450 => x"79",
          2451 => x"73",
          2452 => x"81",
          2453 => x"38",
          2454 => x"33",
          2455 => x"ae",
          2456 => x"70",
          2457 => x"82",
          2458 => x"51",
          2459 => x"54",
          2460 => x"7a",
          2461 => x"74",
          2462 => x"58",
          2463 => x"af",
          2464 => x"77",
          2465 => x"70",
          2466 => x"06",
          2467 => x"51",
          2468 => x"74",
          2469 => x"38",
          2470 => x"a0",
          2471 => x"38",
          2472 => x"0c",
          2473 => x"76",
          2474 => x"a0",
          2475 => x"1c",
          2476 => x"82",
          2477 => x"17",
          2478 => x"19",
          2479 => x"a0",
          2480 => x"8c",
          2481 => x"32",
          2482 => x"80",
          2483 => x"30",
          2484 => x"71",
          2485 => x"53",
          2486 => x"55",
          2487 => x"b5",
          2488 => x"81",
          2489 => x"77",
          2490 => x"51",
          2491 => x"af",
          2492 => x"06",
          2493 => x"5a",
          2494 => x"70",
          2495 => x"55",
          2496 => x"2e",
          2497 => x"83",
          2498 => x"79",
          2499 => x"73",
          2500 => x"bc",
          2501 => x"32",
          2502 => x"80",
          2503 => x"27",
          2504 => x"54",
          2505 => x"a2",
          2506 => x"32",
          2507 => x"ae",
          2508 => x"72",
          2509 => x"9f",
          2510 => x"51",
          2511 => x"74",
          2512 => x"88",
          2513 => x"fe",
          2514 => x"98",
          2515 => x"80",
          2516 => x"75",
          2517 => x"91",
          2518 => x"33",
          2519 => x"51",
          2520 => x"91",
          2521 => x"80",
          2522 => x"78",
          2523 => x"81",
          2524 => x"59",
          2525 => x"d7",
          2526 => x"c8",
          2527 => x"89",
          2528 => x"54",
          2529 => x"86",
          2530 => x"80",
          2531 => x"18",
          2532 => x"34",
          2533 => x"11",
          2534 => x"74",
          2535 => x"58",
          2536 => x"75",
          2537 => x"f0",
          2538 => x"3f",
          2539 => x"08",
          2540 => x"ff",
          2541 => x"73",
          2542 => x"38",
          2543 => x"81",
          2544 => x"54",
          2545 => x"75",
          2546 => x"18",
          2547 => x"39",
          2548 => x"0c",
          2549 => x"80",
          2550 => x"7a",
          2551 => x"81",
          2552 => x"81",
          2553 => x"85",
          2554 => x"54",
          2555 => x"8d",
          2556 => x"86",
          2557 => x"86",
          2558 => x"80",
          2559 => x"1c",
          2560 => x"73",
          2561 => x"0c",
          2562 => x"04",
          2563 => x"78",
          2564 => x"56",
          2565 => x"33",
          2566 => x"72",
          2567 => x"38",
          2568 => x"7a",
          2569 => x"54",
          2570 => x"dc",
          2571 => x"81",
          2572 => x"06",
          2573 => x"2e",
          2574 => x"17",
          2575 => x"0c",
          2576 => x"1a",
          2577 => x"70",
          2578 => x"55",
          2579 => x"09",
          2580 => x"38",
          2581 => x"7a",
          2582 => x"54",
          2583 => x"dc",
          2584 => x"06",
          2585 => x"54",
          2586 => x"53",
          2587 => x"80",
          2588 => x"0c",
          2589 => x"51",
          2590 => x"26",
          2591 => x"80",
          2592 => x"34",
          2593 => x"51",
          2594 => x"91",
          2595 => x"55",
          2596 => x"85",
          2597 => x"39",
          2598 => x"05",
          2599 => x"fb",
          2600 => x"d3",
          2601 => x"91",
          2602 => x"81",
          2603 => x"51",
          2604 => x"91",
          2605 => x"ab",
          2606 => x"55",
          2607 => x"08",
          2608 => x"c2",
          2609 => x"c8",
          2610 => x"09",
          2611 => x"ec",
          2612 => x"2a",
          2613 => x"51",
          2614 => x"2e",
          2615 => x"82",
          2616 => x"06",
          2617 => x"80",
          2618 => x"38",
          2619 => x"ab",
          2620 => x"55",
          2621 => x"73",
          2622 => x"81",
          2623 => x"72",
          2624 => x"55",
          2625 => x"82",
          2626 => x"06",
          2627 => x"ac",
          2628 => x"33",
          2629 => x"70",
          2630 => x"54",
          2631 => x"2e",
          2632 => x"90",
          2633 => x"ff",
          2634 => x"05",
          2635 => x"f4",
          2636 => x"d3",
          2637 => x"17",
          2638 => x"39",
          2639 => x"c8",
          2640 => x"0d",
          2641 => x"0d",
          2642 => x"79",
          2643 => x"54",
          2644 => x"74",
          2645 => x"d0",
          2646 => x"81",
          2647 => x"70",
          2648 => x"30",
          2649 => x"71",
          2650 => x"51",
          2651 => x"70",
          2652 => x"ba",
          2653 => x"06",
          2654 => x"74",
          2655 => x"52",
          2656 => x"26",
          2657 => x"15",
          2658 => x"06",
          2659 => x"59",
          2660 => x"2e",
          2661 => x"80",
          2662 => x"e8",
          2663 => x"10",
          2664 => x"08",
          2665 => x"57",
          2666 => x"81",
          2667 => x"75",
          2668 => x"57",
          2669 => x"12",
          2670 => x"70",
          2671 => x"38",
          2672 => x"81",
          2673 => x"51",
          2674 => x"51",
          2675 => x"89",
          2676 => x"70",
          2677 => x"54",
          2678 => x"74",
          2679 => x"30",
          2680 => x"80",
          2681 => x"2a",
          2682 => x"53",
          2683 => x"b9",
          2684 => x"75",
          2685 => x"30",
          2686 => x"9f",
          2687 => x"2a",
          2688 => x"53",
          2689 => x"2e",
          2690 => x"18",
          2691 => x"25",
          2692 => x"8b",
          2693 => x"24",
          2694 => x"77",
          2695 => x"79",
          2696 => x"91",
          2697 => x"51",
          2698 => x"c8",
          2699 => x"0d",
          2700 => x"0d",
          2701 => x"0b",
          2702 => x"ff",
          2703 => x"0c",
          2704 => x"51",
          2705 => x"84",
          2706 => x"c8",
          2707 => x"38",
          2708 => x"51",
          2709 => x"91",
          2710 => x"83",
          2711 => x"54",
          2712 => x"82",
          2713 => x"09",
          2714 => x"e7",
          2715 => x"b4",
          2716 => x"55",
          2717 => x"2e",
          2718 => x"83",
          2719 => x"73",
          2720 => x"70",
          2721 => x"25",
          2722 => x"51",
          2723 => x"38",
          2724 => x"54",
          2725 => x"2e",
          2726 => x"b5",
          2727 => x"91",
          2728 => x"80",
          2729 => x"de",
          2730 => x"d3",
          2731 => x"91",
          2732 => x"80",
          2733 => x"85",
          2734 => x"84",
          2735 => x"16",
          2736 => x"3f",
          2737 => x"08",
          2738 => x"c8",
          2739 => x"83",
          2740 => x"74",
          2741 => x"0c",
          2742 => x"04",
          2743 => x"60",
          2744 => x"80",
          2745 => x"58",
          2746 => x"0c",
          2747 => x"d5",
          2748 => x"c8",
          2749 => x"56",
          2750 => x"d3",
          2751 => x"87",
          2752 => x"d3",
          2753 => x"10",
          2754 => x"05",
          2755 => x"53",
          2756 => x"80",
          2757 => x"38",
          2758 => x"76",
          2759 => x"75",
          2760 => x"72",
          2761 => x"38",
          2762 => x"51",
          2763 => x"91",
          2764 => x"81",
          2765 => x"81",
          2766 => x"72",
          2767 => x"80",
          2768 => x"73",
          2769 => x"81",
          2770 => x"8a",
          2771 => x"cf",
          2772 => x"86",
          2773 => x"75",
          2774 => x"16",
          2775 => x"81",
          2776 => x"d6",
          2777 => x"d3",
          2778 => x"ff",
          2779 => x"06",
          2780 => x"56",
          2781 => x"38",
          2782 => x"8f",
          2783 => x"2a",
          2784 => x"51",
          2785 => x"72",
          2786 => x"80",
          2787 => x"52",
          2788 => x"3f",
          2789 => x"08",
          2790 => x"57",
          2791 => x"09",
          2792 => x"e4",
          2793 => x"73",
          2794 => x"90",
          2795 => x"10",
          2796 => x"83",
          2797 => x"55",
          2798 => x"57",
          2799 => x"8d",
          2800 => x"16",
          2801 => x"3f",
          2802 => x"08",
          2803 => x"0c",
          2804 => x"83",
          2805 => x"38",
          2806 => x"3d",
          2807 => x"05",
          2808 => x"5b",
          2809 => x"79",
          2810 => x"38",
          2811 => x"51",
          2812 => x"91",
          2813 => x"81",
          2814 => x"81",
          2815 => x"38",
          2816 => x"83",
          2817 => x"38",
          2818 => x"84",
          2819 => x"38",
          2820 => x"81",
          2821 => x"38",
          2822 => x"d9",
          2823 => x"d3",
          2824 => x"ff",
          2825 => x"8d",
          2826 => x"80",
          2827 => x"06",
          2828 => x"80",
          2829 => x"d9",
          2830 => x"d3",
          2831 => x"ff",
          2832 => x"73",
          2833 => x"d8",
          2834 => x"e6",
          2835 => x"c8",
          2836 => x"9c",
          2837 => x"c4",
          2838 => x"16",
          2839 => x"15",
          2840 => x"53",
          2841 => x"81",
          2842 => x"38",
          2843 => x"74",
          2844 => x"c1",
          2845 => x"55",
          2846 => x"16",
          2847 => x"ff",
          2848 => x"72",
          2849 => x"38",
          2850 => x"06",
          2851 => x"2e",
          2852 => x"56",
          2853 => x"80",
          2854 => x"d8",
          2855 => x"d3",
          2856 => x"16",
          2857 => x"c8",
          2858 => x"ff",
          2859 => x"53",
          2860 => x"83",
          2861 => x"c7",
          2862 => x"dd",
          2863 => x"c8",
          2864 => x"ff",
          2865 => x"8d",
          2866 => x"15",
          2867 => x"3f",
          2868 => x"08",
          2869 => x"15",
          2870 => x"3f",
          2871 => x"08",
          2872 => x"06",
          2873 => x"78",
          2874 => x"b3",
          2875 => x"22",
          2876 => x"84",
          2877 => x"56",
          2878 => x"73",
          2879 => x"38",
          2880 => x"52",
          2881 => x"51",
          2882 => x"3f",
          2883 => x"08",
          2884 => x"91",
          2885 => x"80",
          2886 => x"38",
          2887 => x"d3",
          2888 => x"ff",
          2889 => x"26",
          2890 => x"57",
          2891 => x"f5",
          2892 => x"82",
          2893 => x"f5",
          2894 => x"81",
          2895 => x"76",
          2896 => x"db",
          2897 => x"98",
          2898 => x"a0",
          2899 => x"19",
          2900 => x"77",
          2901 => x"0c",
          2902 => x"09",
          2903 => x"38",
          2904 => x"51",
          2905 => x"91",
          2906 => x"83",
          2907 => x"53",
          2908 => x"82",
          2909 => x"15",
          2910 => x"56",
          2911 => x"38",
          2912 => x"51",
          2913 => x"91",
          2914 => x"a8",
          2915 => x"15",
          2916 => x"53",
          2917 => x"15",
          2918 => x"56",
          2919 => x"81",
          2920 => x"15",
          2921 => x"16",
          2922 => x"2e",
          2923 => x"88",
          2924 => x"08",
          2925 => x"39",
          2926 => x"10",
          2927 => x"05",
          2928 => x"98",
          2929 => x"06",
          2930 => x"83",
          2931 => x"2a",
          2932 => x"72",
          2933 => x"26",
          2934 => x"ff",
          2935 => x"0c",
          2936 => x"16",
          2937 => x"0b",
          2938 => x"76",
          2939 => x"81",
          2940 => x"38",
          2941 => x"51",
          2942 => x"91",
          2943 => x"83",
          2944 => x"53",
          2945 => x"09",
          2946 => x"f9",
          2947 => x"52",
          2948 => x"b3",
          2949 => x"c8",
          2950 => x"38",
          2951 => x"08",
          2952 => x"84",
          2953 => x"d5",
          2954 => x"d3",
          2955 => x"ff",
          2956 => x"72",
          2957 => x"2e",
          2958 => x"80",
          2959 => x"15",
          2960 => x"3f",
          2961 => x"08",
          2962 => x"a4",
          2963 => x"81",
          2964 => x"84",
          2965 => x"d5",
          2966 => x"d3",
          2967 => x"8a",
          2968 => x"2e",
          2969 => x"9d",
          2970 => x"15",
          2971 => x"3f",
          2972 => x"08",
          2973 => x"84",
          2974 => x"d5",
          2975 => x"d3",
          2976 => x"16",
          2977 => x"34",
          2978 => x"22",
          2979 => x"72",
          2980 => x"23",
          2981 => x"23",
          2982 => x"16",
          2983 => x"75",
          2984 => x"0c",
          2985 => x"04",
          2986 => x"77",
          2987 => x"73",
          2988 => x"38",
          2989 => x"2e",
          2990 => x"08",
          2991 => x"53",
          2992 => x"a4",
          2993 => x"22",
          2994 => x"57",
          2995 => x"2e",
          2996 => x"94",
          2997 => x"33",
          2998 => x"3f",
          2999 => x"08",
          3000 => x"71",
          3001 => x"55",
          3002 => x"73",
          3003 => x"06",
          3004 => x"08",
          3005 => x"71",
          3006 => x"91",
          3007 => x"87",
          3008 => x"fa",
          3009 => x"ab",
          3010 => x"58",
          3011 => x"05",
          3012 => x"b1",
          3013 => x"c8",
          3014 => x"54",
          3015 => x"d3",
          3016 => x"80",
          3017 => x"d3",
          3018 => x"10",
          3019 => x"05",
          3020 => x"54",
          3021 => x"84",
          3022 => x"34",
          3023 => x"86",
          3024 => x"80",
          3025 => x"10",
          3026 => x"e4",
          3027 => x"0c",
          3028 => x"75",
          3029 => x"38",
          3030 => x"3d",
          3031 => x"05",
          3032 => x"3f",
          3033 => x"08",
          3034 => x"d3",
          3035 => x"3d",
          3036 => x"3d",
          3037 => x"84",
          3038 => x"05",
          3039 => x"89",
          3040 => x"2e",
          3041 => x"76",
          3042 => x"54",
          3043 => x"05",
          3044 => x"84",
          3045 => x"f6",
          3046 => x"d3",
          3047 => x"91",
          3048 => x"84",
          3049 => x"5c",
          3050 => x"3d",
          3051 => x"f0",
          3052 => x"d3",
          3053 => x"91",
          3054 => x"92",
          3055 => x"d7",
          3056 => x"98",
          3057 => x"74",
          3058 => x"38",
          3059 => x"9c",
          3060 => x"80",
          3061 => x"38",
          3062 => x"9c",
          3063 => x"2e",
          3064 => x"8e",
          3065 => x"d4",
          3066 => x"9e",
          3067 => x"c8",
          3068 => x"88",
          3069 => x"39",
          3070 => x"33",
          3071 => x"74",
          3072 => x"38",
          3073 => x"39",
          3074 => x"70",
          3075 => x"55",
          3076 => x"83",
          3077 => x"75",
          3078 => x"76",
          3079 => x"81",
          3080 => x"74",
          3081 => x"a7",
          3082 => x"7a",
          3083 => x"3f",
          3084 => x"08",
          3085 => x"b2",
          3086 => x"8e",
          3087 => x"b9",
          3088 => x"a0",
          3089 => x"34",
          3090 => x"52",
          3091 => x"ce",
          3092 => x"62",
          3093 => x"d2",
          3094 => x"55",
          3095 => x"16",
          3096 => x"2e",
          3097 => x"7a",
          3098 => x"77",
          3099 => x"99",
          3100 => x"53",
          3101 => x"b3",
          3102 => x"c8",
          3103 => x"d3",
          3104 => x"e6",
          3105 => x"7a",
          3106 => x"3f",
          3107 => x"08",
          3108 => x"8c",
          3109 => x"56",
          3110 => x"82",
          3111 => x"b2",
          3112 => x"84",
          3113 => x"06",
          3114 => x"74",
          3115 => x"38",
          3116 => x"39",
          3117 => x"70",
          3118 => x"55",
          3119 => x"8f",
          3120 => x"05",
          3121 => x"55",
          3122 => x"83",
          3123 => x"75",
          3124 => x"76",
          3125 => x"81",
          3126 => x"74",
          3127 => x"38",
          3128 => x"07",
          3129 => x"11",
          3130 => x"0c",
          3131 => x"0c",
          3132 => x"f6",
          3133 => x"74",
          3134 => x"3f",
          3135 => x"08",
          3136 => x"62",
          3137 => x"d0",
          3138 => x"d3",
          3139 => x"19",
          3140 => x"0c",
          3141 => x"84",
          3142 => x"90",
          3143 => x"91",
          3144 => x"9c",
          3145 => x"94",
          3146 => x"80",
          3147 => x"a8",
          3148 => x"98",
          3149 => x"2a",
          3150 => x"51",
          3151 => x"2e",
          3152 => x"8c",
          3153 => x"2e",
          3154 => x"8c",
          3155 => x"19",
          3156 => x"11",
          3157 => x"2b",
          3158 => x"8c",
          3159 => x"5a",
          3160 => x"a5",
          3161 => x"77",
          3162 => x"3f",
          3163 => x"08",
          3164 => x"c8",
          3165 => x"83",
          3166 => x"76",
          3167 => x"81",
          3168 => x"81",
          3169 => x"31",
          3170 => x"70",
          3171 => x"25",
          3172 => x"26",
          3173 => x"55",
          3174 => x"76",
          3175 => x"75",
          3176 => x"78",
          3177 => x"55",
          3178 => x"b9",
          3179 => x"7a",
          3180 => x"3f",
          3181 => x"08",
          3182 => x"56",
          3183 => x"89",
          3184 => x"c8",
          3185 => x"9c",
          3186 => x"81",
          3187 => x"a8",
          3188 => x"81",
          3189 => x"55",
          3190 => x"91",
          3191 => x"80",
          3192 => x"81",
          3193 => x"2e",
          3194 => x"78",
          3195 => x"74",
          3196 => x"0c",
          3197 => x"04",
          3198 => x"7f",
          3199 => x"5f",
          3200 => x"80",
          3201 => x"3d",
          3202 => x"76",
          3203 => x"3f",
          3204 => x"08",
          3205 => x"c8",
          3206 => x"91",
          3207 => x"74",
          3208 => x"38",
          3209 => x"ae",
          3210 => x"33",
          3211 => x"87",
          3212 => x"2e",
          3213 => x"bd",
          3214 => x"91",
          3215 => x"56",
          3216 => x"81",
          3217 => x"34",
          3218 => x"8a",
          3219 => x"91",
          3220 => x"56",
          3221 => x"81",
          3222 => x"34",
          3223 => x"f6",
          3224 => x"91",
          3225 => x"56",
          3226 => x"81",
          3227 => x"34",
          3228 => x"e2",
          3229 => x"08",
          3230 => x"31",
          3231 => x"27",
          3232 => x"59",
          3233 => x"82",
          3234 => x"17",
          3235 => x"ff",
          3236 => x"74",
          3237 => x"7d",
          3238 => x"ff",
          3239 => x"2a",
          3240 => x"7a",
          3241 => x"87",
          3242 => x"08",
          3243 => x"98",
          3244 => x"76",
          3245 => x"3f",
          3246 => x"08",
          3247 => x"27",
          3248 => x"74",
          3249 => x"fb",
          3250 => x"18",
          3251 => x"08",
          3252 => x"d1",
          3253 => x"d3",
          3254 => x"2e",
          3255 => x"91",
          3256 => x"1b",
          3257 => x"5b",
          3258 => x"2e",
          3259 => x"79",
          3260 => x"11",
          3261 => x"56",
          3262 => x"85",
          3263 => x"31",
          3264 => x"77",
          3265 => x"7d",
          3266 => x"52",
          3267 => x"3f",
          3268 => x"08",
          3269 => x"90",
          3270 => x"98",
          3271 => x"74",
          3272 => x"38",
          3273 => x"78",
          3274 => x"7a",
          3275 => x"84",
          3276 => x"17",
          3277 => x"80",
          3278 => x"cc",
          3279 => x"89",
          3280 => x"f9",
          3281 => x"08",
          3282 => x"c9",
          3283 => x"33",
          3284 => x"56",
          3285 => x"25",
          3286 => x"54",
          3287 => x"53",
          3288 => x"7d",
          3289 => x"52",
          3290 => x"3f",
          3291 => x"08",
          3292 => x"90",
          3293 => x"ff",
          3294 => x"90",
          3295 => x"54",
          3296 => x"17",
          3297 => x"11",
          3298 => x"c6",
          3299 => x"d3",
          3300 => x"d7",
          3301 => x"18",
          3302 => x"08",
          3303 => x"84",
          3304 => x"57",
          3305 => x"27",
          3306 => x"56",
          3307 => x"17",
          3308 => x"06",
          3309 => x"52",
          3310 => x"ec",
          3311 => x"31",
          3312 => x"7e",
          3313 => x"94",
          3314 => x"94",
          3315 => x"59",
          3316 => x"38",
          3317 => x"91",
          3318 => x"8f",
          3319 => x"f3",
          3320 => x"62",
          3321 => x"5f",
          3322 => x"7d",
          3323 => x"fc",
          3324 => x"51",
          3325 => x"91",
          3326 => x"55",
          3327 => x"08",
          3328 => x"17",
          3329 => x"80",
          3330 => x"74",
          3331 => x"39",
          3332 => x"70",
          3333 => x"81",
          3334 => x"56",
          3335 => x"80",
          3336 => x"38",
          3337 => x"0b",
          3338 => x"82",
          3339 => x"39",
          3340 => x"18",
          3341 => x"83",
          3342 => x"0b",
          3343 => x"81",
          3344 => x"39",
          3345 => x"18",
          3346 => x"83",
          3347 => x"0b",
          3348 => x"81",
          3349 => x"39",
          3350 => x"18",
          3351 => x"83",
          3352 => x"17",
          3353 => x"74",
          3354 => x"27",
          3355 => x"17",
          3356 => x"78",
          3357 => x"8c",
          3358 => x"08",
          3359 => x"06",
          3360 => x"82",
          3361 => x"8a",
          3362 => x"05",
          3363 => x"06",
          3364 => x"80",
          3365 => x"96",
          3366 => x"08",
          3367 => x"38",
          3368 => x"51",
          3369 => x"91",
          3370 => x"55",
          3371 => x"17",
          3372 => x"51",
          3373 => x"91",
          3374 => x"55",
          3375 => x"82",
          3376 => x"81",
          3377 => x"38",
          3378 => x"fe",
          3379 => x"98",
          3380 => x"17",
          3381 => x"74",
          3382 => x"90",
          3383 => x"98",
          3384 => x"74",
          3385 => x"38",
          3386 => x"17",
          3387 => x"17",
          3388 => x"11",
          3389 => x"c5",
          3390 => x"d3",
          3391 => x"ba",
          3392 => x"33",
          3393 => x"55",
          3394 => x"34",
          3395 => x"52",
          3396 => x"a9",
          3397 => x"c8",
          3398 => x"fe",
          3399 => x"d3",
          3400 => x"79",
          3401 => x"58",
          3402 => x"80",
          3403 => x"1b",
          3404 => x"22",
          3405 => x"74",
          3406 => x"38",
          3407 => x"5a",
          3408 => x"53",
          3409 => x"81",
          3410 => x"55",
          3411 => x"91",
          3412 => x"fd",
          3413 => x"17",
          3414 => x"55",
          3415 => x"9b",
          3416 => x"53",
          3417 => x"29",
          3418 => x"17",
          3419 => x"3f",
          3420 => x"80",
          3421 => x"74",
          3422 => x"79",
          3423 => x"80",
          3424 => x"17",
          3425 => x"a1",
          3426 => x"08",
          3427 => x"27",
          3428 => x"54",
          3429 => x"17",
          3430 => x"11",
          3431 => x"c2",
          3432 => x"d3",
          3433 => x"b0",
          3434 => x"18",
          3435 => x"08",
          3436 => x"84",
          3437 => x"57",
          3438 => x"27",
          3439 => x"56",
          3440 => x"52",
          3441 => x"83",
          3442 => x"a8",
          3443 => x"d8",
          3444 => x"33",
          3445 => x"55",
          3446 => x"34",
          3447 => x"7d",
          3448 => x"0c",
          3449 => x"19",
          3450 => x"94",
          3451 => x"1a",
          3452 => x"5d",
          3453 => x"27",
          3454 => x"55",
          3455 => x"0c",
          3456 => x"38",
          3457 => x"80",
          3458 => x"74",
          3459 => x"80",
          3460 => x"d3",
          3461 => x"3d",
          3462 => x"3d",
          3463 => x"3d",
          3464 => x"70",
          3465 => x"80",
          3466 => x"c8",
          3467 => x"d3",
          3468 => x"aa",
          3469 => x"33",
          3470 => x"70",
          3471 => x"56",
          3472 => x"2e",
          3473 => x"75",
          3474 => x"74",
          3475 => x"38",
          3476 => x"18",
          3477 => x"18",
          3478 => x"11",
          3479 => x"c2",
          3480 => x"55",
          3481 => x"08",
          3482 => x"90",
          3483 => x"ff",
          3484 => x"90",
          3485 => x"18",
          3486 => x"51",
          3487 => x"91",
          3488 => x"57",
          3489 => x"08",
          3490 => x"a4",
          3491 => x"11",
          3492 => x"56",
          3493 => x"17",
          3494 => x"08",
          3495 => x"77",
          3496 => x"fa",
          3497 => x"08",
          3498 => x"51",
          3499 => x"82",
          3500 => x"52",
          3501 => x"c5",
          3502 => x"52",
          3503 => x"c5",
          3504 => x"55",
          3505 => x"16",
          3506 => x"c8",
          3507 => x"d3",
          3508 => x"19",
          3509 => x"06",
          3510 => x"90",
          3511 => x"55",
          3512 => x"c8",
          3513 => x"0d",
          3514 => x"0d",
          3515 => x"54",
          3516 => x"91",
          3517 => x"53",
          3518 => x"08",
          3519 => x"3d",
          3520 => x"73",
          3521 => x"3f",
          3522 => x"08",
          3523 => x"c8",
          3524 => x"91",
          3525 => x"74",
          3526 => x"d3",
          3527 => x"3d",
          3528 => x"3d",
          3529 => x"51",
          3530 => x"8b",
          3531 => x"91",
          3532 => x"24",
          3533 => x"d3",
          3534 => x"d3",
          3535 => x"53",
          3536 => x"c8",
          3537 => x"0d",
          3538 => x"0d",
          3539 => x"3d",
          3540 => x"94",
          3541 => x"84",
          3542 => x"c8",
          3543 => x"d3",
          3544 => x"df",
          3545 => x"63",
          3546 => x"d4",
          3547 => x"9c",
          3548 => x"c8",
          3549 => x"d3",
          3550 => x"38",
          3551 => x"05",
          3552 => x"2b",
          3553 => x"80",
          3554 => x"76",
          3555 => x"0c",
          3556 => x"02",
          3557 => x"70",
          3558 => x"81",
          3559 => x"56",
          3560 => x"93",
          3561 => x"53",
          3562 => x"d7",
          3563 => x"d3",
          3564 => x"15",
          3565 => x"85",
          3566 => x"2e",
          3567 => x"83",
          3568 => x"74",
          3569 => x"0c",
          3570 => x"04",
          3571 => x"a3",
          3572 => x"3d",
          3573 => x"80",
          3574 => x"53",
          3575 => x"b8",
          3576 => x"3d",
          3577 => x"3f",
          3578 => x"08",
          3579 => x"c8",
          3580 => x"38",
          3581 => x"7f",
          3582 => x"4a",
          3583 => x"59",
          3584 => x"81",
          3585 => x"3d",
          3586 => x"40",
          3587 => x"52",
          3588 => x"e4",
          3589 => x"c8",
          3590 => x"d3",
          3591 => x"de",
          3592 => x"7e",
          3593 => x"3f",
          3594 => x"08",
          3595 => x"c8",
          3596 => x"38",
          3597 => x"51",
          3598 => x"91",
          3599 => x"48",
          3600 => x"51",
          3601 => x"91",
          3602 => x"57",
          3603 => x"08",
          3604 => x"7c",
          3605 => x"73",
          3606 => x"3f",
          3607 => x"08",
          3608 => x"c8",
          3609 => x"6c",
          3610 => x"d5",
          3611 => x"d3",
          3612 => x"2e",
          3613 => x"52",
          3614 => x"d1",
          3615 => x"c8",
          3616 => x"d3",
          3617 => x"2e",
          3618 => x"84",
          3619 => x"06",
          3620 => x"57",
          3621 => x"38",
          3622 => x"bc",
          3623 => x"05",
          3624 => x"3f",
          3625 => x"70",
          3626 => x"11",
          3627 => x"57",
          3628 => x"80",
          3629 => x"81",
          3630 => x"81",
          3631 => x"55",
          3632 => x"38",
          3633 => x"78",
          3634 => x"38",
          3635 => x"39",
          3636 => x"99",
          3637 => x"ff",
          3638 => x"08",
          3639 => x"70",
          3640 => x"56",
          3641 => x"33",
          3642 => x"eb",
          3643 => x"a3",
          3644 => x"55",
          3645 => x"34",
          3646 => x"fe",
          3647 => x"81",
          3648 => x"7c",
          3649 => x"06",
          3650 => x"19",
          3651 => x"11",
          3652 => x"74",
          3653 => x"91",
          3654 => x"70",
          3655 => x"bb",
          3656 => x"08",
          3657 => x"52",
          3658 => x"58",
          3659 => x"8d",
          3660 => x"70",
          3661 => x"51",
          3662 => x"f5",
          3663 => x"54",
          3664 => x"a5",
          3665 => x"77",
          3666 => x"38",
          3667 => x"73",
          3668 => x"81",
          3669 => x"81",
          3670 => x"78",
          3671 => x"ba",
          3672 => x"05",
          3673 => x"18",
          3674 => x"38",
          3675 => x"96",
          3676 => x"08",
          3677 => x"5a",
          3678 => x"7a",
          3679 => x"5c",
          3680 => x"26",
          3681 => x"7a",
          3682 => x"d3",
          3683 => x"3d",
          3684 => x"3d",
          3685 => x"90",
          3686 => x"54",
          3687 => x"57",
          3688 => x"91",
          3689 => x"5a",
          3690 => x"08",
          3691 => x"17",
          3692 => x"80",
          3693 => x"79",
          3694 => x"39",
          3695 => x"78",
          3696 => x"90",
          3697 => x"81",
          3698 => x"06",
          3699 => x"74",
          3700 => x"17",
          3701 => x"17",
          3702 => x"70",
          3703 => x"5b",
          3704 => x"82",
          3705 => x"8a",
          3706 => x"89",
          3707 => x"55",
          3708 => x"b6",
          3709 => x"ff",
          3710 => x"96",
          3711 => x"d3",
          3712 => x"17",
          3713 => x"53",
          3714 => x"96",
          3715 => x"d3",
          3716 => x"26",
          3717 => x"30",
          3718 => x"18",
          3719 => x"18",
          3720 => x"18",
          3721 => x"80",
          3722 => x"17",
          3723 => x"be",
          3724 => x"76",
          3725 => x"3f",
          3726 => x"08",
          3727 => x"c8",
          3728 => x"09",
          3729 => x"38",
          3730 => x"18",
          3731 => x"82",
          3732 => x"d3",
          3733 => x"2e",
          3734 => x"8b",
          3735 => x"91",
          3736 => x"55",
          3737 => x"91",
          3738 => x"88",
          3739 => x"98",
          3740 => x"80",
          3741 => x"38",
          3742 => x"80",
          3743 => x"79",
          3744 => x"08",
          3745 => x"0c",
          3746 => x"70",
          3747 => x"81",
          3748 => x"5d",
          3749 => x"2e",
          3750 => x"52",
          3751 => x"be",
          3752 => x"c8",
          3753 => x"d3",
          3754 => x"38",
          3755 => x"08",
          3756 => x"75",
          3757 => x"c2",
          3758 => x"d3",
          3759 => x"75",
          3760 => x"e1",
          3761 => x"27",
          3762 => x"55",
          3763 => x"76",
          3764 => x"82",
          3765 => x"34",
          3766 => x"d8",
          3767 => x"18",
          3768 => x"26",
          3769 => x"94",
          3770 => x"94",
          3771 => x"83",
          3772 => x"74",
          3773 => x"38",
          3774 => x"51",
          3775 => x"91",
          3776 => x"8b",
          3777 => x"91",
          3778 => x"55",
          3779 => x"77",
          3780 => x"d3",
          3781 => x"5b",
          3782 => x"94",
          3783 => x"92",
          3784 => x"08",
          3785 => x"90",
          3786 => x"c0",
          3787 => x"90",
          3788 => x"17",
          3789 => x"06",
          3790 => x"2e",
          3791 => x"9c",
          3792 => x"2e",
          3793 => x"90",
          3794 => x"98",
          3795 => x"74",
          3796 => x"38",
          3797 => x"17",
          3798 => x"17",
          3799 => x"11",
          3800 => x"ff",
          3801 => x"91",
          3802 => x"80",
          3803 => x"81",
          3804 => x"34",
          3805 => x"39",
          3806 => x"80",
          3807 => x"74",
          3808 => x"81",
          3809 => x"a8",
          3810 => x"81",
          3811 => x"55",
          3812 => x"3f",
          3813 => x"08",
          3814 => x"38",
          3815 => x"18",
          3816 => x"90",
          3817 => x"91",
          3818 => x"55",
          3819 => x"9c",
          3820 => x"55",
          3821 => x"c8",
          3822 => x"0d",
          3823 => x"0d",
          3824 => x"54",
          3825 => x"81",
          3826 => x"53",
          3827 => x"05",
          3828 => x"84",
          3829 => x"84",
          3830 => x"c8",
          3831 => x"d3",
          3832 => x"ef",
          3833 => x"0c",
          3834 => x"51",
          3835 => x"91",
          3836 => x"55",
          3837 => x"08",
          3838 => x"ab",
          3839 => x"98",
          3840 => x"80",
          3841 => x"38",
          3842 => x"70",
          3843 => x"81",
          3844 => x"57",
          3845 => x"93",
          3846 => x"08",
          3847 => x"ce",
          3848 => x"d3",
          3849 => x"17",
          3850 => x"85",
          3851 => x"38",
          3852 => x"14",
          3853 => x"23",
          3854 => x"51",
          3855 => x"91",
          3856 => x"55",
          3857 => x"09",
          3858 => x"38",
          3859 => x"80",
          3860 => x"80",
          3861 => x"54",
          3862 => x"c8",
          3863 => x"0d",
          3864 => x"0d",
          3865 => x"fc",
          3866 => x"52",
          3867 => x"3f",
          3868 => x"08",
          3869 => x"c8",
          3870 => x"91",
          3871 => x"74",
          3872 => x"d3",
          3873 => x"3d",
          3874 => x"3d",
          3875 => x"89",
          3876 => x"54",
          3877 => x"54",
          3878 => x"91",
          3879 => x"53",
          3880 => x"08",
          3881 => x"74",
          3882 => x"d3",
          3883 => x"73",
          3884 => x"3f",
          3885 => x"08",
          3886 => x"80",
          3887 => x"ce",
          3888 => x"d3",
          3889 => x"91",
          3890 => x"84",
          3891 => x"06",
          3892 => x"53",
          3893 => x"74",
          3894 => x"d1",
          3895 => x"52",
          3896 => x"e9",
          3897 => x"c8",
          3898 => x"d3",
          3899 => x"2e",
          3900 => x"83",
          3901 => x"72",
          3902 => x"0c",
          3903 => x"04",
          3904 => x"64",
          3905 => x"88",
          3906 => x"95",
          3907 => x"db",
          3908 => x"d3",
          3909 => x"91",
          3910 => x"b5",
          3911 => x"73",
          3912 => x"3f",
          3913 => x"08",
          3914 => x"c8",
          3915 => x"02",
          3916 => x"33",
          3917 => x"55",
          3918 => x"25",
          3919 => x"55",
          3920 => x"80",
          3921 => x"75",
          3922 => x"d4",
          3923 => x"c1",
          3924 => x"d3",
          3925 => x"3d",
          3926 => x"3d",
          3927 => x"55",
          3928 => x"90",
          3929 => x"52",
          3930 => x"da",
          3931 => x"d3",
          3932 => x"91",
          3933 => x"82",
          3934 => x"74",
          3935 => x"98",
          3936 => x"05",
          3937 => x"15",
          3938 => x"93",
          3939 => x"08",
          3940 => x"e9",
          3941 => x"81",
          3942 => x"59",
          3943 => x"80",
          3944 => x"56",
          3945 => x"81",
          3946 => x"06",
          3947 => x"82",
          3948 => x"75",
          3949 => x"f0",
          3950 => x"bc",
          3951 => x"d3",
          3952 => x"2e",
          3953 => x"d3",
          3954 => x"2e",
          3955 => x"d3",
          3956 => x"70",
          3957 => x"08",
          3958 => x"78",
          3959 => x"7d",
          3960 => x"54",
          3961 => x"76",
          3962 => x"80",
          3963 => x"98",
          3964 => x"12",
          3965 => x"54",
          3966 => x"98",
          3967 => x"81",
          3968 => x"58",
          3969 => x"3f",
          3970 => x"08",
          3971 => x"c8",
          3972 => x"38",
          3973 => x"51",
          3974 => x"2e",
          3975 => x"a0",
          3976 => x"b4",
          3977 => x"b5",
          3978 => x"d3",
          3979 => x"ff",
          3980 => x"30",
          3981 => x"19",
          3982 => x"59",
          3983 => x"39",
          3984 => x"05",
          3985 => x"ea",
          3986 => x"c8",
          3987 => x"06",
          3988 => x"80",
          3989 => x"18",
          3990 => x"54",
          3991 => x"06",
          3992 => x"55",
          3993 => x"38",
          3994 => x"7a",
          3995 => x"0c",
          3996 => x"11",
          3997 => x"55",
          3998 => x"16",
          3999 => x"d3",
          4000 => x"3d",
          4001 => x"3d",
          4002 => x"3d",
          4003 => x"70",
          4004 => x"94",
          4005 => x"c8",
          4006 => x"d3",
          4007 => x"38",
          4008 => x"57",
          4009 => x"86",
          4010 => x"81",
          4011 => x"18",
          4012 => x"2a",
          4013 => x"51",
          4014 => x"56",
          4015 => x"81",
          4016 => x"18",
          4017 => x"08",
          4018 => x"38",
          4019 => x"9a",
          4020 => x"88",
          4021 => x"77",
          4022 => x"cf",
          4023 => x"c8",
          4024 => x"0b",
          4025 => x"80",
          4026 => x"18",
          4027 => x"51",
          4028 => x"3f",
          4029 => x"08",
          4030 => x"08",
          4031 => x"30",
          4032 => x"80",
          4033 => x"58",
          4034 => x"c8",
          4035 => x"09",
          4036 => x"38",
          4037 => x"9b",
          4038 => x"75",
          4039 => x"27",
          4040 => x"18",
          4041 => x"52",
          4042 => x"bd",
          4043 => x"d3",
          4044 => x"94",
          4045 => x"19",
          4046 => x"33",
          4047 => x"55",
          4048 => x"34",
          4049 => x"74",
          4050 => x"74",
          4051 => x"38",
          4052 => x"18",
          4053 => x"18",
          4054 => x"11",
          4055 => x"ff",
          4056 => x"91",
          4057 => x"80",
          4058 => x"81",
          4059 => x"90",
          4060 => x"ff",
          4061 => x"90",
          4062 => x"80",
          4063 => x"76",
          4064 => x"76",
          4065 => x"76",
          4066 => x"d3",
          4067 => x"3d",
          4068 => x"3d",
          4069 => x"8c",
          4070 => x"d5",
          4071 => x"9f",
          4072 => x"05",
          4073 => x"51",
          4074 => x"91",
          4075 => x"56",
          4076 => x"08",
          4077 => x"91",
          4078 => x"ff",
          4079 => x"77",
          4080 => x"9f",
          4081 => x"51",
          4082 => x"91",
          4083 => x"91",
          4084 => x"56",
          4085 => x"3f",
          4086 => x"38",
          4087 => x"05",
          4088 => x"2a",
          4089 => x"51",
          4090 => x"80",
          4091 => x"86",
          4092 => x"95",
          4093 => x"98",
          4094 => x"f5",
          4095 => x"f7",
          4096 => x"98",
          4097 => x"73",
          4098 => x"38",
          4099 => x"39",
          4100 => x"05",
          4101 => x"54",
          4102 => x"83",
          4103 => x"75",
          4104 => x"6a",
          4105 => x"c6",
          4106 => x"d3",
          4107 => x"84",
          4108 => x"05",
          4109 => x"2a",
          4110 => x"51",
          4111 => x"73",
          4112 => x"e5",
          4113 => x"9c",
          4114 => x"a5",
          4115 => x"55",
          4116 => x"08",
          4117 => x"d1",
          4118 => x"a0",
          4119 => x"91",
          4120 => x"76",
          4121 => x"a4",
          4122 => x"85",
          4123 => x"89",
          4124 => x"54",
          4125 => x"91",
          4126 => x"56",
          4127 => x"08",
          4128 => x"91",
          4129 => x"52",
          4130 => x"c0",
          4131 => x"c8",
          4132 => x"d3",
          4133 => x"38",
          4134 => x"84",
          4135 => x"70",
          4136 => x"2c",
          4137 => x"56",
          4138 => x"dd",
          4139 => x"a8",
          4140 => x"bd",
          4141 => x"d4",
          4142 => x"a4",
          4143 => x"c8",
          4144 => x"c8",
          4145 => x"91",
          4146 => x"07",
          4147 => x"30",
          4148 => x"9f",
          4149 => x"52",
          4150 => x"56",
          4151 => x"9b",
          4152 => x"ac",
          4153 => x"89",
          4154 => x"76",
          4155 => x"d4",
          4156 => x"ba",
          4157 => x"d3",
          4158 => x"75",
          4159 => x"51",
          4160 => x"3f",
          4161 => x"08",
          4162 => x"b0",
          4163 => x"e1",
          4164 => x"d3",
          4165 => x"3d",
          4166 => x"3d",
          4167 => x"98",
          4168 => x"52",
          4169 => x"d3",
          4170 => x"d3",
          4171 => x"91",
          4172 => x"82",
          4173 => x"5d",
          4174 => x"3d",
          4175 => x"cd",
          4176 => x"d3",
          4177 => x"91",
          4178 => x"83",
          4179 => x"74",
          4180 => x"81",
          4181 => x"38",
          4182 => x"05",
          4183 => x"2a",
          4184 => x"51",
          4185 => x"80",
          4186 => x"86",
          4187 => x"2e",
          4188 => x"81",
          4189 => x"59",
          4190 => x"3d",
          4191 => x"ff",
          4192 => x"91",
          4193 => x"56",
          4194 => x"d3",
          4195 => x"2e",
          4196 => x"83",
          4197 => x"75",
          4198 => x"81",
          4199 => x"82",
          4200 => x"2e",
          4201 => x"83",
          4202 => x"82",
          4203 => x"57",
          4204 => x"38",
          4205 => x"51",
          4206 => x"3f",
          4207 => x"08",
          4208 => x"c8",
          4209 => x"38",
          4210 => x"52",
          4211 => x"ff",
          4212 => x"77",
          4213 => x"b4",
          4214 => x"54",
          4215 => x"15",
          4216 => x"80",
          4217 => x"ff",
          4218 => x"75",
          4219 => x"52",
          4220 => x"aa",
          4221 => x"b4",
          4222 => x"d4",
          4223 => x"af",
          4224 => x"54",
          4225 => x"d5",
          4226 => x"53",
          4227 => x"52",
          4228 => x"8a",
          4229 => x"81",
          4230 => x"34",
          4231 => x"05",
          4232 => x"3f",
          4233 => x"08",
          4234 => x"c8",
          4235 => x"76",
          4236 => x"05",
          4237 => x"c1",
          4238 => x"63",
          4239 => x"c2",
          4240 => x"54",
          4241 => x"15",
          4242 => x"81",
          4243 => x"34",
          4244 => x"b1",
          4245 => x"d3",
          4246 => x"8e",
          4247 => x"75",
          4248 => x"c4",
          4249 => x"b7",
          4250 => x"91",
          4251 => x"98",
          4252 => x"db",
          4253 => x"3d",
          4254 => x"cd",
          4255 => x"53",
          4256 => x"84",
          4257 => x"3d",
          4258 => x"3f",
          4259 => x"08",
          4260 => x"c8",
          4261 => x"38",
          4262 => x"3d",
          4263 => x"3d",
          4264 => x"ca",
          4265 => x"d3",
          4266 => x"91",
          4267 => x"82",
          4268 => x"81",
          4269 => x"81",
          4270 => x"73",
          4271 => x"38",
          4272 => x"82",
          4273 => x"53",
          4274 => x"52",
          4275 => x"88",
          4276 => x"ad",
          4277 => x"53",
          4278 => x"05",
          4279 => x"70",
          4280 => x"ad",
          4281 => x"3d",
          4282 => x"51",
          4283 => x"91",
          4284 => x"55",
          4285 => x"08",
          4286 => x"6e",
          4287 => x"06",
          4288 => x"55",
          4289 => x"08",
          4290 => x"88",
          4291 => x"2e",
          4292 => x"81",
          4293 => x"3d",
          4294 => x"51",
          4295 => x"91",
          4296 => x"55",
          4297 => x"08",
          4298 => x"67",
          4299 => x"a7",
          4300 => x"05",
          4301 => x"51",
          4302 => x"3f",
          4303 => x"33",
          4304 => x"8b",
          4305 => x"84",
          4306 => x"06",
          4307 => x"73",
          4308 => x"a0",
          4309 => x"8b",
          4310 => x"54",
          4311 => x"15",
          4312 => x"33",
          4313 => x"70",
          4314 => x"55",
          4315 => x"2e",
          4316 => x"6d",
          4317 => x"d5",
          4318 => x"77",
          4319 => x"e5",
          4320 => x"c8",
          4321 => x"51",
          4322 => x"3f",
          4323 => x"d3",
          4324 => x"2e",
          4325 => x"d3",
          4326 => x"77",
          4327 => x"a7",
          4328 => x"c8",
          4329 => x"19",
          4330 => x"d3",
          4331 => x"38",
          4332 => x"54",
          4333 => x"09",
          4334 => x"38",
          4335 => x"52",
          4336 => x"bf",
          4337 => x"54",
          4338 => x"15",
          4339 => x"38",
          4340 => x"05",
          4341 => x"3f",
          4342 => x"08",
          4343 => x"c8",
          4344 => x"77",
          4345 => x"a6",
          4346 => x"c8",
          4347 => x"91",
          4348 => x"a7",
          4349 => x"ed",
          4350 => x"80",
          4351 => x"02",
          4352 => x"df",
          4353 => x"57",
          4354 => x"3d",
          4355 => x"96",
          4356 => x"c8",
          4357 => x"c8",
          4358 => x"d3",
          4359 => x"d4",
          4360 => x"65",
          4361 => x"d4",
          4362 => x"e0",
          4363 => x"c8",
          4364 => x"d3",
          4365 => x"38",
          4366 => x"05",
          4367 => x"06",
          4368 => x"2e",
          4369 => x"55",
          4370 => x"75",
          4371 => x"71",
          4372 => x"33",
          4373 => x"74",
          4374 => x"57",
          4375 => x"8b",
          4376 => x"54",
          4377 => x"15",
          4378 => x"ff",
          4379 => x"91",
          4380 => x"55",
          4381 => x"c8",
          4382 => x"0d",
          4383 => x"0d",
          4384 => x"53",
          4385 => x"05",
          4386 => x"51",
          4387 => x"91",
          4388 => x"55",
          4389 => x"08",
          4390 => x"77",
          4391 => x"94",
          4392 => x"51",
          4393 => x"91",
          4394 => x"55",
          4395 => x"08",
          4396 => x"80",
          4397 => x"81",
          4398 => x"73",
          4399 => x"38",
          4400 => x"a9",
          4401 => x"22",
          4402 => x"70",
          4403 => x"07",
          4404 => x"7f",
          4405 => x"ff",
          4406 => x"77",
          4407 => x"83",
          4408 => x"51",
          4409 => x"3f",
          4410 => x"08",
          4411 => x"d3",
          4412 => x"3d",
          4413 => x"3d",
          4414 => x"5c",
          4415 => x"98",
          4416 => x"52",
          4417 => x"cb",
          4418 => x"d3",
          4419 => x"d3",
          4420 => x"70",
          4421 => x"08",
          4422 => x"7b",
          4423 => x"07",
          4424 => x"06",
          4425 => x"56",
          4426 => x"2e",
          4427 => x"7b",
          4428 => x"80",
          4429 => x"70",
          4430 => x"b7",
          4431 => x"d3",
          4432 => x"91",
          4433 => x"80",
          4434 => x"52",
          4435 => x"bc",
          4436 => x"d3",
          4437 => x"91",
          4438 => x"bb",
          4439 => x"c8",
          4440 => x"c8",
          4441 => x"58",
          4442 => x"81",
          4443 => x"56",
          4444 => x"33",
          4445 => x"18",
          4446 => x"27",
          4447 => x"19",
          4448 => x"34",
          4449 => x"8f",
          4450 => x"79",
          4451 => x"51",
          4452 => x"a0",
          4453 => x"75",
          4454 => x"81",
          4455 => x"80",
          4456 => x"56",
          4457 => x"77",
          4458 => x"7c",
          4459 => x"07",
          4460 => x"06",
          4461 => x"55",
          4462 => x"bc",
          4463 => x"11",
          4464 => x"ff",
          4465 => x"91",
          4466 => x"56",
          4467 => x"08",
          4468 => x"70",
          4469 => x"80",
          4470 => x"83",
          4471 => x"80",
          4472 => x"84",
          4473 => x"a7",
          4474 => x"b4",
          4475 => x"a6",
          4476 => x"d3",
          4477 => x"0c",
          4478 => x"c8",
          4479 => x"0d",
          4480 => x"0d",
          4481 => x"3d",
          4482 => x"52",
          4483 => x"c9",
          4484 => x"d3",
          4485 => x"91",
          4486 => x"83",
          4487 => x"53",
          4488 => x"3d",
          4489 => x"51",
          4490 => x"3f",
          4491 => x"71",
          4492 => x"55",
          4493 => x"27",
          4494 => x"74",
          4495 => x"05",
          4496 => x"ff",
          4497 => x"ff",
          4498 => x"91",
          4499 => x"80",
          4500 => x"6a",
          4501 => x"53",
          4502 => x"a7",
          4503 => x"d3",
          4504 => x"2e",
          4505 => x"88",
          4506 => x"6b",
          4507 => x"56",
          4508 => x"56",
          4509 => x"54",
          4510 => x"8a",
          4511 => x"70",
          4512 => x"06",
          4513 => x"ff",
          4514 => x"38",
          4515 => x"16",
          4516 => x"80",
          4517 => x"75",
          4518 => x"f8",
          4519 => x"f7",
          4520 => x"c8",
          4521 => x"81",
          4522 => x"88",
          4523 => x"26",
          4524 => x"39",
          4525 => x"86",
          4526 => x"82",
          4527 => x"ff",
          4528 => x"38",
          4529 => x"05",
          4530 => x"76",
          4531 => x"55",
          4532 => x"81",
          4533 => x"3d",
          4534 => x"bc",
          4535 => x"74",
          4536 => x"6b",
          4537 => x"56",
          4538 => x"26",
          4539 => x"89",
          4540 => x"86",
          4541 => x"e5",
          4542 => x"38",
          4543 => x"a8",
          4544 => x"05",
          4545 => x"70",
          4546 => x"56",
          4547 => x"2e",
          4548 => x"94",
          4549 => x"57",
          4550 => x"8c",
          4551 => x"70",
          4552 => x"73",
          4553 => x"38",
          4554 => x"41",
          4555 => x"3d",
          4556 => x"ff",
          4557 => x"91",
          4558 => x"54",
          4559 => x"08",
          4560 => x"81",
          4561 => x"ff",
          4562 => x"91",
          4563 => x"54",
          4564 => x"08",
          4565 => x"80",
          4566 => x"8b",
          4567 => x"ff",
          4568 => x"65",
          4569 => x"c0",
          4570 => x"65",
          4571 => x"34",
          4572 => x"0b",
          4573 => x"77",
          4574 => x"92",
          4575 => x"c8",
          4576 => x"df",
          4577 => x"c8",
          4578 => x"09",
          4579 => x"d3",
          4580 => x"76",
          4581 => x"cb",
          4582 => x"9a",
          4583 => x"51",
          4584 => x"3f",
          4585 => x"08",
          4586 => x"c8",
          4587 => x"a0",
          4588 => x"c8",
          4589 => x"51",
          4590 => x"3f",
          4591 => x"0b",
          4592 => x"8b",
          4593 => x"ff",
          4594 => x"65",
          4595 => x"d8",
          4596 => x"81",
          4597 => x"34",
          4598 => x"a6",
          4599 => x"d3",
          4600 => x"73",
          4601 => x"d3",
          4602 => x"3d",
          4603 => x"3d",
          4604 => x"02",
          4605 => x"cf",
          4606 => x"3d",
          4607 => x"72",
          4608 => x"58",
          4609 => x"91",
          4610 => x"57",
          4611 => x"08",
          4612 => x"18",
          4613 => x"80",
          4614 => x"76",
          4615 => x"39",
          4616 => x"95",
          4617 => x"08",
          4618 => x"18",
          4619 => x"2a",
          4620 => x"51",
          4621 => x"90",
          4622 => x"82",
          4623 => x"57",
          4624 => x"81",
          4625 => x"39",
          4626 => x"22",
          4627 => x"70",
          4628 => x"58",
          4629 => x"f9",
          4630 => x"16",
          4631 => x"30",
          4632 => x"9f",
          4633 => x"c8",
          4634 => x"8c",
          4635 => x"52",
          4636 => x"80",
          4637 => x"27",
          4638 => x"14",
          4639 => x"83",
          4640 => x"78",
          4641 => x"80",
          4642 => x"77",
          4643 => x"d7",
          4644 => x"c8",
          4645 => x"61",
          4646 => x"98",
          4647 => x"26",
          4648 => x"55",
          4649 => x"ff",
          4650 => x"ff",
          4651 => x"38",
          4652 => x"81",
          4653 => x"7e",
          4654 => x"85",
          4655 => x"80",
          4656 => x"2e",
          4657 => x"c1",
          4658 => x"76",
          4659 => x"7b",
          4660 => x"38",
          4661 => x"55",
          4662 => x"b3",
          4663 => x"54",
          4664 => x"09",
          4665 => x"38",
          4666 => x"53",
          4667 => x"51",
          4668 => x"3f",
          4669 => x"08",
          4670 => x"c8",
          4671 => x"74",
          4672 => x"18",
          4673 => x"75",
          4674 => x"39",
          4675 => x"76",
          4676 => x"7f",
          4677 => x"0c",
          4678 => x"2e",
          4679 => x"88",
          4680 => x"8c",
          4681 => x"18",
          4682 => x"07",
          4683 => x"19",
          4684 => x"11",
          4685 => x"55",
          4686 => x"08",
          4687 => x"38",
          4688 => x"7e",
          4689 => x"0c",
          4690 => x"33",
          4691 => x"55",
          4692 => x"34",
          4693 => x"91",
          4694 => x"91",
          4695 => x"ea",
          4696 => x"02",
          4697 => x"e7",
          4698 => x"3d",
          4699 => x"ff",
          4700 => x"91",
          4701 => x"56",
          4702 => x"0b",
          4703 => x"08",
          4704 => x"38",
          4705 => x"08",
          4706 => x"d3",
          4707 => x"74",
          4708 => x"87",
          4709 => x"55",
          4710 => x"75",
          4711 => x"5a",
          4712 => x"51",
          4713 => x"3f",
          4714 => x"08",
          4715 => x"70",
          4716 => x"56",
          4717 => x"8c",
          4718 => x"82",
          4719 => x"06",
          4720 => x"57",
          4721 => x"38",
          4722 => x"05",
          4723 => x"79",
          4724 => x"dd",
          4725 => x"c8",
          4726 => x"66",
          4727 => x"38",
          4728 => x"80",
          4729 => x"66",
          4730 => x"06",
          4731 => x"2e",
          4732 => x"47",
          4733 => x"77",
          4734 => x"38",
          4735 => x"92",
          4736 => x"80",
          4737 => x"38",
          4738 => x"06",
          4739 => x"2e",
          4740 => x"57",
          4741 => x"7d",
          4742 => x"fe",
          4743 => x"91",
          4744 => x"6c",
          4745 => x"53",
          4746 => x"f6",
          4747 => x"d3",
          4748 => x"91",
          4749 => x"29",
          4750 => x"62",
          4751 => x"91",
          4752 => x"30",
          4753 => x"c8",
          4754 => x"25",
          4755 => x"59",
          4756 => x"41",
          4757 => x"8a",
          4758 => x"3d",
          4759 => x"81",
          4760 => x"ff",
          4761 => x"81",
          4762 => x"c8",
          4763 => x"38",
          4764 => x"70",
          4765 => x"55",
          4766 => x"64",
          4767 => x"06",
          4768 => x"44",
          4769 => x"66",
          4770 => x"38",
          4771 => x"46",
          4772 => x"ff",
          4773 => x"bc",
          4774 => x"77",
          4775 => x"8a",
          4776 => x"81",
          4777 => x"06",
          4778 => x"80",
          4779 => x"7c",
          4780 => x"74",
          4781 => x"38",
          4782 => x"55",
          4783 => x"83",
          4784 => x"7c",
          4785 => x"93",
          4786 => x"74",
          4787 => x"84",
          4788 => x"61",
          4789 => x"81",
          4790 => x"38",
          4791 => x"65",
          4792 => x"5c",
          4793 => x"91",
          4794 => x"71",
          4795 => x"56",
          4796 => x"2e",
          4797 => x"77",
          4798 => x"81",
          4799 => x"71",
          4800 => x"22",
          4801 => x"5b",
          4802 => x"86",
          4803 => x"27",
          4804 => x"52",
          4805 => x"f4",
          4806 => x"d3",
          4807 => x"d3",
          4808 => x"10",
          4809 => x"87",
          4810 => x"fe",
          4811 => x"91",
          4812 => x"5c",
          4813 => x"0b",
          4814 => x"17",
          4815 => x"ff",
          4816 => x"27",
          4817 => x"8e",
          4818 => x"39",
          4819 => x"65",
          4820 => x"5c",
          4821 => x"91",
          4822 => x"71",
          4823 => x"56",
          4824 => x"2e",
          4825 => x"77",
          4826 => x"81",
          4827 => x"71",
          4828 => x"22",
          4829 => x"5b",
          4830 => x"86",
          4831 => x"27",
          4832 => x"52",
          4833 => x"f3",
          4834 => x"d3",
          4835 => x"84",
          4836 => x"d3",
          4837 => x"f5",
          4838 => x"81",
          4839 => x"c8",
          4840 => x"11",
          4841 => x"83",
          4842 => x"42",
          4843 => x"1e",
          4844 => x"fe",
          4845 => x"91",
          4846 => x"5c",
          4847 => x"5b",
          4848 => x"51",
          4849 => x"3f",
          4850 => x"08",
          4851 => x"06",
          4852 => x"7c",
          4853 => x"68",
          4854 => x"69",
          4855 => x"06",
          4856 => x"58",
          4857 => x"61",
          4858 => x"81",
          4859 => x"76",
          4860 => x"41",
          4861 => x"76",
          4862 => x"90",
          4863 => x"65",
          4864 => x"74",
          4865 => x"be",
          4866 => x"31",
          4867 => x"53",
          4868 => x"52",
          4869 => x"9e",
          4870 => x"c8",
          4871 => x"83",
          4872 => x"06",
          4873 => x"d3",
          4874 => x"ff",
          4875 => x"38",
          4876 => x"78",
          4877 => x"77",
          4878 => x"8e",
          4879 => x"39",
          4880 => x"09",
          4881 => x"d3",
          4882 => x"f5",
          4883 => x"38",
          4884 => x"78",
          4885 => x"80",
          4886 => x"38",
          4887 => x"f1",
          4888 => x"2a",
          4889 => x"74",
          4890 => x"38",
          4891 => x"e1",
          4892 => x"38",
          4893 => x"81",
          4894 => x"fc",
          4895 => x"57",
          4896 => x"75",
          4897 => x"93",
          4898 => x"38",
          4899 => x"81",
          4900 => x"fc",
          4901 => x"57",
          4902 => x"80",
          4903 => x"2e",
          4904 => x"83",
          4905 => x"75",
          4906 => x"75",
          4907 => x"57",
          4908 => x"38",
          4909 => x"52",
          4910 => x"9a",
          4911 => x"53",
          4912 => x"52",
          4913 => x"99",
          4914 => x"52",
          4915 => x"ff",
          4916 => x"78",
          4917 => x"34",
          4918 => x"ff",
          4919 => x"1f",
          4920 => x"f7",
          4921 => x"90",
          4922 => x"83",
          4923 => x"70",
          4924 => x"80",
          4925 => x"55",
          4926 => x"ff",
          4927 => x"65",
          4928 => x"26",
          4929 => x"80",
          4930 => x"52",
          4931 => x"ff",
          4932 => x"8a",
          4933 => x"a0",
          4934 => x"98",
          4935 => x"7f",
          4936 => x"bf",
          4937 => x"51",
          4938 => x"3f",
          4939 => x"9a",
          4940 => x"98",
          4941 => x"52",
          4942 => x"ff",
          4943 => x"61",
          4944 => x"81",
          4945 => x"38",
          4946 => x"0a",
          4947 => x"1f",
          4948 => x"a5",
          4949 => x"a4",
          4950 => x"98",
          4951 => x"52",
          4952 => x"ff",
          4953 => x"81",
          4954 => x"51",
          4955 => x"3f",
          4956 => x"1f",
          4957 => x"e3",
          4958 => x"7f",
          4959 => x"34",
          4960 => x"c2",
          4961 => x"53",
          4962 => x"52",
          4963 => x"51",
          4964 => x"3f",
          4965 => x"88",
          4966 => x"a7",
          4967 => x"97",
          4968 => x"83",
          4969 => x"52",
          4970 => x"ff",
          4971 => x"ff",
          4972 => x"05",
          4973 => x"a6",
          4974 => x"53",
          4975 => x"52",
          4976 => x"ff",
          4977 => x"82",
          4978 => x"83",
          4979 => x"ff",
          4980 => x"81",
          4981 => x"7e",
          4982 => x"ff",
          4983 => x"81",
          4984 => x"c8",
          4985 => x"38",
          4986 => x"09",
          4987 => x"f0",
          4988 => x"63",
          4989 => x"7e",
          4990 => x"ff",
          4991 => x"7d",
          4992 => x"7e",
          4993 => x"c4",
          4994 => x"85",
          4995 => x"7e",
          4996 => x"e5",
          4997 => x"85",
          4998 => x"83",
          4999 => x"ff",
          5000 => x"ff",
          5001 => x"e8",
          5002 => x"96",
          5003 => x"52",
          5004 => x"51",
          5005 => x"3f",
          5006 => x"52",
          5007 => x"51",
          5008 => x"3f",
          5009 => x"87",
          5010 => x"52",
          5011 => x"93",
          5012 => x"54",
          5013 => x"53",
          5014 => x"51",
          5015 => x"3f",
          5016 => x"52",
          5017 => x"96",
          5018 => x"56",
          5019 => x"83",
          5020 => x"06",
          5021 => x"52",
          5022 => x"95",
          5023 => x"52",
          5024 => x"ff",
          5025 => x"f0",
          5026 => x"1f",
          5027 => x"e9",
          5028 => x"87",
          5029 => x"55",
          5030 => x"83",
          5031 => x"74",
          5032 => x"ff",
          5033 => x"7b",
          5034 => x"74",
          5035 => x"38",
          5036 => x"54",
          5037 => x"52",
          5038 => x"92",
          5039 => x"d3",
          5040 => x"86",
          5041 => x"80",
          5042 => x"ff",
          5043 => x"76",
          5044 => x"31",
          5045 => x"d1",
          5046 => x"5b",
          5047 => x"ff",
          5048 => x"55",
          5049 => x"83",
          5050 => x"60",
          5051 => x"26",
          5052 => x"57",
          5053 => x"53",
          5054 => x"51",
          5055 => x"3f",
          5056 => x"08",
          5057 => x"76",
          5058 => x"31",
          5059 => x"db",
          5060 => x"61",
          5061 => x"38",
          5062 => x"83",
          5063 => x"8a",
          5064 => x"61",
          5065 => x"38",
          5066 => x"83",
          5067 => x"58",
          5068 => x"38",
          5069 => x"52",
          5070 => x"95",
          5071 => x"d4",
          5072 => x"fe",
          5073 => x"94",
          5074 => x"be",
          5075 => x"76",
          5076 => x"81",
          5077 => x"0b",
          5078 => x"77",
          5079 => x"76",
          5080 => x"63",
          5081 => x"80",
          5082 => x"76",
          5083 => x"c6",
          5084 => x"85",
          5085 => x"d3",
          5086 => x"2a",
          5087 => x"74",
          5088 => x"91",
          5089 => x"87",
          5090 => x"52",
          5091 => x"51",
          5092 => x"3f",
          5093 => x"ca",
          5094 => x"93",
          5095 => x"54",
          5096 => x"52",
          5097 => x"90",
          5098 => x"57",
          5099 => x"08",
          5100 => x"53",
          5101 => x"51",
          5102 => x"3f",
          5103 => x"d3",
          5104 => x"38",
          5105 => x"57",
          5106 => x"57",
          5107 => x"57",
          5108 => x"57",
          5109 => x"c8",
          5110 => x"0d",
          5111 => x"0d",
          5112 => x"93",
          5113 => x"38",
          5114 => x"91",
          5115 => x"52",
          5116 => x"91",
          5117 => x"ff",
          5118 => x"81",
          5119 => x"c2",
          5120 => x"80",
          5121 => x"c9",
          5122 => x"98",
          5123 => x"93",
          5124 => x"39",
          5125 => x"51",
          5126 => x"3f",
          5127 => x"91",
          5128 => x"fe",
          5129 => x"81",
          5130 => x"c2",
          5131 => x"ff",
          5132 => x"9d",
          5133 => x"e0",
          5134 => x"e7",
          5135 => x"39",
          5136 => x"51",
          5137 => x"3f",
          5138 => x"91",
          5139 => x"fe",
          5140 => x"80",
          5141 => x"c3",
          5142 => x"ff",
          5143 => x"f1",
          5144 => x"b8",
          5145 => x"bb",
          5146 => x"39",
          5147 => x"51",
          5148 => x"3f",
          5149 => x"91",
          5150 => x"fe",
          5151 => x"80",
          5152 => x"c4",
          5153 => x"ff",
          5154 => x"c5",
          5155 => x"a8",
          5156 => x"8f",
          5157 => x"91",
          5158 => x"fe",
          5159 => x"b1",
          5160 => x"dc",
          5161 => x"fb",
          5162 => x"91",
          5163 => x"fe",
          5164 => x"9d",
          5165 => x"8c",
          5166 => x"e7",
          5167 => x"91",
          5168 => x"fe",
          5169 => x"89",
          5170 => x"b0",
          5171 => x"d3",
          5172 => x"0d",
          5173 => x"0d",
          5174 => x"56",
          5175 => x"26",
          5176 => x"52",
          5177 => x"29",
          5178 => x"ca",
          5179 => x"c8",
          5180 => x"39",
          5181 => x"74",
          5182 => x"ba",
          5183 => x"c8",
          5184 => x"51",
          5185 => x"3f",
          5186 => x"08",
          5187 => x"79",
          5188 => x"91",
          5189 => x"ff",
          5190 => x"87",
          5191 => x"fe",
          5192 => x"81",
          5193 => x"81",
          5194 => x"02",
          5195 => x"e3",
          5196 => x"73",
          5197 => x"07",
          5198 => x"ff",
          5199 => x"54",
          5200 => x"57",
          5201 => x"75",
          5202 => x"81",
          5203 => x"81",
          5204 => x"d8",
          5205 => x"bc",
          5206 => x"d3",
          5207 => x"91",
          5208 => x"bb",
          5209 => x"c8",
          5210 => x"98",
          5211 => x"d3",
          5212 => x"81",
          5213 => x"d4",
          5214 => x"84",
          5215 => x"52",
          5216 => x"51",
          5217 => x"91",
          5218 => x"58",
          5219 => x"08",
          5220 => x"80",
          5221 => x"7a",
          5222 => x"58",
          5223 => x"81",
          5224 => x"d8",
          5225 => x"c1",
          5226 => x"70",
          5227 => x"25",
          5228 => x"9f",
          5229 => x"51",
          5230 => x"74",
          5231 => x"38",
          5232 => x"53",
          5233 => x"88",
          5234 => x"51",
          5235 => x"77",
          5236 => x"d3",
          5237 => x"96",
          5238 => x"f8",
          5239 => x"b7",
          5240 => x"ff",
          5241 => x"80",
          5242 => x"7a",
          5243 => x"3f",
          5244 => x"08",
          5245 => x"80",
          5246 => x"76",
          5247 => x"38",
          5248 => x"55",
          5249 => x"d3",
          5250 => x"52",
          5251 => x"2d",
          5252 => x"08",
          5253 => x"75",
          5254 => x"d3",
          5255 => x"3d",
          5256 => x"3d",
          5257 => x"05",
          5258 => x"ec",
          5259 => x"f4",
          5260 => x"81",
          5261 => x"cb",
          5262 => x"52",
          5263 => x"d6",
          5264 => x"80",
          5265 => x"8c",
          5266 => x"33",
          5267 => x"94",
          5268 => x"c9",
          5269 => x"2e",
          5270 => x"f6",
          5271 => x"3d",
          5272 => x"3d",
          5273 => x"96",
          5274 => x"fe",
          5275 => x"81",
          5276 => x"ff",
          5277 => x"b0",
          5278 => x"f5",
          5279 => x"fe",
          5280 => x"72",
          5281 => x"81",
          5282 => x"71",
          5283 => x"38",
          5284 => x"ee",
          5285 => x"c6",
          5286 => x"f0",
          5287 => x"51",
          5288 => x"3f",
          5289 => x"70",
          5290 => x"52",
          5291 => x"95",
          5292 => x"fe",
          5293 => x"91",
          5294 => x"fe",
          5295 => x"80",
          5296 => x"af",
          5297 => x"2a",
          5298 => x"51",
          5299 => x"2e",
          5300 => x"51",
          5301 => x"3f",
          5302 => x"51",
          5303 => x"3f",
          5304 => x"ee",
          5305 => x"84",
          5306 => x"06",
          5307 => x"80",
          5308 => x"81",
          5309 => x"fb",
          5310 => x"84",
          5311 => x"f1",
          5312 => x"fe",
          5313 => x"72",
          5314 => x"81",
          5315 => x"71",
          5316 => x"38",
          5317 => x"ed",
          5318 => x"c7",
          5319 => x"ef",
          5320 => x"51",
          5321 => x"3f",
          5322 => x"70",
          5323 => x"52",
          5324 => x"95",
          5325 => x"fe",
          5326 => x"91",
          5327 => x"fe",
          5328 => x"80",
          5329 => x"ab",
          5330 => x"2a",
          5331 => x"51",
          5332 => x"2e",
          5333 => x"51",
          5334 => x"3f",
          5335 => x"51",
          5336 => x"3f",
          5337 => x"ed",
          5338 => x"88",
          5339 => x"06",
          5340 => x"80",
          5341 => x"81",
          5342 => x"f7",
          5343 => x"d4",
          5344 => x"ed",
          5345 => x"fe",
          5346 => x"fe",
          5347 => x"84",
          5348 => x"fa",
          5349 => x"70",
          5350 => x"56",
          5351 => x"2e",
          5352 => x"8e",
          5353 => x"0c",
          5354 => x"53",
          5355 => x"81",
          5356 => x"75",
          5357 => x"72",
          5358 => x"38",
          5359 => x"30",
          5360 => x"75",
          5361 => x"72",
          5362 => x"33",
          5363 => x"2e",
          5364 => x"88",
          5365 => x"70",
          5366 => x"34",
          5367 => x"90",
          5368 => x"88",
          5369 => x"53",
          5370 => x"54",
          5371 => x"3f",
          5372 => x"08",
          5373 => x"14",
          5374 => x"81",
          5375 => x"38",
          5376 => x"81",
          5377 => x"53",
          5378 => x"d2",
          5379 => x"72",
          5380 => x"0c",
          5381 => x"04",
          5382 => x"80",
          5383 => x"c8",
          5384 => x"5d",
          5385 => x"5a",
          5386 => x"51",
          5387 => x"3f",
          5388 => x"08",
          5389 => x"59",
          5390 => x"09",
          5391 => x"38",
          5392 => x"52",
          5393 => x"52",
          5394 => x"e7",
          5395 => x"78",
          5396 => x"1b",
          5397 => x"ab",
          5398 => x"c8",
          5399 => x"80",
          5400 => x"91",
          5401 => x"fe",
          5402 => x"85",
          5403 => x"5e",
          5404 => x"d0",
          5405 => x"ab",
          5406 => x"70",
          5407 => x"f8",
          5408 => x"80",
          5409 => x"fe",
          5410 => x"79",
          5411 => x"fe",
          5412 => x"b4",
          5413 => x"05",
          5414 => x"3f",
          5415 => x"08",
          5416 => x"90",
          5417 => x"78",
          5418 => x"85",
          5419 => x"10",
          5420 => x"88",
          5421 => x"08",
          5422 => x"fe",
          5423 => x"fe",
          5424 => x"fe",
          5425 => x"91",
          5426 => x"8c",
          5427 => x"d4",
          5428 => x"c9",
          5429 => x"39",
          5430 => x"f0",
          5431 => x"f8",
          5432 => x"fe",
          5433 => x"d3",
          5434 => x"2e",
          5435 => x"60",
          5436 => x"80",
          5437 => x"05",
          5438 => x"80",
          5439 => x"51",
          5440 => x"3f",
          5441 => x"08",
          5442 => x"59",
          5443 => x"91",
          5444 => x"fe",
          5445 => x"81",
          5446 => x"39",
          5447 => x"51",
          5448 => x"3f",
          5449 => x"b4",
          5450 => x"11",
          5451 => x"05",
          5452 => x"f4",
          5453 => x"c8",
          5454 => x"fe",
          5455 => x"53",
          5456 => x"80",
          5457 => x"51",
          5458 => x"3f",
          5459 => x"08",
          5460 => x"8c",
          5461 => x"c5",
          5462 => x"39",
          5463 => x"f4",
          5464 => x"f8",
          5465 => x"fd",
          5466 => x"d3",
          5467 => x"2e",
          5468 => x"89",
          5469 => x"38",
          5470 => x"f0",
          5471 => x"f8",
          5472 => x"fd",
          5473 => x"d3",
          5474 => x"38",
          5475 => x"08",
          5476 => x"91",
          5477 => x"96",
          5478 => x"59",
          5479 => x"3f",
          5480 => x"33",
          5481 => x"60",
          5482 => x"91",
          5483 => x"51",
          5484 => x"3f",
          5485 => x"08",
          5486 => x"38",
          5487 => x"08",
          5488 => x"3f",
          5489 => x"91",
          5490 => x"fe",
          5491 => x"81",
          5492 => x"39",
          5493 => x"f8",
          5494 => x"e4",
          5495 => x"d3",
          5496 => x"3d",
          5497 => x"52",
          5498 => x"fa",
          5499 => x"91",
          5500 => x"52",
          5501 => x"a7",
          5502 => x"c8",
          5503 => x"fc",
          5504 => x"d3",
          5505 => x"f3",
          5506 => x"e5",
          5507 => x"fe",
          5508 => x"fe",
          5509 => x"91",
          5510 => x"b5",
          5511 => x"05",
          5512 => x"e4",
          5513 => x"d3",
          5514 => x"3d",
          5515 => x"52",
          5516 => x"b2",
          5517 => x"c8",
          5518 => x"fe",
          5519 => x"59",
          5520 => x"3f",
          5521 => x"58",
          5522 => x"57",
          5523 => x"55",
          5524 => x"08",
          5525 => x"54",
          5526 => x"52",
          5527 => x"fb",
          5528 => x"c8",
          5529 => x"fc",
          5530 => x"d3",
          5531 => x"f2",
          5532 => x"fd",
          5533 => x"98",
          5534 => x"a7",
          5535 => x"fe",
          5536 => x"fb",
          5537 => x"c9",
          5538 => x"f3",
          5539 => x"51",
          5540 => x"3f",
          5541 => x"84",
          5542 => x"87",
          5543 => x"0c",
          5544 => x"0b",
          5545 => x"94",
          5546 => x"c8",
          5547 => x"f3",
          5548 => x"39",
          5549 => x"51",
          5550 => x"3f",
          5551 => x"0b",
          5552 => x"84",
          5553 => x"83",
          5554 => x"94",
          5555 => x"a1",
          5556 => x"fe",
          5557 => x"fe",
          5558 => x"fe",
          5559 => x"91",
          5560 => x"80",
          5561 => x"38",
          5562 => x"c9",
          5563 => x"f8",
          5564 => x"59",
          5565 => x"3d",
          5566 => x"53",
          5567 => x"51",
          5568 => x"3f",
          5569 => x"08",
          5570 => x"e5",
          5571 => x"91",
          5572 => x"fe",
          5573 => x"60",
          5574 => x"91",
          5575 => x"5e",
          5576 => x"08",
          5577 => x"c9",
          5578 => x"c8",
          5579 => x"ca",
          5580 => x"f7",
          5581 => x"b9",
          5582 => x"c4",
          5583 => x"e3",
          5584 => x"bc",
          5585 => x"39",
          5586 => x"51",
          5587 => x"3f",
          5588 => x"a0",
          5589 => x"84",
          5590 => x"39",
          5591 => x"51",
          5592 => x"2e",
          5593 => x"7c",
          5594 => x"78",
          5595 => x"cb",
          5596 => x"fe",
          5597 => x"fe",
          5598 => x"91",
          5599 => x"91",
          5600 => x"55",
          5601 => x"54",
          5602 => x"ca",
          5603 => x"3d",
          5604 => x"fe",
          5605 => x"91",
          5606 => x"91",
          5607 => x"80",
          5608 => x"05",
          5609 => x"80",
          5610 => x"80",
          5611 => x"80",
          5612 => x"f4",
          5613 => x"d3",
          5614 => x"7c",
          5615 => x"81",
          5616 => x"78",
          5617 => x"ff",
          5618 => x"06",
          5619 => x"91",
          5620 => x"fe",
          5621 => x"f9",
          5622 => x"3d",
          5623 => x"91",
          5624 => x"9b",
          5625 => x"0b",
          5626 => x"8c",
          5627 => x"86",
          5628 => x"c0",
          5629 => x"8c",
          5630 => x"87",
          5631 => x"0c",
          5632 => x"0b",
          5633 => x"94",
          5634 => x"8d",
          5635 => x"d8",
          5636 => x"80",
          5637 => x"dc",
          5638 => x"87",
          5639 => x"cd",
          5640 => x"9c",
          5641 => x"c9",
          5642 => x"a8",
          5643 => x"f3",
          5644 => x"e2",
          5645 => x"b0",
          5646 => x"f3",
          5647 => x"d8",
          5648 => x"00",
          5649 => x"5d",
          5650 => x"30",
          5651 => x"39",
          5652 => x"42",
          5653 => x"4b",
          5654 => x"54",
          5655 => x"cf",
          5656 => x"c0",
          5657 => x"d7",
          5658 => x"df",
          5659 => x"df",
          5660 => x"df",
          5661 => x"df",
          5662 => x"df",
          5663 => x"df",
          5664 => x"df",
          5665 => x"df",
          5666 => x"df",
          5667 => x"df",
          5668 => x"d3",
          5669 => x"df",
          5670 => x"df",
          5671 => x"df",
          5672 => x"53",
          5673 => x"df",
          5674 => x"d7",
          5675 => x"df",
          5676 => x"df",
          5677 => x"db",
          5678 => x"bf",
          5679 => x"f3",
          5680 => x"fe",
          5681 => x"09",
          5682 => x"14",
          5683 => x"1f",
          5684 => x"2a",
          5685 => x"35",
          5686 => x"40",
          5687 => x"4b",
          5688 => x"56",
          5689 => x"61",
          5690 => x"6c",
          5691 => x"77",
          5692 => x"82",
          5693 => x"8d",
          5694 => x"97",
          5695 => x"a1",
          5696 => x"ab",
          5697 => x"b5",
          5698 => x"71",
          5699 => x"5c",
          5700 => x"b9",
          5701 => x"5c",
          5702 => x"27",
          5703 => x"5c",
          5704 => x"5c",
          5705 => x"5c",
          5706 => x"5c",
          5707 => x"5c",
          5708 => x"5c",
          5709 => x"5c",
          5710 => x"5c",
          5711 => x"5c",
          5712 => x"5c",
          5713 => x"5c",
          5714 => x"5c",
          5715 => x"5c",
          5716 => x"5c",
          5717 => x"5c",
          5718 => x"5c",
          5719 => x"5c",
          5720 => x"5c",
          5721 => x"5c",
          5722 => x"5c",
          5723 => x"5c",
          5724 => x"5c",
          5725 => x"5c",
          5726 => x"5c",
          5727 => x"5c",
          5728 => x"5c",
          5729 => x"5c",
          5730 => x"5c",
          5731 => x"5c",
          5732 => x"5c",
          5733 => x"5c",
          5734 => x"5c",
          5735 => x"5c",
          5736 => x"5c",
          5737 => x"5c",
          5738 => x"5c",
          5739 => x"5c",
          5740 => x"5c",
          5741 => x"d4",
          5742 => x"5c",
          5743 => x"5c",
          5744 => x"5c",
          5745 => x"5c",
          5746 => x"0d",
          5747 => x"5c",
          5748 => x"5c",
          5749 => x"5c",
          5750 => x"5c",
          5751 => x"5c",
          5752 => x"5c",
          5753 => x"5c",
          5754 => x"5c",
          5755 => x"5c",
          5756 => x"5c",
          5757 => x"5c",
          5758 => x"5c",
          5759 => x"5c",
          5760 => x"5c",
          5761 => x"5c",
          5762 => x"5c",
          5763 => x"5c",
          5764 => x"5c",
          5765 => x"5c",
          5766 => x"5c",
          5767 => x"5c",
          5768 => x"5c",
          5769 => x"5c",
          5770 => x"5c",
          5771 => x"5c",
          5772 => x"5c",
          5773 => x"5c",
          5774 => x"5c",
          5775 => x"5c",
          5776 => x"5c",
          5777 => x"5c",
          5778 => x"75",
          5779 => x"86",
          5780 => x"5c",
          5781 => x"5c",
          5782 => x"97",
          5783 => x"b4",
          5784 => x"5c",
          5785 => x"5c",
          5786 => x"5c",
          5787 => x"5c",
          5788 => x"5c",
          5789 => x"5c",
          5790 => x"5c",
          5791 => x"5c",
          5792 => x"5c",
          5793 => x"5c",
          5794 => x"5c",
          5795 => x"5c",
          5796 => x"5c",
          5797 => x"5c",
          5798 => x"5c",
          5799 => x"5c",
          5800 => x"5c",
          5801 => x"5c",
          5802 => x"5c",
          5803 => x"5c",
          5804 => x"5c",
          5805 => x"5c",
          5806 => x"5c",
          5807 => x"5c",
          5808 => x"5c",
          5809 => x"5c",
          5810 => x"5c",
          5811 => x"5c",
          5812 => x"5c",
          5813 => x"5c",
          5814 => x"5c",
          5815 => x"5c",
          5816 => x"5c",
          5817 => x"5c",
          5818 => x"d1",
          5819 => x"f6",
          5820 => x"5c",
          5821 => x"5c",
          5822 => x"5c",
          5823 => x"5c",
          5824 => x"5c",
          5825 => x"5c",
          5826 => x"5c",
          5827 => x"5c",
          5828 => x"39",
          5829 => x"48",
          5830 => x"5c",
          5831 => x"55",
          5832 => x"5c",
          5833 => x"71",
          5834 => x"25",
          5835 => x"64",
          5836 => x"3a",
          5837 => x"25",
          5838 => x"64",
          5839 => x"00",
          5840 => x"20",
          5841 => x"66",
          5842 => x"72",
          5843 => x"6f",
          5844 => x"00",
          5845 => x"72",
          5846 => x"53",
          5847 => x"63",
          5848 => x"69",
          5849 => x"00",
          5850 => x"65",
          5851 => x"65",
          5852 => x"6d",
          5853 => x"6d",
          5854 => x"65",
          5855 => x"00",
          5856 => x"20",
          5857 => x"4e",
          5858 => x"41",
          5859 => x"53",
          5860 => x"74",
          5861 => x"38",
          5862 => x"53",
          5863 => x"3d",
          5864 => x"58",
          5865 => x"00",
          5866 => x"20",
          5867 => x"4d",
          5868 => x"74",
          5869 => x"3d",
          5870 => x"58",
          5871 => x"69",
          5872 => x"25",
          5873 => x"29",
          5874 => x"00",
          5875 => x"20",
          5876 => x"20",
          5877 => x"61",
          5878 => x"25",
          5879 => x"2c",
          5880 => x"7a",
          5881 => x"30",
          5882 => x"2e",
          5883 => x"00",
          5884 => x"20",
          5885 => x"54",
          5886 => x"00",
          5887 => x"20",
          5888 => x"0a",
          5889 => x"00",
          5890 => x"20",
          5891 => x"0a",
          5892 => x"00",
          5893 => x"20",
          5894 => x"43",
          5895 => x"20",
          5896 => x"76",
          5897 => x"73",
          5898 => x"32",
          5899 => x"0a",
          5900 => x"00",
          5901 => x"20",
          5902 => x"45",
          5903 => x"50",
          5904 => x"4f",
          5905 => x"4f",
          5906 => x"52",
          5907 => x"00",
          5908 => x"20",
          5909 => x"45",
          5910 => x"28",
          5911 => x"65",
          5912 => x"25",
          5913 => x"29",
          5914 => x"00",
          5915 => x"72",
          5916 => x"65",
          5917 => x"00",
          5918 => x"20",
          5919 => x"20",
          5920 => x"65",
          5921 => x"65",
          5922 => x"72",
          5923 => x"64",
          5924 => x"73",
          5925 => x"25",
          5926 => x"0a",
          5927 => x"00",
          5928 => x"20",
          5929 => x"20",
          5930 => x"6f",
          5931 => x"53",
          5932 => x"74",
          5933 => x"64",
          5934 => x"73",
          5935 => x"25",
          5936 => x"0a",
          5937 => x"00",
          5938 => x"20",
          5939 => x"63",
          5940 => x"74",
          5941 => x"20",
          5942 => x"72",
          5943 => x"20",
          5944 => x"20",
          5945 => x"25",
          5946 => x"0a",
          5947 => x"00",
          5948 => x"20",
          5949 => x"20",
          5950 => x"20",
          5951 => x"20",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"25",
          5956 => x"0a",
          5957 => x"00",
          5958 => x"20",
          5959 => x"74",
          5960 => x"43",
          5961 => x"6b",
          5962 => x"65",
          5963 => x"20",
          5964 => x"20",
          5965 => x"25",
          5966 => x"0a",
          5967 => x"00",
          5968 => x"6c",
          5969 => x"00",
          5970 => x"69",
          5971 => x"00",
          5972 => x"78",
          5973 => x"00",
          5974 => x"00",
          5975 => x"6d",
          5976 => x"00",
          5977 => x"6e",
          5978 => x"00",
          5979 => x"00",
          5980 => x"2c",
          5981 => x"3d",
          5982 => x"5d",
          5983 => x"00",
          5984 => x"00",
          5985 => x"33",
          5986 => x"00",
          5987 => x"00",
          5988 => x"00",
          5989 => x"00",
          5990 => x"00",
          5991 => x"00",
          5992 => x"00",
          5993 => x"00",
          5994 => x"00",
          5995 => x"00",
          5996 => x"00",
          5997 => x"4d",
          5998 => x"53",
          5999 => x"00",
          6000 => x"4e",
          6001 => x"20",
          6002 => x"46",
          6003 => x"32",
          6004 => x"00",
          6005 => x"4e",
          6006 => x"20",
          6007 => x"46",
          6008 => x"20",
          6009 => x"00",
          6010 => x"6c",
          6011 => x"00",
          6012 => x"00",
          6013 => x"00",
          6014 => x"41",
          6015 => x"80",
          6016 => x"49",
          6017 => x"8f",
          6018 => x"4f",
          6019 => x"55",
          6020 => x"9b",
          6021 => x"9f",
          6022 => x"55",
          6023 => x"a7",
          6024 => x"ab",
          6025 => x"af",
          6026 => x"b3",
          6027 => x"b7",
          6028 => x"bb",
          6029 => x"bf",
          6030 => x"c3",
          6031 => x"c7",
          6032 => x"cb",
          6033 => x"cf",
          6034 => x"d3",
          6035 => x"d7",
          6036 => x"db",
          6037 => x"df",
          6038 => x"e3",
          6039 => x"e7",
          6040 => x"eb",
          6041 => x"ef",
          6042 => x"f3",
          6043 => x"f7",
          6044 => x"fb",
          6045 => x"ff",
          6046 => x"3b",
          6047 => x"2f",
          6048 => x"3a",
          6049 => x"7c",
          6050 => x"00",
          6051 => x"04",
          6052 => x"40",
          6053 => x"00",
          6054 => x"00",
          6055 => x"02",
          6056 => x"08",
          6057 => x"20",
          6058 => x"00",
          6059 => x"31",
          6060 => x"00",
          6061 => x"31",
          6062 => x"00",
          6063 => x"41",
          6064 => x"00",
          6065 => x"4b",
          6066 => x"20",
          6067 => x"54",
          6068 => x"53",
          6069 => x"00",
          6070 => x"4b",
          6071 => x"46",
          6072 => x"20",
          6073 => x"54",
          6074 => x"53",
          6075 => x"00",
          6076 => x"45",
          6077 => x"54",
          6078 => x"43",
          6079 => x"52",
          6080 => x"00",
          6081 => x"4f",
          6082 => x"00",
          6083 => x"44",
          6084 => x"45",
          6085 => x"00",
          6086 => x"54",
          6087 => x"00",
          6088 => x"43",
          6089 => x"4f",
          6090 => x"00",
          6091 => x"43",
          6092 => x"4d",
          6093 => x"44",
          6094 => x"00",
          6095 => x"6d",
          6096 => x"00",
          6097 => x"69",
          6098 => x"00",
          6099 => x"61",
          6100 => x"00",
          6101 => x"63",
          6102 => x"00",
          6103 => x"6d",
          6104 => x"00",
          6105 => x"69",
          6106 => x"00",
          6107 => x"61",
          6108 => x"00",
          6109 => x"69",
          6110 => x"00",
          6111 => x"6c",
          6112 => x"00",
          6113 => x"6e",
          6114 => x"00",
          6115 => x"69",
          6116 => x"00",
          6117 => x"65",
          6118 => x"00",
          6119 => x"6f",
          6120 => x"00",
          6121 => x"65",
          6122 => x"00",
          6123 => x"61",
          6124 => x"00",
          6125 => x"73",
          6126 => x"74",
          6127 => x"00",
          6128 => x"69",
          6129 => x"00",
          6130 => x"75",
          6131 => x"00",
          6132 => x"6c",
          6133 => x"00",
          6134 => x"74",
          6135 => x"00",
          6136 => x"6d",
          6137 => x"00",
          6138 => x"6e",
          6139 => x"00",
          6140 => x"6c",
          6141 => x"00",
          6142 => x"64",
          6143 => x"00",
          6144 => x"61",
          6145 => x"00",
          6146 => x"72",
          6147 => x"00",
          6148 => x"74",
          6149 => x"00",
          6150 => x"00",
          6151 => x"6e",
          6152 => x"00",
          6153 => x"72",
          6154 => x"00",
          6155 => x"61",
          6156 => x"00",
          6157 => x"65",
          6158 => x"00",
          6159 => x"76",
          6160 => x"00",
          6161 => x"6d",
          6162 => x"00",
          6163 => x"00",
          6164 => x"69",
          6165 => x"00",
          6166 => x"6f",
          6167 => x"72",
          6168 => x"00",
          6169 => x"62",
          6170 => x"00",
          6171 => x"66",
          6172 => x"00",
          6173 => x"72",
          6174 => x"00",
          6175 => x"6d",
          6176 => x"00",
          6177 => x"00",
          6178 => x"00",
          6179 => x"00",
          6180 => x"00",
          6181 => x"00",
          6182 => x"00",
          6183 => x"00",
          6184 => x"00",
          6185 => x"00",
          6186 => x"79",
          6187 => x"00",
          6188 => x"65",
          6189 => x"6b",
          6190 => x"00",
          6191 => x"6c",
          6192 => x"00",
          6193 => x"00",
          6194 => x"74",
          6195 => x"00",
          6196 => x"65",
          6197 => x"00",
          6198 => x"70",
          6199 => x"00",
          6200 => x"6f",
          6201 => x"00",
          6202 => x"65",
          6203 => x"00",
          6204 => x"74",
          6205 => x"00",
          6206 => x"6b",
          6207 => x"72",
          6208 => x"00",
          6209 => x"65",
          6210 => x"6c",
          6211 => x"72",
          6212 => x"0a",
          6213 => x"00",
          6214 => x"6b",
          6215 => x"74",
          6216 => x"61",
          6217 => x"0a",
          6218 => x"00",
          6219 => x"66",
          6220 => x"20",
          6221 => x"6e",
          6222 => x"00",
          6223 => x"70",
          6224 => x"20",
          6225 => x"6e",
          6226 => x"00",
          6227 => x"61",
          6228 => x"20",
          6229 => x"65",
          6230 => x"65",
          6231 => x"00",
          6232 => x"65",
          6233 => x"64",
          6234 => x"65",
          6235 => x"00",
          6236 => x"65",
          6237 => x"72",
          6238 => x"79",
          6239 => x"69",
          6240 => x"2e",
          6241 => x"00",
          6242 => x"65",
          6243 => x"6e",
          6244 => x"20",
          6245 => x"61",
          6246 => x"2e",
          6247 => x"00",
          6248 => x"69",
          6249 => x"72",
          6250 => x"20",
          6251 => x"74",
          6252 => x"65",
          6253 => x"00",
          6254 => x"76",
          6255 => x"75",
          6256 => x"72",
          6257 => x"20",
          6258 => x"61",
          6259 => x"2e",
          6260 => x"00",
          6261 => x"6b",
          6262 => x"74",
          6263 => x"61",
          6264 => x"64",
          6265 => x"00",
          6266 => x"63",
          6267 => x"61",
          6268 => x"6c",
          6269 => x"69",
          6270 => x"79",
          6271 => x"6d",
          6272 => x"75",
          6273 => x"6f",
          6274 => x"69",
          6275 => x"0a",
          6276 => x"00",
          6277 => x"6d",
          6278 => x"61",
          6279 => x"74",
          6280 => x"0a",
          6281 => x"00",
          6282 => x"65",
          6283 => x"2c",
          6284 => x"65",
          6285 => x"69",
          6286 => x"63",
          6287 => x"65",
          6288 => x"64",
          6289 => x"00",
          6290 => x"65",
          6291 => x"20",
          6292 => x"6b",
          6293 => x"0a",
          6294 => x"00",
          6295 => x"75",
          6296 => x"63",
          6297 => x"74",
          6298 => x"6d",
          6299 => x"2e",
          6300 => x"00",
          6301 => x"20",
          6302 => x"79",
          6303 => x"65",
          6304 => x"69",
          6305 => x"2e",
          6306 => x"00",
          6307 => x"61",
          6308 => x"65",
          6309 => x"69",
          6310 => x"72",
          6311 => x"74",
          6312 => x"00",
          6313 => x"63",
          6314 => x"2e",
          6315 => x"00",
          6316 => x"6e",
          6317 => x"20",
          6318 => x"6f",
          6319 => x"00",
          6320 => x"75",
          6321 => x"74",
          6322 => x"25",
          6323 => x"74",
          6324 => x"75",
          6325 => x"74",
          6326 => x"73",
          6327 => x"0a",
          6328 => x"00",
          6329 => x"64",
          6330 => x"00",
          6331 => x"54",
          6332 => x"00",
          6333 => x"20",
          6334 => x"28",
          6335 => x"00",
          6336 => x"30",
          6337 => x"30",
          6338 => x"00",
          6339 => x"33",
          6340 => x"00",
          6341 => x"55",
          6342 => x"65",
          6343 => x"30",
          6344 => x"20",
          6345 => x"25",
          6346 => x"2a",
          6347 => x"00",
          6348 => x"54",
          6349 => x"6e",
          6350 => x"72",
          6351 => x"20",
          6352 => x"64",
          6353 => x"0a",
          6354 => x"00",
          6355 => x"65",
          6356 => x"6e",
          6357 => x"72",
          6358 => x"0a",
          6359 => x"00",
          6360 => x"20",
          6361 => x"65",
          6362 => x"70",
          6363 => x"00",
          6364 => x"54",
          6365 => x"44",
          6366 => x"74",
          6367 => x"75",
          6368 => x"00",
          6369 => x"54",
          6370 => x"52",
          6371 => x"74",
          6372 => x"75",
          6373 => x"00",
          6374 => x"54",
          6375 => x"58",
          6376 => x"74",
          6377 => x"75",
          6378 => x"00",
          6379 => x"54",
          6380 => x"58",
          6381 => x"74",
          6382 => x"75",
          6383 => x"00",
          6384 => x"54",
          6385 => x"58",
          6386 => x"74",
          6387 => x"75",
          6388 => x"00",
          6389 => x"54",
          6390 => x"58",
          6391 => x"74",
          6392 => x"75",
          6393 => x"00",
          6394 => x"74",
          6395 => x"20",
          6396 => x"74",
          6397 => x"72",
          6398 => x"0a",
          6399 => x"00",
          6400 => x"62",
          6401 => x"67",
          6402 => x"6d",
          6403 => x"2e",
          6404 => x"00",
          6405 => x"00",
          6406 => x"6c",
          6407 => x"74",
          6408 => x"6e",
          6409 => x"61",
          6410 => x"65",
          6411 => x"20",
          6412 => x"64",
          6413 => x"20",
          6414 => x"61",
          6415 => x"69",
          6416 => x"20",
          6417 => x"75",
          6418 => x"79",
          6419 => x"00",
          6420 => x"00",
          6421 => x"20",
          6422 => x"6b",
          6423 => x"21",
          6424 => x"00",
          6425 => x"74",
          6426 => x"69",
          6427 => x"2e",
          6428 => x"00",
          6429 => x"6c",
          6430 => x"74",
          6431 => x"6e",
          6432 => x"61",
          6433 => x"65",
          6434 => x"00",
          6435 => x"25",
          6436 => x"00",
          6437 => x"00",
          6438 => x"61",
          6439 => x"6e",
          6440 => x"6e",
          6441 => x"72",
          6442 => x"73",
          6443 => x"00",
          6444 => x"62",
          6445 => x"67",
          6446 => x"74",
          6447 => x"75",
          6448 => x"0a",
          6449 => x"00",
          6450 => x"61",
          6451 => x"64",
          6452 => x"72",
          6453 => x"69",
          6454 => x"00",
          6455 => x"62",
          6456 => x"67",
          6457 => x"72",
          6458 => x"69",
          6459 => x"00",
          6460 => x"63",
          6461 => x"6e",
          6462 => x"6f",
          6463 => x"40",
          6464 => x"38",
          6465 => x"2e",
          6466 => x"00",
          6467 => x"6c",
          6468 => x"20",
          6469 => x"65",
          6470 => x"25",
          6471 => x"20",
          6472 => x"0a",
          6473 => x"00",
          6474 => x"6c",
          6475 => x"74",
          6476 => x"65",
          6477 => x"6f",
          6478 => x"28",
          6479 => x"2e",
          6480 => x"00",
          6481 => x"74",
          6482 => x"69",
          6483 => x"61",
          6484 => x"69",
          6485 => x"69",
          6486 => x"2e",
          6487 => x"00",
          6488 => x"64",
          6489 => x"62",
          6490 => x"69",
          6491 => x"2e",
          6492 => x"00",
          6493 => x"00",
          6494 => x"00",
          6495 => x"5c",
          6496 => x"25",
          6497 => x"73",
          6498 => x"00",
          6499 => x"20",
          6500 => x"6d",
          6501 => x"2e",
          6502 => x"00",
          6503 => x"6e",
          6504 => x"2e",
          6505 => x"00",
          6506 => x"62",
          6507 => x"67",
          6508 => x"74",
          6509 => x"75",
          6510 => x"2e",
          6511 => x"00",
          6512 => x"00",
          6513 => x"00",
          6514 => x"ff",
          6515 => x"00",
          6516 => x"ff",
          6517 => x"00",
          6518 => x"ff",
          6519 => x"00",
          6520 => x"00",
          6521 => x"00",
          6522 => x"00",
          6523 => x"00",
          6524 => x"01",
          6525 => x"01",
          6526 => x"01",
          6527 => x"00",
          6528 => x"00",
          6529 => x"00",
          6530 => x"3c",
          6531 => x"00",
          6532 => x"00",
          6533 => x"00",
          6534 => x"44",
          6535 => x"00",
          6536 => x"00",
          6537 => x"00",
          6538 => x"4c",
          6539 => x"00",
          6540 => x"00",
          6541 => x"00",
          6542 => x"54",
          6543 => x"00",
          6544 => x"00",
          6545 => x"00",
          6546 => x"5c",
          6547 => x"00",
          6548 => x"00",
          6549 => x"00",
          6550 => x"64",
          6551 => x"00",
          6552 => x"00",
          6553 => x"00",
          6554 => x"6c",
          6555 => x"00",
          6556 => x"00",
          6557 => x"00",
          6558 => x"74",
          6559 => x"00",
          6560 => x"00",
          6561 => x"00",
          6562 => x"7c",
          6563 => x"00",
          6564 => x"00",
          6565 => x"00",
          6566 => x"84",
          6567 => x"00",
          6568 => x"00",
          6569 => x"00",
          6570 => x"8c",
          6571 => x"00",
          6572 => x"00",
          6573 => x"00",
          6574 => x"94",
          6575 => x"00",
          6576 => x"00",
          6577 => x"00",
          6578 => x"9c",
          6579 => x"00",
          6580 => x"00",
          6581 => x"00",
          6582 => x"a4",
          6583 => x"00",
          6584 => x"00",
          6585 => x"00",
          6586 => x"ac",
          6587 => x"00",
          6588 => x"00",
          6589 => x"00",
          6590 => x"b4",
          6591 => x"00",
          6592 => x"00",
          6593 => x"00",
          6594 => x"c0",
          6595 => x"00",
          6596 => x"00",
          6597 => x"00",
          6598 => x"c8",
          6599 => x"00",
          6600 => x"00",
          6601 => x"00",
          6602 => x"d0",
          6603 => x"00",
          6604 => x"00",
          6605 => x"00",
          6606 => x"d8",
          6607 => x"00",
          6608 => x"00",
          6609 => x"00",
          6610 => x"e0",
          6611 => x"00",
          6612 => x"00",
          6613 => x"00",
          6614 => x"e8",
          6615 => x"00",
          6616 => x"00",
          6617 => x"00",
          6618 => x"f0",
          6619 => x"00",
          6620 => x"00",
          6621 => x"00",
          6622 => x"f8",
          6623 => x"00",
          6624 => x"00",
          6625 => x"00",
          6626 => x"00",
          6627 => x"00",
          6628 => x"00",
          6629 => x"00",
          6630 => x"08",
          6631 => x"00",
          6632 => x"00",
          6633 => x"00",
          6634 => x"10",
          6635 => x"00",
          6636 => x"00",
          6637 => x"00",
          6638 => x"18",
          6639 => x"00",
          6640 => x"00",
          6641 => x"00",
          6642 => x"1c",
          6643 => x"00",
          6644 => x"00",
          6645 => x"00",
          6646 => x"24",
          6647 => x"00",
          6648 => x"00",
          6649 => x"00",
          6650 => x"2c",
          6651 => x"00",
          6652 => x"00",
          6653 => x"00",
          6654 => x"34",
          6655 => x"00",
          6656 => x"00",
          6657 => x"00",
          6658 => x"3c",
          6659 => x"00",
          6660 => x"00",
          6661 => x"00",
          6662 => x"44",
          6663 => x"00",
          6664 => x"00",
          6665 => x"00",
          6666 => x"4c",
          6667 => x"00",
          6668 => x"00",
          6669 => x"00",
          6670 => x"50",
          6671 => x"00",
          6672 => x"00",
          6673 => x"00",
          6674 => x"58",
          6675 => x"00",
          6676 => x"00",
          6677 => x"00",
          6678 => x"64",
          6679 => x"00",
          6680 => x"00",
          6681 => x"00",
          6682 => x"6c",
          6683 => x"00",
          6684 => x"00",
          6685 => x"00",
          6686 => x"74",
          6687 => x"00",
          6688 => x"00",
          6689 => x"00",
          6690 => x"7c",
          6691 => x"00",
          6692 => x"00",
          6693 => x"00",
          6694 => x"84",
          6695 => x"00",
          6696 => x"00",
          6697 => x"00",
          6698 => x"88",
          6699 => x"00",
          6700 => x"00",
          6701 => x"00",
          6702 => x"8c",
          6703 => x"00",
          6704 => x"00",
          6705 => x"00",
          6706 => x"90",
          6707 => x"00",
          6708 => x"00",
          6709 => x"00",
          6710 => x"94",
          6711 => x"00",
          6712 => x"00",
          6713 => x"00",
          6714 => x"98",
          6715 => x"00",
          6716 => x"00",
          6717 => x"00",
          6718 => x"9c",
          6719 => x"00",
          6720 => x"00",
          6721 => x"00",
          6722 => x"a0",
          6723 => x"00",
          6724 => x"00",
          6725 => x"00",
          6726 => x"a4",
          6727 => x"00",
          6728 => x"00",
          6729 => x"00",
          6730 => x"a8",
          6731 => x"00",
          6732 => x"00",
          6733 => x"00",
          6734 => x"b0",
          6735 => x"00",
          6736 => x"00",
          6737 => x"00",
          6738 => x"bc",
          6739 => x"00",
          6740 => x"00",
          6741 => x"00",
          6742 => x"c4",
          6743 => x"00",
          6744 => x"00",
          6745 => x"00",
          6746 => x"c8",
          6747 => x"00",
          6748 => x"00",
          6749 => x"00",
          6750 => x"d0",
          6751 => x"00",
          6752 => x"00",
          6753 => x"00",
          6754 => x"d8",
          6755 => x"00",
          6756 => x"00",
          6757 => x"00",
          6758 => x"e0",
          6759 => x"00",
          6760 => x"00",
          6761 => x"00",
          6762 => x"e8",
          6763 => x"00",
          6764 => x"00",
          6765 => x"00",
          6766 => x"f0",
          6767 => x"00",
          6768 => x"00",
          6769 => x"00",
        others => X"00"
    );

    shared variable RAM1 : ramArray :=
    (
             0 => x"90",
             1 => x"0b",
             2 => x"95",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"90",
             9 => x"0b",
            10 => x"85",
            11 => x"90",
            12 => x"0b",
            13 => x"a5",
            14 => x"90",
            15 => x"0b",
            16 => x"c5",
            17 => x"90",
            18 => x"0b",
            19 => x"e5",
            20 => x"90",
            21 => x"0b",
            22 => x"85",
            23 => x"90",
            24 => x"0b",
            25 => x"a5",
            26 => x"90",
            27 => x"0b",
            28 => x"c5",
            29 => x"90",
            30 => x"0b",
            31 => x"e5",
            32 => x"90",
            33 => x"0b",
            34 => x"85",
            35 => x"90",
            36 => x"0b",
            37 => x"a5",
            38 => x"90",
            39 => x"0b",
            40 => x"c5",
            41 => x"90",
            42 => x"0b",
            43 => x"e5",
            44 => x"90",
            45 => x"0b",
            46 => x"85",
            47 => x"90",
            48 => x"0b",
            49 => x"a5",
            50 => x"90",
            51 => x"0b",
            52 => x"c5",
            53 => x"90",
            54 => x"0b",
            55 => x"e5",
            56 => x"90",
            57 => x"0b",
            58 => x"85",
            59 => x"90",
            60 => x"0b",
            61 => x"a5",
            62 => x"90",
            63 => x"0b",
            64 => x"c5",
            65 => x"90",
            66 => x"0b",
            67 => x"e5",
            68 => x"90",
            69 => x"0b",
            70 => x"85",
            71 => x"90",
            72 => x"0b",
            73 => x"a5",
            74 => x"90",
            75 => x"0b",
            76 => x"c5",
            77 => x"90",
            78 => x"0b",
            79 => x"e5",
            80 => x"90",
            81 => x"0b",
            82 => x"85",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"84",
           129 => x"d3",
           130 => x"95",
           131 => x"d3",
           132 => x"80",
           133 => x"d3",
           134 => x"9f",
           135 => x"d3",
           136 => x"80",
           137 => x"d3",
           138 => x"a0",
           139 => x"d3",
           140 => x"80",
           141 => x"d3",
           142 => x"a0",
           143 => x"d3",
           144 => x"80",
           145 => x"d3",
           146 => x"a6",
           147 => x"d3",
           148 => x"80",
           149 => x"d3",
           150 => x"a8",
           151 => x"d3",
           152 => x"80",
           153 => x"d3",
           154 => x"a0",
           155 => x"d3",
           156 => x"80",
           157 => x"d3",
           158 => x"a8",
           159 => x"d3",
           160 => x"80",
           161 => x"d3",
           162 => x"aa",
           163 => x"d3",
           164 => x"80",
           165 => x"d3",
           166 => x"a6",
           167 => x"d3",
           168 => x"80",
           169 => x"d3",
           170 => x"a6",
           171 => x"d3",
           172 => x"80",
           173 => x"d3",
           174 => x"a6",
           175 => x"d3",
           176 => x"80",
           177 => x"d3",
           178 => x"97",
           179 => x"d3",
           180 => x"80",
           181 => x"d3",
           182 => x"97",
           183 => x"d3",
           184 => x"80",
           185 => x"d3",
           186 => x"8f",
           187 => x"d3",
           188 => x"80",
           189 => x"d3",
           190 => x"91",
           191 => x"d3",
           192 => x"80",
           193 => x"d3",
           194 => x"92",
           195 => x"d3",
           196 => x"80",
           197 => x"d3",
           198 => x"de",
           199 => x"d3",
           200 => x"80",
           201 => x"d3",
           202 => x"ed",
           203 => x"d3",
           204 => x"80",
           205 => x"d3",
           206 => x"e3",
           207 => x"d3",
           208 => x"80",
           209 => x"d3",
           210 => x"e7",
           211 => x"d3",
           212 => x"80",
           213 => x"d3",
           214 => x"f3",
           215 => x"d3",
           216 => x"80",
           217 => x"d3",
           218 => x"fd",
           219 => x"d3",
           220 => x"80",
           221 => x"d3",
           222 => x"ec",
           223 => x"d3",
           224 => x"80",
           225 => x"d3",
           226 => x"f7",
           227 => x"d3",
           228 => x"80",
           229 => x"d3",
           230 => x"f8",
           231 => x"d3",
           232 => x"80",
           233 => x"d3",
           234 => x"f9",
           235 => x"d3",
           236 => x"80",
           237 => x"d3",
           238 => x"82",
           239 => x"d3",
           240 => x"80",
           241 => x"d3",
           242 => x"ff",
           243 => x"d3",
           244 => x"80",
           245 => x"d3",
           246 => x"84",
           247 => x"d3",
           248 => x"80",
           249 => x"d3",
           250 => x"fa",
           251 => x"d3",
           252 => x"80",
           253 => x"d3",
           254 => x"87",
           255 => x"d3",
           256 => x"80",
           257 => x"d3",
           258 => x"88",
           259 => x"d3",
           260 => x"80",
           261 => x"d3",
           262 => x"ee",
           263 => x"d3",
           264 => x"80",
           265 => x"d3",
           266 => x"ee",
           267 => x"d3",
           268 => x"80",
           269 => x"d3",
           270 => x"ef",
           271 => x"d3",
           272 => x"80",
           273 => x"d3",
           274 => x"fa",
           275 => x"d3",
           276 => x"80",
           277 => x"d3",
           278 => x"89",
           279 => x"d3",
           280 => x"80",
           281 => x"d3",
           282 => x"8c",
           283 => x"d3",
           284 => x"80",
           285 => x"d3",
           286 => x"8f",
           287 => x"d3",
           288 => x"80",
           289 => x"d3",
           290 => x"de",
           291 => x"d3",
           292 => x"80",
           293 => x"d3",
           294 => x"92",
           295 => x"d3",
           296 => x"80",
           297 => x"d3",
           298 => x"ad",
           299 => x"d3",
           300 => x"80",
           301 => x"d3",
           302 => x"af",
           303 => x"d3",
           304 => x"80",
           305 => x"d3",
           306 => x"b1",
           307 => x"d3",
           308 => x"80",
           309 => x"d3",
           310 => x"90",
           311 => x"d3",
           312 => x"80",
           313 => x"d3",
           314 => x"90",
           315 => x"d3",
           316 => x"80",
           317 => x"d3",
           318 => x"93",
           319 => x"d3",
           320 => x"80",
           321 => x"d3",
           322 => x"9f",
           323 => x"d3",
           324 => x"80",
           325 => x"d3",
           326 => x"f6",
           327 => x"38",
           328 => x"84",
           329 => x"0b",
           330 => x"98",
           331 => x"80",
           332 => x"da",
           333 => x"91",
           334 => x"02",
           335 => x"0c",
           336 => x"80",
           337 => x"d4",
           338 => x"08",
           339 => x"d4",
           340 => x"08",
           341 => x"3f",
           342 => x"08",
           343 => x"c8",
           344 => x"3d",
           345 => x"d4",
           346 => x"d3",
           347 => x"91",
           348 => x"fd",
           349 => x"53",
           350 => x"08",
           351 => x"52",
           352 => x"08",
           353 => x"51",
           354 => x"d3",
           355 => x"91",
           356 => x"54",
           357 => x"91",
           358 => x"04",
           359 => x"08",
           360 => x"d4",
           361 => x"0d",
           362 => x"d3",
           363 => x"05",
           364 => x"91",
           365 => x"f8",
           366 => x"d3",
           367 => x"05",
           368 => x"d4",
           369 => x"08",
           370 => x"91",
           371 => x"fc",
           372 => x"2e",
           373 => x"0b",
           374 => x"08",
           375 => x"24",
           376 => x"d3",
           377 => x"05",
           378 => x"d3",
           379 => x"05",
           380 => x"d4",
           381 => x"08",
           382 => x"d4",
           383 => x"0c",
           384 => x"91",
           385 => x"fc",
           386 => x"2e",
           387 => x"91",
           388 => x"8c",
           389 => x"d3",
           390 => x"05",
           391 => x"38",
           392 => x"08",
           393 => x"91",
           394 => x"8c",
           395 => x"91",
           396 => x"88",
           397 => x"d3",
           398 => x"05",
           399 => x"d4",
           400 => x"08",
           401 => x"d4",
           402 => x"0c",
           403 => x"08",
           404 => x"81",
           405 => x"d4",
           406 => x"0c",
           407 => x"08",
           408 => x"81",
           409 => x"d4",
           410 => x"0c",
           411 => x"91",
           412 => x"90",
           413 => x"2e",
           414 => x"d3",
           415 => x"05",
           416 => x"d3",
           417 => x"05",
           418 => x"39",
           419 => x"08",
           420 => x"70",
           421 => x"08",
           422 => x"51",
           423 => x"08",
           424 => x"91",
           425 => x"85",
           426 => x"d3",
           427 => x"fc",
           428 => x"79",
           429 => x"05",
           430 => x"57",
           431 => x"83",
           432 => x"38",
           433 => x"51",
           434 => x"a4",
           435 => x"52",
           436 => x"93",
           437 => x"70",
           438 => x"34",
           439 => x"71",
           440 => x"81",
           441 => x"74",
           442 => x"0c",
           443 => x"04",
           444 => x"2b",
           445 => x"71",
           446 => x"51",
           447 => x"72",
           448 => x"72",
           449 => x"05",
           450 => x"71",
           451 => x"53",
           452 => x"70",
           453 => x"0c",
           454 => x"84",
           455 => x"f0",
           456 => x"8f",
           457 => x"83",
           458 => x"38",
           459 => x"84",
           460 => x"fc",
           461 => x"83",
           462 => x"70",
           463 => x"39",
           464 => x"77",
           465 => x"07",
           466 => x"54",
           467 => x"38",
           468 => x"08",
           469 => x"71",
           470 => x"80",
           471 => x"75",
           472 => x"33",
           473 => x"06",
           474 => x"80",
           475 => x"72",
           476 => x"75",
           477 => x"06",
           478 => x"12",
           479 => x"33",
           480 => x"06",
           481 => x"52",
           482 => x"72",
           483 => x"81",
           484 => x"81",
           485 => x"71",
           486 => x"c8",
           487 => x"87",
           488 => x"71",
           489 => x"fb",
           490 => x"06",
           491 => x"82",
           492 => x"51",
           493 => x"97",
           494 => x"84",
           495 => x"54",
           496 => x"75",
           497 => x"38",
           498 => x"52",
           499 => x"80",
           500 => x"c8",
           501 => x"0d",
           502 => x"0d",
           503 => x"52",
           504 => x"52",
           505 => x"91",
           506 => x"81",
           507 => x"07",
           508 => x"52",
           509 => x"e8",
           510 => x"d3",
           511 => x"3d",
           512 => x"3d",
           513 => x"08",
           514 => x"55",
           515 => x"80",
           516 => x"33",
           517 => x"2e",
           518 => x"8c",
           519 => x"70",
           520 => x"70",
           521 => x"38",
           522 => x"39",
           523 => x"80",
           524 => x"53",
           525 => x"83",
           526 => x"70",
           527 => x"2a",
           528 => x"51",
           529 => x"71",
           530 => x"a0",
           531 => x"06",
           532 => x"72",
           533 => x"54",
           534 => x"0c",
           535 => x"91",
           536 => x"86",
           537 => x"fc",
           538 => x"53",
           539 => x"2e",
           540 => x"3d",
           541 => x"72",
           542 => x"3f",
           543 => x"08",
           544 => x"53",
           545 => x"53",
           546 => x"c8",
           547 => x"0d",
           548 => x"0d",
           549 => x"33",
           550 => x"5c",
           551 => x"8b",
           552 => x"38",
           553 => x"ff",
           554 => x"5b",
           555 => x"81",
           556 => x"1c",
           557 => x"5b",
           558 => x"81",
           559 => x"1c",
           560 => x"5b",
           561 => x"81",
           562 => x"1c",
           563 => x"5b",
           564 => x"81",
           565 => x"1c",
           566 => x"5b",
           567 => x"26",
           568 => x"8a",
           569 => x"87",
           570 => x"e7",
           571 => x"38",
           572 => x"59",
           573 => x"58",
           574 => x"57",
           575 => x"56",
           576 => x"55",
           577 => x"54",
           578 => x"53",
           579 => x"91",
           580 => x"94",
           581 => x"c0",
           582 => x"81",
           583 => x"22",
           584 => x"bc",
           585 => x"33",
           586 => x"b8",
           587 => x"33",
           588 => x"b4",
           589 => x"33",
           590 => x"b0",
           591 => x"33",
           592 => x"ac",
           593 => x"33",
           594 => x"a8",
           595 => x"22",
           596 => x"a4",
           597 => x"22",
           598 => x"a0",
           599 => x"0c",
           600 => x"91",
           601 => x"8d",
           602 => x"f5",
           603 => x"5a",
           604 => x"9c",
           605 => x"0c",
           606 => x"bc",
           607 => x"7a",
           608 => x"98",
           609 => x"7a",
           610 => x"87",
           611 => x"08",
           612 => x"1b",
           613 => x"98",
           614 => x"7a",
           615 => x"87",
           616 => x"08",
           617 => x"1b",
           618 => x"98",
           619 => x"7a",
           620 => x"87",
           621 => x"08",
           622 => x"1b",
           623 => x"98",
           624 => x"7a",
           625 => x"80",
           626 => x"1a",
           627 => x"1a",
           628 => x"1a",
           629 => x"1a",
           630 => x"1a",
           631 => x"1a",
           632 => x"1a",
           633 => x"22",
           634 => x"a8",
           635 => x"3f",
           636 => x"04",
           637 => x"02",
           638 => x"70",
           639 => x"2a",
           640 => x"70",
           641 => x"cb",
           642 => x"3d",
           643 => x"3d",
           644 => x"0b",
           645 => x"33",
           646 => x"c0",
           647 => x"72",
           648 => x"38",
           649 => x"94",
           650 => x"70",
           651 => x"81",
           652 => x"52",
           653 => x"8c",
           654 => x"2a",
           655 => x"51",
           656 => x"38",
           657 => x"81",
           658 => x"06",
           659 => x"80",
           660 => x"71",
           661 => x"81",
           662 => x"70",
           663 => x"0b",
           664 => x"c0",
           665 => x"c0",
           666 => x"70",
           667 => x"38",
           668 => x"90",
           669 => x"0c",
           670 => x"c8",
           671 => x"0d",
           672 => x"0d",
           673 => x"33",
           674 => x"cb",
           675 => x"54",
           676 => x"84",
           677 => x"2e",
           678 => x"c0",
           679 => x"70",
           680 => x"2a",
           681 => x"51",
           682 => x"80",
           683 => x"71",
           684 => x"81",
           685 => x"70",
           686 => x"96",
           687 => x"70",
           688 => x"51",
           689 => x"8d",
           690 => x"2a",
           691 => x"51",
           692 => x"bc",
           693 => x"91",
           694 => x"51",
           695 => x"80",
           696 => x"2e",
           697 => x"c0",
           698 => x"73",
           699 => x"3d",
           700 => x"3d",
           701 => x"80",
           702 => x"56",
           703 => x"80",
           704 => x"70",
           705 => x"33",
           706 => x"cb",
           707 => x"55",
           708 => x"84",
           709 => x"2e",
           710 => x"c0",
           711 => x"70",
           712 => x"2a",
           713 => x"51",
           714 => x"80",
           715 => x"71",
           716 => x"81",
           717 => x"70",
           718 => x"96",
           719 => x"70",
           720 => x"51",
           721 => x"8d",
           722 => x"2a",
           723 => x"51",
           724 => x"bc",
           725 => x"91",
           726 => x"51",
           727 => x"80",
           728 => x"2e",
           729 => x"c0",
           730 => x"74",
           731 => x"16",
           732 => x"56",
           733 => x"38",
           734 => x"c8",
           735 => x"0d",
           736 => x"0d",
           737 => x"cb",
           738 => x"87",
           739 => x"51",
           740 => x"86",
           741 => x"94",
           742 => x"08",
           743 => x"70",
           744 => x"51",
           745 => x"2e",
           746 => x"0b",
           747 => x"33",
           748 => x"94",
           749 => x"80",
           750 => x"87",
           751 => x"52",
           752 => x"81",
           753 => x"d3",
           754 => x"83",
           755 => x"ff",
           756 => x"0b",
           757 => x"33",
           758 => x"94",
           759 => x"80",
           760 => x"87",
           761 => x"52",
           762 => x"82",
           763 => x"06",
           764 => x"ff",
           765 => x"2e",
           766 => x"0b",
           767 => x"33",
           768 => x"94",
           769 => x"80",
           770 => x"87",
           771 => x"52",
           772 => x"98",
           773 => x"2c",
           774 => x"71",
           775 => x"0c",
           776 => x"04",
           777 => x"87",
           778 => x"70",
           779 => x"2a",
           780 => x"52",
           781 => x"2e",
           782 => x"91",
           783 => x"87",
           784 => x"08",
           785 => x"11",
           786 => x"a0",
           787 => x"52",
           788 => x"c0",
           789 => x"71",
           790 => x"11",
           791 => x"90",
           792 => x"52",
           793 => x"c0",
           794 => x"71",
           795 => x"11",
           796 => x"98",
           797 => x"52",
           798 => x"c0",
           799 => x"71",
           800 => x"11",
           801 => x"a8",
           802 => x"52",
           803 => x"c0",
           804 => x"71",
           805 => x"08",
           806 => x"a4",
           807 => x"12",
           808 => x"84",
           809 => x"51",
           810 => x"13",
           811 => x"52",
           812 => x"c0",
           813 => x"70",
           814 => x"51",
           815 => x"80",
           816 => x"81",
           817 => x"34",
           818 => x"c0",
           819 => x"70",
           820 => x"06",
           821 => x"70",
           822 => x"38",
           823 => x"91",
           824 => x"80",
           825 => x"9e",
           826 => x"80",
           827 => x"51",
           828 => x"80",
           829 => x"81",
           830 => x"cb",
           831 => x"0b",
           832 => x"88",
           833 => x"80",
           834 => x"52",
           835 => x"83",
           836 => x"71",
           837 => x"34",
           838 => x"c0",
           839 => x"70",
           840 => x"51",
           841 => x"80",
           842 => x"81",
           843 => x"cb",
           844 => x"0b",
           845 => x"88",
           846 => x"80",
           847 => x"52",
           848 => x"83",
           849 => x"71",
           850 => x"34",
           851 => x"c0",
           852 => x"70",
           853 => x"51",
           854 => x"80",
           855 => x"81",
           856 => x"cb",
           857 => x"0b",
           858 => x"88",
           859 => x"80",
           860 => x"52",
           861 => x"83",
           862 => x"71",
           863 => x"34",
           864 => x"52",
           865 => x"88",
           866 => x"80",
           867 => x"86",
           868 => x"52",
           869 => x"70",
           870 => x"34",
           871 => x"73",
           872 => x"06",
           873 => x"70",
           874 => x"38",
           875 => x"74",
           876 => x"87",
           877 => x"08",
           878 => x"51",
           879 => x"80",
           880 => x"81",
           881 => x"cb",
           882 => x"c0",
           883 => x"70",
           884 => x"51",
           885 => x"fc",
           886 => x"0d",
           887 => x"0d",
           888 => x"51",
           889 => x"91",
           890 => x"54",
           891 => x"88",
           892 => x"d4",
           893 => x"3f",
           894 => x"51",
           895 => x"91",
           896 => x"33",
           897 => x"80",
           898 => x"d7",
           899 => x"91",
           900 => x"52",
           901 => x"51",
           902 => x"91",
           903 => x"33",
           904 => x"80",
           905 => x"de",
           906 => x"da",
           907 => x"91",
           908 => x"89",
           909 => x"cb",
           910 => x"55",
           911 => x"38",
           912 => x"54",
           913 => x"93",
           914 => x"d8",
           915 => x"fc",
           916 => x"54",
           917 => x"51",
           918 => x"91",
           919 => x"54",
           920 => x"88",
           921 => x"f0",
           922 => x"3f",
           923 => x"33",
           924 => x"2e",
           925 => x"b7",
           926 => x"a8",
           927 => x"f7",
           928 => x"80",
           929 => x"91",
           930 => x"83",
           931 => x"cb",
           932 => x"55",
           933 => x"2e",
           934 => x"15",
           935 => x"b8",
           936 => x"fa",
           937 => x"fa",
           938 => x"80",
           939 => x"91",
           940 => x"82",
           941 => x"cb",
           942 => x"55",
           943 => x"2e",
           944 => x"15",
           945 => x"b8",
           946 => x"d2",
           947 => x"ec",
           948 => x"3f",
           949 => x"70",
           950 => x"05",
           951 => x"91",
           952 => x"55",
           953 => x"3f",
           954 => x"91",
           955 => x"88",
           956 => x"15",
           957 => x"b9",
           958 => x"a2",
           959 => x"22",
           960 => x"f0",
           961 => x"3f",
           962 => x"52",
           963 => x"51",
           964 => x"86",
           965 => x"ff",
           966 => x"8e",
           967 => x"71",
           968 => x"38",
           969 => x"0b",
           970 => x"c4",
           971 => x"08",
           972 => x"c0",
           973 => x"3f",
           974 => x"ba",
           975 => x"b2",
           976 => x"91",
           977 => x"f7",
           978 => x"39",
           979 => x"51",
           980 => x"91",
           981 => x"dc",
           982 => x"3f",
           983 => x"ba",
           984 => x"8e",
           985 => x"0d",
           986 => x"80",
           987 => x"0b",
           988 => x"84",
           989 => x"3d",
           990 => x"96",
           991 => x"52",
           992 => x"0c",
           993 => x"70",
           994 => x"0c",
           995 => x"3d",
           996 => x"3d",
           997 => x"96",
           998 => x"91",
           999 => x"52",
          1000 => x"73",
          1001 => x"cc",
          1002 => x"70",
          1003 => x"0c",
          1004 => x"83",
          1005 => x"91",
          1006 => x"87",
          1007 => x"0c",
          1008 => x"0d",
          1009 => x"33",
          1010 => x"2e",
          1011 => x"85",
          1012 => x"ed",
          1013 => x"e0",
          1014 => x"95",
          1015 => x"e0",
          1016 => x"72",
          1017 => x"e0",
          1018 => x"91",
          1019 => x"92",
          1020 => x"d8",
          1021 => x"8a",
          1022 => x"91",
          1023 => x"52",
          1024 => x"3d",
          1025 => x"3d",
          1026 => x"05",
          1027 => x"d8",
          1028 => x"d3",
          1029 => x"51",
          1030 => x"72",
          1031 => x"0c",
          1032 => x"04",
          1033 => x"74",
          1034 => x"53",
          1035 => x"91",
          1036 => x"81",
          1037 => x"51",
          1038 => x"72",
          1039 => x"f1",
          1040 => x"0d",
          1041 => x"0d",
          1042 => x"d8",
          1043 => x"d3",
          1044 => x"33",
          1045 => x"71",
          1046 => x"38",
          1047 => x"05",
          1048 => x"fe",
          1049 => x"33",
          1050 => x"38",
          1051 => x"d8",
          1052 => x"0d",
          1053 => x"0d",
          1054 => x"59",
          1055 => x"05",
          1056 => x"75",
          1057 => x"92",
          1058 => x"2e",
          1059 => x"51",
          1060 => x"e8",
          1061 => x"7a",
          1062 => x"5c",
          1063 => x"5a",
          1064 => x"09",
          1065 => x"38",
          1066 => x"81",
          1067 => x"57",
          1068 => x"75",
          1069 => x"81",
          1070 => x"82",
          1071 => x"05",
          1072 => x"5d",
          1073 => x"09",
          1074 => x"38",
          1075 => x"71",
          1076 => x"81",
          1077 => x"59",
          1078 => x"9f",
          1079 => x"53",
          1080 => x"97",
          1081 => x"29",
          1082 => x"79",
          1083 => x"5b",
          1084 => x"55",
          1085 => x"73",
          1086 => x"75",
          1087 => x"70",
          1088 => x"07",
          1089 => x"80",
          1090 => x"30",
          1091 => x"80",
          1092 => x"53",
          1093 => x"54",
          1094 => x"2e",
          1095 => x"84",
          1096 => x"81",
          1097 => x"57",
          1098 => x"2e",
          1099 => x"75",
          1100 => x"76",
          1101 => x"e0",
          1102 => x"ff",
          1103 => x"ff",
          1104 => x"72",
          1105 => x"98",
          1106 => x"10",
          1107 => x"05",
          1108 => x"04",
          1109 => x"71",
          1110 => x"53",
          1111 => x"54",
          1112 => x"2e",
          1113 => x"14",
          1114 => x"33",
          1115 => x"72",
          1116 => x"81",
          1117 => x"06",
          1118 => x"a3",
          1119 => x"15",
          1120 => x"7a",
          1121 => x"7c",
          1122 => x"06",
          1123 => x"fc",
          1124 => x"8b",
          1125 => x"15",
          1126 => x"73",
          1127 => x"74",
          1128 => x"3f",
          1129 => x"55",
          1130 => x"27",
          1131 => x"a0",
          1132 => x"3f",
          1133 => x"55",
          1134 => x"26",
          1135 => x"bc",
          1136 => x"1d",
          1137 => x"53",
          1138 => x"f5",
          1139 => x"39",
          1140 => x"39",
          1141 => x"39",
          1142 => x"39",
          1143 => x"39",
          1144 => x"dd",
          1145 => x"39",
          1146 => x"70",
          1147 => x"53",
          1148 => x"8b",
          1149 => x"1d",
          1150 => x"5d",
          1151 => x"74",
          1152 => x"09",
          1153 => x"38",
          1154 => x"71",
          1155 => x"53",
          1156 => x"84",
          1157 => x"59",
          1158 => x"80",
          1159 => x"30",
          1160 => x"80",
          1161 => x"7b",
          1162 => x"52",
          1163 => x"80",
          1164 => x"76",
          1165 => x"07",
          1166 => x"58",
          1167 => x"51",
          1168 => x"91",
          1169 => x"81",
          1170 => x"53",
          1171 => x"e5",
          1172 => x"d3",
          1173 => x"89",
          1174 => x"38",
          1175 => x"70",
          1176 => x"57",
          1177 => x"80",
          1178 => x"38",
          1179 => x"81",
          1180 => x"53",
          1181 => x"05",
          1182 => x"16",
          1183 => x"74",
          1184 => x"77",
          1185 => x"07",
          1186 => x"9f",
          1187 => x"51",
          1188 => x"72",
          1189 => x"7c",
          1190 => x"81",
          1191 => x"72",
          1192 => x"38",
          1193 => x"05",
          1194 => x"ad",
          1195 => x"18",
          1196 => x"81",
          1197 => x"b0",
          1198 => x"38",
          1199 => x"81",
          1200 => x"06",
          1201 => x"a3",
          1202 => x"15",
          1203 => x"7a",
          1204 => x"7c",
          1205 => x"06",
          1206 => x"f9",
          1207 => x"8b",
          1208 => x"15",
          1209 => x"73",
          1210 => x"ff",
          1211 => x"e0",
          1212 => x"33",
          1213 => x"f9",
          1214 => x"ef",
          1215 => x"15",
          1216 => x"7a",
          1217 => x"38",
          1218 => x"b5",
          1219 => x"15",
          1220 => x"73",
          1221 => x"fa",
          1222 => x"3d",
          1223 => x"3d",
          1224 => x"70",
          1225 => x"52",
          1226 => x"73",
          1227 => x"3f",
          1228 => x"04",
          1229 => x"74",
          1230 => x"0c",
          1231 => x"05",
          1232 => x"fa",
          1233 => x"d3",
          1234 => x"80",
          1235 => x"0b",
          1236 => x"0c",
          1237 => x"04",
          1238 => x"91",
          1239 => x"76",
          1240 => x"0c",
          1241 => x"05",
          1242 => x"53",
          1243 => x"72",
          1244 => x"0c",
          1245 => x"04",
          1246 => x"78",
          1247 => x"80",
          1248 => x"dc",
          1249 => x"80",
          1250 => x"39",
          1251 => x"f3",
          1252 => x"91",
          1253 => x"52",
          1254 => x"d3",
          1255 => x"ff",
          1256 => x"80",
          1257 => x"73",
          1258 => x"ca",
          1259 => x"32",
          1260 => x"30",
          1261 => x"9f",
          1262 => x"25",
          1263 => x"51",
          1264 => x"2e",
          1265 => x"15",
          1266 => x"06",
          1267 => x"f1",
          1268 => x"9f",
          1269 => x"bb",
          1270 => x"52",
          1271 => x"ff",
          1272 => x"15",
          1273 => x"34",
          1274 => x"81",
          1275 => x"55",
          1276 => x"ff",
          1277 => x"17",
          1278 => x"34",
          1279 => x"c1",
          1280 => x"72",
          1281 => x"0c",
          1282 => x"04",
          1283 => x"91",
          1284 => x"75",
          1285 => x"0c",
          1286 => x"52",
          1287 => x"3f",
          1288 => x"dc",
          1289 => x"0d",
          1290 => x"0d",
          1291 => x"55",
          1292 => x"0c",
          1293 => x"33",
          1294 => x"73",
          1295 => x"81",
          1296 => x"74",
          1297 => x"75",
          1298 => x"70",
          1299 => x"73",
          1300 => x"38",
          1301 => x"09",
          1302 => x"38",
          1303 => x"11",
          1304 => x"08",
          1305 => x"54",
          1306 => x"2e",
          1307 => x"80",
          1308 => x"08",
          1309 => x"0c",
          1310 => x"33",
          1311 => x"80",
          1312 => x"38",
          1313 => x"2e",
          1314 => x"a1",
          1315 => x"81",
          1316 => x"75",
          1317 => x"56",
          1318 => x"c1",
          1319 => x"08",
          1320 => x"0c",
          1321 => x"33",
          1322 => x"b1",
          1323 => x"a0",
          1324 => x"82",
          1325 => x"53",
          1326 => x"57",
          1327 => x"9d",
          1328 => x"39",
          1329 => x"80",
          1330 => x"26",
          1331 => x"8b",
          1332 => x"80",
          1333 => x"56",
          1334 => x"8a",
          1335 => x"a0",
          1336 => x"c5",
          1337 => x"74",
          1338 => x"e0",
          1339 => x"ff",
          1340 => x"d0",
          1341 => x"ff",
          1342 => x"90",
          1343 => x"38",
          1344 => x"81",
          1345 => x"53",
          1346 => x"c5",
          1347 => x"27",
          1348 => x"76",
          1349 => x"08",
          1350 => x"0c",
          1351 => x"33",
          1352 => x"73",
          1353 => x"bd",
          1354 => x"2e",
          1355 => x"30",
          1356 => x"0c",
          1357 => x"91",
          1358 => x"8a",
          1359 => x"f8",
          1360 => x"7c",
          1361 => x"70",
          1362 => x"08",
          1363 => x"54",
          1364 => x"2e",
          1365 => x"92",
          1366 => x"81",
          1367 => x"74",
          1368 => x"55",
          1369 => x"2e",
          1370 => x"ad",
          1371 => x"06",
          1372 => x"75",
          1373 => x"0c",
          1374 => x"33",
          1375 => x"73",
          1376 => x"81",
          1377 => x"38",
          1378 => x"05",
          1379 => x"08",
          1380 => x"53",
          1381 => x"2e",
          1382 => x"80",
          1383 => x"81",
          1384 => x"90",
          1385 => x"76",
          1386 => x"70",
          1387 => x"57",
          1388 => x"82",
          1389 => x"05",
          1390 => x"08",
          1391 => x"54",
          1392 => x"81",
          1393 => x"27",
          1394 => x"d0",
          1395 => x"56",
          1396 => x"73",
          1397 => x"80",
          1398 => x"14",
          1399 => x"72",
          1400 => x"e8",
          1401 => x"80",
          1402 => x"39",
          1403 => x"dc",
          1404 => x"80",
          1405 => x"27",
          1406 => x"80",
          1407 => x"89",
          1408 => x"70",
          1409 => x"55",
          1410 => x"70",
          1411 => x"55",
          1412 => x"27",
          1413 => x"14",
          1414 => x"06",
          1415 => x"74",
          1416 => x"73",
          1417 => x"38",
          1418 => x"14",
          1419 => x"05",
          1420 => x"08",
          1421 => x"54",
          1422 => x"26",
          1423 => x"77",
          1424 => x"38",
          1425 => x"75",
          1426 => x"56",
          1427 => x"c8",
          1428 => x"0d",
          1429 => x"0d",
          1430 => x"33",
          1431 => x"70",
          1432 => x"38",
          1433 => x"11",
          1434 => x"91",
          1435 => x"83",
          1436 => x"fd",
          1437 => x"97",
          1438 => x"84",
          1439 => x"33",
          1440 => x"51",
          1441 => x"80",
          1442 => x"90",
          1443 => x"92",
          1444 => x"88",
          1445 => x"2e",
          1446 => x"88",
          1447 => x"0c",
          1448 => x"87",
          1449 => x"05",
          1450 => x"0c",
          1451 => x"c0",
          1452 => x"70",
          1453 => x"98",
          1454 => x"08",
          1455 => x"51",
          1456 => x"2e",
          1457 => x"08",
          1458 => x"38",
          1459 => x"87",
          1460 => x"05",
          1461 => x"80",
          1462 => x"51",
          1463 => x"87",
          1464 => x"08",
          1465 => x"2e",
          1466 => x"91",
          1467 => x"34",
          1468 => x"13",
          1469 => x"91",
          1470 => x"85",
          1471 => x"f2",
          1472 => x"63",
          1473 => x"05",
          1474 => x"33",
          1475 => x"58",
          1476 => x"5b",
          1477 => x"91",
          1478 => x"81",
          1479 => x"52",
          1480 => x"38",
          1481 => x"5d",
          1482 => x"8c",
          1483 => x"87",
          1484 => x"11",
          1485 => x"84",
          1486 => x"5c",
          1487 => x"85",
          1488 => x"c0",
          1489 => x"7c",
          1490 => x"84",
          1491 => x"08",
          1492 => x"70",
          1493 => x"53",
          1494 => x"2e",
          1495 => x"08",
          1496 => x"70",
          1497 => x"34",
          1498 => x"73",
          1499 => x"71",
          1500 => x"38",
          1501 => x"71",
          1502 => x"08",
          1503 => x"2e",
          1504 => x"84",
          1505 => x"38",
          1506 => x"87",
          1507 => x"1e",
          1508 => x"70",
          1509 => x"52",
          1510 => x"ff",
          1511 => x"39",
          1512 => x"81",
          1513 => x"ff",
          1514 => x"5c",
          1515 => x"90",
          1516 => x"80",
          1517 => x"71",
          1518 => x"7d",
          1519 => x"38",
          1520 => x"80",
          1521 => x"80",
          1522 => x"81",
          1523 => x"73",
          1524 => x"0c",
          1525 => x"04",
          1526 => x"60",
          1527 => x"8c",
          1528 => x"33",
          1529 => x"57",
          1530 => x"5a",
          1531 => x"91",
          1532 => x"81",
          1533 => x"52",
          1534 => x"38",
          1535 => x"c0",
          1536 => x"84",
          1537 => x"92",
          1538 => x"c0",
          1539 => x"72",
          1540 => x"5a",
          1541 => x"0c",
          1542 => x"80",
          1543 => x"0c",
          1544 => x"0c",
          1545 => x"08",
          1546 => x"70",
          1547 => x"53",
          1548 => x"2e",
          1549 => x"70",
          1550 => x"33",
          1551 => x"13",
          1552 => x"2a",
          1553 => x"51",
          1554 => x"2e",
          1555 => x"08",
          1556 => x"38",
          1557 => x"71",
          1558 => x"38",
          1559 => x"2e",
          1560 => x"75",
          1561 => x"92",
          1562 => x"72",
          1563 => x"06",
          1564 => x"f7",
          1565 => x"5a",
          1566 => x"1c",
          1567 => x"06",
          1568 => x"5d",
          1569 => x"80",
          1570 => x"73",
          1571 => x"06",
          1572 => x"38",
          1573 => x"fe",
          1574 => x"fc",
          1575 => x"52",
          1576 => x"83",
          1577 => x"71",
          1578 => x"d3",
          1579 => x"3d",
          1580 => x"3d",
          1581 => x"84",
          1582 => x"33",
          1583 => x"b3",
          1584 => x"54",
          1585 => x"fb",
          1586 => x"d3",
          1587 => x"06",
          1588 => x"71",
          1589 => x"54",
          1590 => x"a2",
          1591 => x"24",
          1592 => x"80",
          1593 => x"a7",
          1594 => x"2e",
          1595 => x"39",
          1596 => x"87",
          1597 => x"05",
          1598 => x"52",
          1599 => x"80",
          1600 => x"80",
          1601 => x"81",
          1602 => x"80",
          1603 => x"84",
          1604 => x"d3",
          1605 => x"3d",
          1606 => x"3d",
          1607 => x"33",
          1608 => x"70",
          1609 => x"07",
          1610 => x"0c",
          1611 => x"83",
          1612 => x"fd",
          1613 => x"83",
          1614 => x"12",
          1615 => x"2b",
          1616 => x"07",
          1617 => x"71",
          1618 => x"71",
          1619 => x"91",
          1620 => x"51",
          1621 => x"52",
          1622 => x"04",
          1623 => x"73",
          1624 => x"92",
          1625 => x"52",
          1626 => x"81",
          1627 => x"70",
          1628 => x"70",
          1629 => x"3d",
          1630 => x"3d",
          1631 => x"52",
          1632 => x"70",
          1633 => x"34",
          1634 => x"51",
          1635 => x"81",
          1636 => x"70",
          1637 => x"70",
          1638 => x"05",
          1639 => x"88",
          1640 => x"72",
          1641 => x"0d",
          1642 => x"0d",
          1643 => x"54",
          1644 => x"80",
          1645 => x"71",
          1646 => x"53",
          1647 => x"81",
          1648 => x"ff",
          1649 => x"ef",
          1650 => x"0d",
          1651 => x"0d",
          1652 => x"54",
          1653 => x"72",
          1654 => x"54",
          1655 => x"51",
          1656 => x"84",
          1657 => x"fc",
          1658 => x"77",
          1659 => x"53",
          1660 => x"05",
          1661 => x"70",
          1662 => x"33",
          1663 => x"ff",
          1664 => x"52",
          1665 => x"2e",
          1666 => x"80",
          1667 => x"71",
          1668 => x"0c",
          1669 => x"04",
          1670 => x"74",
          1671 => x"53",
          1672 => x"80",
          1673 => x"70",
          1674 => x"38",
          1675 => x"33",
          1676 => x"80",
          1677 => x"70",
          1678 => x"81",
          1679 => x"71",
          1680 => x"c8",
          1681 => x"0d",
          1682 => x"91",
          1683 => x"04",
          1684 => x"d3",
          1685 => x"f9",
          1686 => x"56",
          1687 => x"17",
          1688 => x"74",
          1689 => x"d7",
          1690 => x"b0",
          1691 => x"b4",
          1692 => x"81",
          1693 => x"57",
          1694 => x"91",
          1695 => x"78",
          1696 => x"06",
          1697 => x"d3",
          1698 => x"17",
          1699 => x"08",
          1700 => x"31",
          1701 => x"17",
          1702 => x"38",
          1703 => x"55",
          1704 => x"09",
          1705 => x"38",
          1706 => x"16",
          1707 => x"08",
          1708 => x"52",
          1709 => x"51",
          1710 => x"83",
          1711 => x"77",
          1712 => x"0c",
          1713 => x"04",
          1714 => x"78",
          1715 => x"80",
          1716 => x"08",
          1717 => x"38",
          1718 => x"fb",
          1719 => x"c8",
          1720 => x"d3",
          1721 => x"38",
          1722 => x"53",
          1723 => x"81",
          1724 => x"f8",
          1725 => x"d3",
          1726 => x"2e",
          1727 => x"55",
          1728 => x"b0",
          1729 => x"91",
          1730 => x"88",
          1731 => x"f8",
          1732 => x"70",
          1733 => x"bf",
          1734 => x"c8",
          1735 => x"d3",
          1736 => x"91",
          1737 => x"55",
          1738 => x"09",
          1739 => x"f0",
          1740 => x"33",
          1741 => x"2e",
          1742 => x"80",
          1743 => x"80",
          1744 => x"c8",
          1745 => x"17",
          1746 => x"fd",
          1747 => x"d4",
          1748 => x"b2",
          1749 => x"84",
          1750 => x"85",
          1751 => x"75",
          1752 => x"3f",
          1753 => x"e4",
          1754 => x"98",
          1755 => x"8a",
          1756 => x"08",
          1757 => x"17",
          1758 => x"3f",
          1759 => x"52",
          1760 => x"51",
          1761 => x"a0",
          1762 => x"05",
          1763 => x"0c",
          1764 => x"75",
          1765 => x"33",
          1766 => x"3f",
          1767 => x"34",
          1768 => x"52",
          1769 => x"51",
          1770 => x"91",
          1771 => x"80",
          1772 => x"81",
          1773 => x"d3",
          1774 => x"3d",
          1775 => x"3d",
          1776 => x"1a",
          1777 => x"fe",
          1778 => x"54",
          1779 => x"73",
          1780 => x"8a",
          1781 => x"76",
          1782 => x"08",
          1783 => x"75",
          1784 => x"0c",
          1785 => x"04",
          1786 => x"7a",
          1787 => x"56",
          1788 => x"75",
          1789 => x"98",
          1790 => x"26",
          1791 => x"56",
          1792 => x"ff",
          1793 => x"56",
          1794 => x"80",
          1795 => x"82",
          1796 => x"72",
          1797 => x"38",
          1798 => x"72",
          1799 => x"8e",
          1800 => x"39",
          1801 => x"15",
          1802 => x"a4",
          1803 => x"53",
          1804 => x"fd",
          1805 => x"d3",
          1806 => x"9f",
          1807 => x"ff",
          1808 => x"11",
          1809 => x"70",
          1810 => x"18",
          1811 => x"76",
          1812 => x"53",
          1813 => x"91",
          1814 => x"80",
          1815 => x"83",
          1816 => x"b4",
          1817 => x"88",
          1818 => x"77",
          1819 => x"84",
          1820 => x"5a",
          1821 => x"80",
          1822 => x"9f",
          1823 => x"80",
          1824 => x"88",
          1825 => x"08",
          1826 => x"51",
          1827 => x"91",
          1828 => x"80",
          1829 => x"15",
          1830 => x"74",
          1831 => x"51",
          1832 => x"91",
          1833 => x"83",
          1834 => x"56",
          1835 => x"87",
          1836 => x"08",
          1837 => x"51",
          1838 => x"91",
          1839 => x"9b",
          1840 => x"2b",
          1841 => x"74",
          1842 => x"51",
          1843 => x"91",
          1844 => x"f0",
          1845 => x"83",
          1846 => x"75",
          1847 => x"0c",
          1848 => x"04",
          1849 => x"7b",
          1850 => x"55",
          1851 => x"81",
          1852 => x"af",
          1853 => x"16",
          1854 => x"a7",
          1855 => x"53",
          1856 => x"81",
          1857 => x"77",
          1858 => x"72",
          1859 => x"38",
          1860 => x"72",
          1861 => x"c9",
          1862 => x"39",
          1863 => x"14",
          1864 => x"a4",
          1865 => x"53",
          1866 => x"fb",
          1867 => x"d3",
          1868 => x"91",
          1869 => x"81",
          1870 => x"83",
          1871 => x"b4",
          1872 => x"76",
          1873 => x"5b",
          1874 => x"57",
          1875 => x"8f",
          1876 => x"2b",
          1877 => x"78",
          1878 => x"71",
          1879 => x"76",
          1880 => x"0b",
          1881 => x"78",
          1882 => x"16",
          1883 => x"74",
          1884 => x"3f",
          1885 => x"08",
          1886 => x"c8",
          1887 => x"38",
          1888 => x"06",
          1889 => x"75",
          1890 => x"84",
          1891 => x"51",
          1892 => x"38",
          1893 => x"78",
          1894 => x"06",
          1895 => x"06",
          1896 => x"78",
          1897 => x"83",
          1898 => x"f7",
          1899 => x"2a",
          1900 => x"05",
          1901 => x"fa",
          1902 => x"d3",
          1903 => x"91",
          1904 => x"80",
          1905 => x"83",
          1906 => x"52",
          1907 => x"ff",
          1908 => x"b4",
          1909 => x"84",
          1910 => x"83",
          1911 => x"c3",
          1912 => x"2a",
          1913 => x"05",
          1914 => x"f9",
          1915 => x"d3",
          1916 => x"91",
          1917 => x"ab",
          1918 => x"0a",
          1919 => x"2b",
          1920 => x"76",
          1921 => x"70",
          1922 => x"56",
          1923 => x"91",
          1924 => x"8f",
          1925 => x"07",
          1926 => x"f6",
          1927 => x"0b",
          1928 => x"76",
          1929 => x"0c",
          1930 => x"04",
          1931 => x"79",
          1932 => x"08",
          1933 => x"57",
          1934 => x"88",
          1935 => x"08",
          1936 => x"38",
          1937 => x"8e",
          1938 => x"2e",
          1939 => x"53",
          1940 => x"51",
          1941 => x"91",
          1942 => x"56",
          1943 => x"08",
          1944 => x"93",
          1945 => x"80",
          1946 => x"56",
          1947 => x"91",
          1948 => x"56",
          1949 => x"73",
          1950 => x"fa",
          1951 => x"d3",
          1952 => x"91",
          1953 => x"80",
          1954 => x"38",
          1955 => x"08",
          1956 => x"38",
          1957 => x"08",
          1958 => x"38",
          1959 => x"52",
          1960 => x"c0",
          1961 => x"c8",
          1962 => x"98",
          1963 => x"05",
          1964 => x"08",
          1965 => x"38",
          1966 => x"81",
          1967 => x"0c",
          1968 => x"81",
          1969 => x"84",
          1970 => x"54",
          1971 => x"76",
          1972 => x"38",
          1973 => x"91",
          1974 => x"89",
          1975 => x"f5",
          1976 => x"7f",
          1977 => x"5c",
          1978 => x"38",
          1979 => x"58",
          1980 => x"88",
          1981 => x"08",
          1982 => x"38",
          1983 => x"39",
          1984 => x"51",
          1985 => x"81",
          1986 => x"d3",
          1987 => x"82",
          1988 => x"d3",
          1989 => x"91",
          1990 => x"ff",
          1991 => x"38",
          1992 => x"08",
          1993 => x"08",
          1994 => x"08",
          1995 => x"38",
          1996 => x"55",
          1997 => x"75",
          1998 => x"38",
          1999 => x"7b",
          2000 => x"06",
          2001 => x"81",
          2002 => x"19",
          2003 => x"83",
          2004 => x"76",
          2005 => x"f9",
          2006 => x"d3",
          2007 => x"80",
          2008 => x"c8",
          2009 => x"09",
          2010 => x"38",
          2011 => x"08",
          2012 => x"32",
          2013 => x"72",
          2014 => x"70",
          2015 => x"53",
          2016 => x"54",
          2017 => x"38",
          2018 => x"95",
          2019 => x"08",
          2020 => x"27",
          2021 => x"98",
          2022 => x"83",
          2023 => x"80",
          2024 => x"de",
          2025 => x"81",
          2026 => x"19",
          2027 => x"89",
          2028 => x"76",
          2029 => x"b6",
          2030 => x"7b",
          2031 => x"3f",
          2032 => x"08",
          2033 => x"c8",
          2034 => x"b6",
          2035 => x"91",
          2036 => x"81",
          2037 => x"06",
          2038 => x"d3",
          2039 => x"75",
          2040 => x"30",
          2041 => x"80",
          2042 => x"07",
          2043 => x"54",
          2044 => x"38",
          2045 => x"09",
          2046 => x"ab",
          2047 => x"80",
          2048 => x"53",
          2049 => x"51",
          2050 => x"91",
          2051 => x"91",
          2052 => x"30",
          2053 => x"c8",
          2054 => x"25",
          2055 => x"7f",
          2056 => x"72",
          2057 => x"51",
          2058 => x"80",
          2059 => x"76",
          2060 => x"78",
          2061 => x"3f",
          2062 => x"08",
          2063 => x"38",
          2064 => x"0c",
          2065 => x"fe",
          2066 => x"19",
          2067 => x"89",
          2068 => x"08",
          2069 => x"1a",
          2070 => x"33",
          2071 => x"73",
          2072 => x"94",
          2073 => x"75",
          2074 => x"38",
          2075 => x"55",
          2076 => x"55",
          2077 => x"57",
          2078 => x"91",
          2079 => x"8d",
          2080 => x"f7",
          2081 => x"70",
          2082 => x"cb",
          2083 => x"91",
          2084 => x"80",
          2085 => x"52",
          2086 => x"a2",
          2087 => x"c8",
          2088 => x"c8",
          2089 => x"0c",
          2090 => x"53",
          2091 => x"17",
          2092 => x"f2",
          2093 => x"59",
          2094 => x"56",
          2095 => x"16",
          2096 => x"22",
          2097 => x"27",
          2098 => x"54",
          2099 => x"78",
          2100 => x"33",
          2101 => x"3f",
          2102 => x"08",
          2103 => x"38",
          2104 => x"18",
          2105 => x"74",
          2106 => x"38",
          2107 => x"55",
          2108 => x"c8",
          2109 => x"0d",
          2110 => x"0d",
          2111 => x"08",
          2112 => x"74",
          2113 => x"26",
          2114 => x"9f",
          2115 => x"80",
          2116 => x"82",
          2117 => x"39",
          2118 => x"0c",
          2119 => x"54",
          2120 => x"75",
          2121 => x"73",
          2122 => x"a8",
          2123 => x"73",
          2124 => x"85",
          2125 => x"0b",
          2126 => x"5a",
          2127 => x"27",
          2128 => x"a8",
          2129 => x"18",
          2130 => x"39",
          2131 => x"70",
          2132 => x"58",
          2133 => x"b6",
          2134 => x"76",
          2135 => x"3f",
          2136 => x"08",
          2137 => x"c8",
          2138 => x"bf",
          2139 => x"91",
          2140 => x"27",
          2141 => x"16",
          2142 => x"c8",
          2143 => x"38",
          2144 => x"c1",
          2145 => x"31",
          2146 => x"27",
          2147 => x"52",
          2148 => x"aa",
          2149 => x"c8",
          2150 => x"0c",
          2151 => x"0c",
          2152 => x"17",
          2153 => x"9d",
          2154 => x"81",
          2155 => x"74",
          2156 => x"18",
          2157 => x"18",
          2158 => x"ff",
          2159 => x"05",
          2160 => x"80",
          2161 => x"d3",
          2162 => x"3d",
          2163 => x"3d",
          2164 => x"71",
          2165 => x"08",
          2166 => x"59",
          2167 => x"80",
          2168 => x"86",
          2169 => x"98",
          2170 => x"53",
          2171 => x"80",
          2172 => x"38",
          2173 => x"06",
          2174 => x"c1",
          2175 => x"08",
          2176 => x"16",
          2177 => x"08",
          2178 => x"85",
          2179 => x"22",
          2180 => x"73",
          2181 => x"38",
          2182 => x"0c",
          2183 => x"ad",
          2184 => x"22",
          2185 => x"89",
          2186 => x"53",
          2187 => x"38",
          2188 => x"52",
          2189 => x"b0",
          2190 => x"c8",
          2191 => x"53",
          2192 => x"d3",
          2193 => x"81",
          2194 => x"53",
          2195 => x"08",
          2196 => x"f9",
          2197 => x"08",
          2198 => x"08",
          2199 => x"38",
          2200 => x"77",
          2201 => x"84",
          2202 => x"39",
          2203 => x"52",
          2204 => x"eb",
          2205 => x"c8",
          2206 => x"53",
          2207 => x"08",
          2208 => x"c9",
          2209 => x"91",
          2210 => x"81",
          2211 => x"81",
          2212 => x"c8",
          2213 => x"b5",
          2214 => x"c8",
          2215 => x"51",
          2216 => x"81",
          2217 => x"c8",
          2218 => x"73",
          2219 => x"73",
          2220 => x"f2",
          2221 => x"d3",
          2222 => x"16",
          2223 => x"16",
          2224 => x"ff",
          2225 => x"05",
          2226 => x"80",
          2227 => x"d3",
          2228 => x"3d",
          2229 => x"3d",
          2230 => x"71",
          2231 => x"56",
          2232 => x"51",
          2233 => x"91",
          2234 => x"54",
          2235 => x"08",
          2236 => x"91",
          2237 => x"57",
          2238 => x"52",
          2239 => x"c8",
          2240 => x"c8",
          2241 => x"d3",
          2242 => x"c7",
          2243 => x"c8",
          2244 => x"08",
          2245 => x"54",
          2246 => x"e5",
          2247 => x"06",
          2248 => x"55",
          2249 => x"80",
          2250 => x"51",
          2251 => x"2e",
          2252 => x"17",
          2253 => x"2e",
          2254 => x"39",
          2255 => x"52",
          2256 => x"8a",
          2257 => x"c8",
          2258 => x"d3",
          2259 => x"2e",
          2260 => x"73",
          2261 => x"81",
          2262 => x"87",
          2263 => x"d3",
          2264 => x"3d",
          2265 => x"3d",
          2266 => x"11",
          2267 => x"aa",
          2268 => x"c8",
          2269 => x"ff",
          2270 => x"33",
          2271 => x"71",
          2272 => x"81",
          2273 => x"94",
          2274 => x"8e",
          2275 => x"c8",
          2276 => x"73",
          2277 => x"91",
          2278 => x"85",
          2279 => x"fc",
          2280 => x"79",
          2281 => x"ff",
          2282 => x"12",
          2283 => x"eb",
          2284 => x"70",
          2285 => x"72",
          2286 => x"81",
          2287 => x"73",
          2288 => x"94",
          2289 => x"94",
          2290 => x"0d",
          2291 => x"0d",
          2292 => x"56",
          2293 => x"5a",
          2294 => x"08",
          2295 => x"86",
          2296 => x"08",
          2297 => x"ed",
          2298 => x"d3",
          2299 => x"91",
          2300 => x"80",
          2301 => x"16",
          2302 => x"56",
          2303 => x"38",
          2304 => x"e2",
          2305 => x"08",
          2306 => x"70",
          2307 => x"81",
          2308 => x"51",
          2309 => x"86",
          2310 => x"81",
          2311 => x"30",
          2312 => x"70",
          2313 => x"06",
          2314 => x"51",
          2315 => x"73",
          2316 => x"38",
          2317 => x"96",
          2318 => x"df",
          2319 => x"72",
          2320 => x"81",
          2321 => x"81",
          2322 => x"2e",
          2323 => x"52",
          2324 => x"fa",
          2325 => x"c8",
          2326 => x"d3",
          2327 => x"38",
          2328 => x"fe",
          2329 => x"80",
          2330 => x"80",
          2331 => x"0c",
          2332 => x"c8",
          2333 => x"0d",
          2334 => x"0d",
          2335 => x"59",
          2336 => x"75",
          2337 => x"3f",
          2338 => x"08",
          2339 => x"c8",
          2340 => x"38",
          2341 => x"57",
          2342 => x"98",
          2343 => x"77",
          2344 => x"3f",
          2345 => x"08",
          2346 => x"c8",
          2347 => x"38",
          2348 => x"70",
          2349 => x"73",
          2350 => x"38",
          2351 => x"8b",
          2352 => x"06",
          2353 => x"86",
          2354 => x"15",
          2355 => x"2a",
          2356 => x"51",
          2357 => x"93",
          2358 => x"a0",
          2359 => x"51",
          2360 => x"91",
          2361 => x"80",
          2362 => x"80",
          2363 => x"f9",
          2364 => x"d3",
          2365 => x"91",
          2366 => x"80",
          2367 => x"38",
          2368 => x"91",
          2369 => x"8a",
          2370 => x"fb",
          2371 => x"70",
          2372 => x"81",
          2373 => x"fb",
          2374 => x"d3",
          2375 => x"91",
          2376 => x"b4",
          2377 => x"08",
          2378 => x"eb",
          2379 => x"d3",
          2380 => x"91",
          2381 => x"a0",
          2382 => x"91",
          2383 => x"52",
          2384 => x"51",
          2385 => x"8b",
          2386 => x"52",
          2387 => x"51",
          2388 => x"81",
          2389 => x"34",
          2390 => x"c8",
          2391 => x"0d",
          2392 => x"0d",
          2393 => x"98",
          2394 => x"70",
          2395 => x"ea",
          2396 => x"d3",
          2397 => x"91",
          2398 => x"8d",
          2399 => x"08",
          2400 => x"34",
          2401 => x"16",
          2402 => x"d3",
          2403 => x"3d",
          2404 => x"3d",
          2405 => x"57",
          2406 => x"89",
          2407 => x"17",
          2408 => x"81",
          2409 => x"70",
          2410 => x"17",
          2411 => x"33",
          2412 => x"54",
          2413 => x"2e",
          2414 => x"85",
          2415 => x"06",
          2416 => x"e5",
          2417 => x"2e",
          2418 => x"8e",
          2419 => x"88",
          2420 => x"0b",
          2421 => x"81",
          2422 => x"15",
          2423 => x"72",
          2424 => x"81",
          2425 => x"74",
          2426 => x"75",
          2427 => x"52",
          2428 => x"13",
          2429 => x"08",
          2430 => x"33",
          2431 => x"9c",
          2432 => x"05",
          2433 => x"3f",
          2434 => x"08",
          2435 => x"17",
          2436 => x"51",
          2437 => x"91",
          2438 => x"86",
          2439 => x"17",
          2440 => x"51",
          2441 => x"91",
          2442 => x"84",
          2443 => x"3d",
          2444 => x"3d",
          2445 => x"08",
          2446 => x"5d",
          2447 => x"53",
          2448 => x"51",
          2449 => x"80",
          2450 => x"88",
          2451 => x"5a",
          2452 => x"09",
          2453 => x"df",
          2454 => x"70",
          2455 => x"71",
          2456 => x"30",
          2457 => x"73",
          2458 => x"51",
          2459 => x"57",
          2460 => x"38",
          2461 => x"75",
          2462 => x"18",
          2463 => x"75",
          2464 => x"30",
          2465 => x"32",
          2466 => x"73",
          2467 => x"53",
          2468 => x"55",
          2469 => x"89",
          2470 => x"75",
          2471 => x"e4",
          2472 => x"7c",
          2473 => x"a0",
          2474 => x"38",
          2475 => x"8b",
          2476 => x"54",
          2477 => x"78",
          2478 => x"81",
          2479 => x"54",
          2480 => x"82",
          2481 => x"af",
          2482 => x"77",
          2483 => x"70",
          2484 => x"25",
          2485 => x"07",
          2486 => x"51",
          2487 => x"2e",
          2488 => x"39",
          2489 => x"80",
          2490 => x"33",
          2491 => x"73",
          2492 => x"81",
          2493 => x"81",
          2494 => x"1a",
          2495 => x"55",
          2496 => x"dc",
          2497 => x"06",
          2498 => x"55",
          2499 => x"54",
          2500 => x"81",
          2501 => x"ae",
          2502 => x"70",
          2503 => x"7d",
          2504 => x"51",
          2505 => x"2e",
          2506 => x"8b",
          2507 => x"77",
          2508 => x"30",
          2509 => x"71",
          2510 => x"53",
          2511 => x"55",
          2512 => x"38",
          2513 => x"5a",
          2514 => x"75",
          2515 => x"73",
          2516 => x"38",
          2517 => x"06",
          2518 => x"11",
          2519 => x"75",
          2520 => x"3f",
          2521 => x"08",
          2522 => x"38",
          2523 => x"33",
          2524 => x"54",
          2525 => x"e5",
          2526 => x"d3",
          2527 => x"2e",
          2528 => x"1a",
          2529 => x"26",
          2530 => x"54",
          2531 => x"7a",
          2532 => x"74",
          2533 => x"7b",
          2534 => x"74",
          2535 => x"18",
          2536 => x"39",
          2537 => x"ba",
          2538 => x"ec",
          2539 => x"c8",
          2540 => x"38",
          2541 => x"54",
          2542 => x"89",
          2543 => x"70",
          2544 => x"57",
          2545 => x"54",
          2546 => x"81",
          2547 => x"e7",
          2548 => x"7c",
          2549 => x"77",
          2550 => x"38",
          2551 => x"73",
          2552 => x"09",
          2553 => x"38",
          2554 => x"84",
          2555 => x"27",
          2556 => x"39",
          2557 => x"39",
          2558 => x"39",
          2559 => x"8b",
          2560 => x"54",
          2561 => x"c8",
          2562 => x"0d",
          2563 => x"0d",
          2564 => x"58",
          2565 => x"70",
          2566 => x"55",
          2567 => x"83",
          2568 => x"80",
          2569 => x"51",
          2570 => x"80",
          2571 => x"38",
          2572 => x"74",
          2573 => x"80",
          2574 => x"94",
          2575 => x"17",
          2576 => x"81",
          2577 => x"7a",
          2578 => x"54",
          2579 => x"2e",
          2580 => x"83",
          2581 => x"80",
          2582 => x"51",
          2583 => x"80",
          2584 => x"81",
          2585 => x"81",
          2586 => x"07",
          2587 => x"38",
          2588 => x"17",
          2589 => x"33",
          2590 => x"9f",
          2591 => x"ff",
          2592 => x"17",
          2593 => x"75",
          2594 => x"3f",
          2595 => x"08",
          2596 => x"39",
          2597 => x"a5",
          2598 => x"84",
          2599 => x"51",
          2600 => x"91",
          2601 => x"55",
          2602 => x"08",
          2603 => x"75",
          2604 => x"3f",
          2605 => x"08",
          2606 => x"55",
          2607 => x"c8",
          2608 => x"80",
          2609 => x"d3",
          2610 => x"2e",
          2611 => x"80",
          2612 => x"85",
          2613 => x"06",
          2614 => x"80",
          2615 => x"73",
          2616 => x"81",
          2617 => x"72",
          2618 => x"ad",
          2619 => x"0b",
          2620 => x"80",
          2621 => x"39",
          2622 => x"70",
          2623 => x"53",
          2624 => x"85",
          2625 => x"73",
          2626 => x"81",
          2627 => x"72",
          2628 => x"16",
          2629 => x"2a",
          2630 => x"51",
          2631 => x"80",
          2632 => x"38",
          2633 => x"83",
          2634 => x"b4",
          2635 => x"51",
          2636 => x"91",
          2637 => x"88",
          2638 => x"dd",
          2639 => x"d3",
          2640 => x"3d",
          2641 => x"3d",
          2642 => x"ff",
          2643 => x"72",
          2644 => x"5a",
          2645 => x"81",
          2646 => x"70",
          2647 => x"33",
          2648 => x"70",
          2649 => x"26",
          2650 => x"06",
          2651 => x"53",
          2652 => x"72",
          2653 => x"81",
          2654 => x"38",
          2655 => x"11",
          2656 => x"89",
          2657 => x"82",
          2658 => x"ff",
          2659 => x"51",
          2660 => x"77",
          2661 => x"38",
          2662 => x"bb",
          2663 => x"77",
          2664 => x"70",
          2665 => x"57",
          2666 => x"70",
          2667 => x"33",
          2668 => x"05",
          2669 => x"9f",
          2670 => x"54",
          2671 => x"89",
          2672 => x"70",
          2673 => x"55",
          2674 => x"13",
          2675 => x"26",
          2676 => x"13",
          2677 => x"06",
          2678 => x"30",
          2679 => x"70",
          2680 => x"07",
          2681 => x"9f",
          2682 => x"55",
          2683 => x"ff",
          2684 => x"30",
          2685 => x"70",
          2686 => x"07",
          2687 => x"9f",
          2688 => x"55",
          2689 => x"80",
          2690 => x"81",
          2691 => x"78",
          2692 => x"38",
          2693 => x"83",
          2694 => x"77",
          2695 => x"5a",
          2696 => x"39",
          2697 => x"33",
          2698 => x"d3",
          2699 => x"3d",
          2700 => x"3d",
          2701 => x"80",
          2702 => x"34",
          2703 => x"17",
          2704 => x"75",
          2705 => x"3f",
          2706 => x"d3",
          2707 => x"84",
          2708 => x"16",
          2709 => x"3f",
          2710 => x"08",
          2711 => x"06",
          2712 => x"73",
          2713 => x"2e",
          2714 => x"80",
          2715 => x"0b",
          2716 => x"55",
          2717 => x"e9",
          2718 => x"06",
          2719 => x"55",
          2720 => x"32",
          2721 => x"80",
          2722 => x"51",
          2723 => x"8e",
          2724 => x"33",
          2725 => x"e8",
          2726 => x"06",
          2727 => x"53",
          2728 => x"52",
          2729 => x"51",
          2730 => x"91",
          2731 => x"55",
          2732 => x"08",
          2733 => x"38",
          2734 => x"bb",
          2735 => x"86",
          2736 => x"a3",
          2737 => x"c8",
          2738 => x"d3",
          2739 => x"2e",
          2740 => x"55",
          2741 => x"c8",
          2742 => x"0d",
          2743 => x"0d",
          2744 => x"05",
          2745 => x"33",
          2746 => x"74",
          2747 => x"fc",
          2748 => x"d3",
          2749 => x"8b",
          2750 => x"91",
          2751 => x"24",
          2752 => x"91",
          2753 => x"10",
          2754 => x"e4",
          2755 => x"56",
          2756 => x"74",
          2757 => x"88",
          2758 => x"0c",
          2759 => x"06",
          2760 => x"57",
          2761 => x"af",
          2762 => x"33",
          2763 => x"3f",
          2764 => x"08",
          2765 => x"70",
          2766 => x"54",
          2767 => x"76",
          2768 => x"38",
          2769 => x"70",
          2770 => x"53",
          2771 => x"86",
          2772 => x"56",
          2773 => x"80",
          2774 => x"81",
          2775 => x"52",
          2776 => x"51",
          2777 => x"91",
          2778 => x"81",
          2779 => x"81",
          2780 => x"83",
          2781 => x"a8",
          2782 => x"2e",
          2783 => x"82",
          2784 => x"06",
          2785 => x"56",
          2786 => x"38",
          2787 => x"75",
          2788 => x"9e",
          2789 => x"c8",
          2790 => x"06",
          2791 => x"2e",
          2792 => x"80",
          2793 => x"54",
          2794 => x"15",
          2795 => x"10",
          2796 => x"05",
          2797 => x"33",
          2798 => x"80",
          2799 => x"2e",
          2800 => x"fa",
          2801 => x"eb",
          2802 => x"c8",
          2803 => x"78",
          2804 => x"54",
          2805 => x"d0",
          2806 => x"8f",
          2807 => x"10",
          2808 => x"08",
          2809 => x"57",
          2810 => x"90",
          2811 => x"74",
          2812 => x"3f",
          2813 => x"08",
          2814 => x"57",
          2815 => x"89",
          2816 => x"54",
          2817 => x"d3",
          2818 => x"76",
          2819 => x"90",
          2820 => x"76",
          2821 => x"88",
          2822 => x"51",
          2823 => x"91",
          2824 => x"83",
          2825 => x"53",
          2826 => x"84",
          2827 => x"81",
          2828 => x"38",
          2829 => x"51",
          2830 => x"91",
          2831 => x"83",
          2832 => x"54",
          2833 => x"80",
          2834 => x"d9",
          2835 => x"d3",
          2836 => x"73",
          2837 => x"80",
          2838 => x"82",
          2839 => x"c4",
          2840 => x"05",
          2841 => x"72",
          2842 => x"b4",
          2843 => x"33",
          2844 => x"80",
          2845 => x"52",
          2846 => x"8a",
          2847 => x"83",
          2848 => x"53",
          2849 => x"8b",
          2850 => x"73",
          2851 => x"80",
          2852 => x"8d",
          2853 => x"39",
          2854 => x"51",
          2855 => x"91",
          2856 => x"88",
          2857 => x"d3",
          2858 => x"ff",
          2859 => x"06",
          2860 => x"72",
          2861 => x"80",
          2862 => x"d8",
          2863 => x"d3",
          2864 => x"ff",
          2865 => x"72",
          2866 => x"d4",
          2867 => x"e3",
          2868 => x"c8",
          2869 => x"c2",
          2870 => x"be",
          2871 => x"c8",
          2872 => x"ff",
          2873 => x"56",
          2874 => x"83",
          2875 => x"15",
          2876 => x"71",
          2877 => x"59",
          2878 => x"77",
          2879 => x"a0",
          2880 => x"22",
          2881 => x"31",
          2882 => x"ab",
          2883 => x"c8",
          2884 => x"56",
          2885 => x"08",
          2886 => x"84",
          2887 => x"91",
          2888 => x"80",
          2889 => x"f5",
          2890 => x"83",
          2891 => x"ff",
          2892 => x"38",
          2893 => x"9f",
          2894 => x"38",
          2895 => x"56",
          2896 => x"82",
          2897 => x"13",
          2898 => x"79",
          2899 => x"79",
          2900 => x"0c",
          2901 => x"16",
          2902 => x"2e",
          2903 => x"b7",
          2904 => x"15",
          2905 => x"3f",
          2906 => x"08",
          2907 => x"06",
          2908 => x"72",
          2909 => x"88",
          2910 => x"8d",
          2911 => x"a0",
          2912 => x"15",
          2913 => x"3f",
          2914 => x"08",
          2915 => x"98",
          2916 => x"2b",
          2917 => x"88",
          2918 => x"8d",
          2919 => x"2e",
          2920 => x"a4",
          2921 => x"a8",
          2922 => x"82",
          2923 => x"06",
          2924 => x"15",
          2925 => x"94",
          2926 => x"08",
          2927 => x"08",
          2928 => x"2a",
          2929 => x"81",
          2930 => x"53",
          2931 => x"89",
          2932 => x"56",
          2933 => x"08",
          2934 => x"38",
          2935 => x"16",
          2936 => x"8c",
          2937 => x"80",
          2938 => x"34",
          2939 => x"09",
          2940 => x"92",
          2941 => x"15",
          2942 => x"3f",
          2943 => x"08",
          2944 => x"06",
          2945 => x"2e",
          2946 => x"80",
          2947 => x"1a",
          2948 => x"d9",
          2949 => x"d3",
          2950 => x"ea",
          2951 => x"c8",
          2952 => x"34",
          2953 => x"51",
          2954 => x"91",
          2955 => x"83",
          2956 => x"53",
          2957 => x"d5",
          2958 => x"06",
          2959 => x"b4",
          2960 => x"ef",
          2961 => x"c8",
          2962 => x"85",
          2963 => x"09",
          2964 => x"38",
          2965 => x"51",
          2966 => x"91",
          2967 => x"86",
          2968 => x"f2",
          2969 => x"06",
          2970 => x"9c",
          2971 => x"c3",
          2972 => x"c8",
          2973 => x"0c",
          2974 => x"51",
          2975 => x"91",
          2976 => x"8c",
          2977 => x"75",
          2978 => x"f4",
          2979 => x"53",
          2980 => x"f4",
          2981 => x"16",
          2982 => x"94",
          2983 => x"56",
          2984 => x"c8",
          2985 => x"0d",
          2986 => x"0d",
          2987 => x"55",
          2988 => x"b5",
          2989 => x"80",
          2990 => x"73",
          2991 => x"53",
          2992 => x"2e",
          2993 => x"14",
          2994 => x"22",
          2995 => x"76",
          2996 => x"06",
          2997 => x"13",
          2998 => x"f9",
          2999 => x"c8",
          3000 => x"52",
          3001 => x"71",
          3002 => x"74",
          3003 => x"81",
          3004 => x"73",
          3005 => x"73",
          3006 => x"74",
          3007 => x"0c",
          3008 => x"04",
          3009 => x"02",
          3010 => x"7a",
          3011 => x"fc",
          3012 => x"f4",
          3013 => x"d3",
          3014 => x"8b",
          3015 => x"91",
          3016 => x"24",
          3017 => x"91",
          3018 => x"10",
          3019 => x"e4",
          3020 => x"51",
          3021 => x"2e",
          3022 => x"74",
          3023 => x"2e",
          3024 => x"54",
          3025 => x"74",
          3026 => x"d3",
          3027 => x"71",
          3028 => x"54",
          3029 => x"92",
          3030 => x"89",
          3031 => x"84",
          3032 => x"f9",
          3033 => x"c8",
          3034 => x"91",
          3035 => x"88",
          3036 => x"eb",
          3037 => x"02",
          3038 => x"e7",
          3039 => x"58",
          3040 => x"80",
          3041 => x"38",
          3042 => x"70",
          3043 => x"d0",
          3044 => x"3d",
          3045 => x"57",
          3046 => x"91",
          3047 => x"56",
          3048 => x"08",
          3049 => x"7a",
          3050 => x"97",
          3051 => x"51",
          3052 => x"91",
          3053 => x"56",
          3054 => x"08",
          3055 => x"80",
          3056 => x"70",
          3057 => x"59",
          3058 => x"83",
          3059 => x"76",
          3060 => x"74",
          3061 => x"c3",
          3062 => x"2e",
          3063 => x"84",
          3064 => x"06",
          3065 => x"3d",
          3066 => x"ea",
          3067 => x"d3",
          3068 => x"76",
          3069 => x"a0",
          3070 => x"05",
          3071 => x"55",
          3072 => x"85",
          3073 => x"90",
          3074 => x"2a",
          3075 => x"51",
          3076 => x"2e",
          3077 => x"56",
          3078 => x"38",
          3079 => x"70",
          3080 => x"55",
          3081 => x"81",
          3082 => x"52",
          3083 => x"b6",
          3084 => x"c8",
          3085 => x"88",
          3086 => x"62",
          3087 => x"d2",
          3088 => x"55",
          3089 => x"16",
          3090 => x"62",
          3091 => x"e6",
          3092 => x"52",
          3093 => x"51",
          3094 => x"7a",
          3095 => x"83",
          3096 => x"80",
          3097 => x"38",
          3098 => x"08",
          3099 => x"54",
          3100 => x"05",
          3101 => x"db",
          3102 => x"d3",
          3103 => x"91",
          3104 => x"82",
          3105 => x"52",
          3106 => x"bc",
          3107 => x"c8",
          3108 => x"1b",
          3109 => x"56",
          3110 => x"75",
          3111 => x"02",
          3112 => x"70",
          3113 => x"81",
          3114 => x"59",
          3115 => x"85",
          3116 => x"9c",
          3117 => x"2a",
          3118 => x"51",
          3119 => x"2e",
          3120 => x"b2",
          3121 => x"06",
          3122 => x"2e",
          3123 => x"56",
          3124 => x"38",
          3125 => x"70",
          3126 => x"55",
          3127 => x"86",
          3128 => x"c0",
          3129 => x"b0",
          3130 => x"1a",
          3131 => x"1a",
          3132 => x"81",
          3133 => x"52",
          3134 => x"ea",
          3135 => x"c8",
          3136 => x"0c",
          3137 => x"51",
          3138 => x"91",
          3139 => x"8c",
          3140 => x"78",
          3141 => x"22",
          3142 => x"76",
          3143 => x"75",
          3144 => x"75",
          3145 => x"75",
          3146 => x"84",
          3147 => x"52",
          3148 => x"d1",
          3149 => x"85",
          3150 => x"06",
          3151 => x"80",
          3152 => x"38",
          3153 => x"80",
          3154 => x"38",
          3155 => x"94",
          3156 => x"8a",
          3157 => x"89",
          3158 => x"08",
          3159 => x"5d",
          3160 => x"55",
          3161 => x"52",
          3162 => x"fc",
          3163 => x"c8",
          3164 => x"d3",
          3165 => x"26",
          3166 => x"56",
          3167 => x"09",
          3168 => x"38",
          3169 => x"7a",
          3170 => x"30",
          3171 => x"80",
          3172 => x"7d",
          3173 => x"51",
          3174 => x"38",
          3175 => x"0c",
          3176 => x"38",
          3177 => x"06",
          3178 => x"2e",
          3179 => x"52",
          3180 => x"8a",
          3181 => x"c8",
          3182 => x"82",
          3183 => x"78",
          3184 => x"d3",
          3185 => x"70",
          3186 => x"55",
          3187 => x"53",
          3188 => x"7a",
          3189 => x"52",
          3190 => x"3f",
          3191 => x"08",
          3192 => x"38",
          3193 => x"80",
          3194 => x"80",
          3195 => x"55",
          3196 => x"c8",
          3197 => x"0d",
          3198 => x"0d",
          3199 => x"63",
          3200 => x"57",
          3201 => x"8f",
          3202 => x"52",
          3203 => x"99",
          3204 => x"c8",
          3205 => x"d3",
          3206 => x"38",
          3207 => x"55",
          3208 => x"86",
          3209 => x"83",
          3210 => x"17",
          3211 => x"55",
          3212 => x"80",
          3213 => x"38",
          3214 => x"0b",
          3215 => x"82",
          3216 => x"39",
          3217 => x"18",
          3218 => x"83",
          3219 => x"0b",
          3220 => x"82",
          3221 => x"39",
          3222 => x"18",
          3223 => x"82",
          3224 => x"0b",
          3225 => x"81",
          3226 => x"39",
          3227 => x"18",
          3228 => x"82",
          3229 => x"17",
          3230 => x"08",
          3231 => x"79",
          3232 => x"74",
          3233 => x"2e",
          3234 => x"94",
          3235 => x"83",
          3236 => x"56",
          3237 => x"38",
          3238 => x"22",
          3239 => x"89",
          3240 => x"55",
          3241 => x"75",
          3242 => x"17",
          3243 => x"39",
          3244 => x"52",
          3245 => x"b0",
          3246 => x"c8",
          3247 => x"75",
          3248 => x"38",
          3249 => x"fe",
          3250 => x"98",
          3251 => x"17",
          3252 => x"51",
          3253 => x"91",
          3254 => x"80",
          3255 => x"38",
          3256 => x"08",
          3257 => x"2a",
          3258 => x"80",
          3259 => x"38",
          3260 => x"8a",
          3261 => x"56",
          3262 => x"27",
          3263 => x"7b",
          3264 => x"54",
          3265 => x"52",
          3266 => x"33",
          3267 => x"ef",
          3268 => x"c8",
          3269 => x"38",
          3270 => x"70",
          3271 => x"56",
          3272 => x"9b",
          3273 => x"08",
          3274 => x"74",
          3275 => x"38",
          3276 => x"a8",
          3277 => x"84",
          3278 => x"51",
          3279 => x"79",
          3280 => x"80",
          3281 => x"17",
          3282 => x"80",
          3283 => x"17",
          3284 => x"2b",
          3285 => x"80",
          3286 => x"81",
          3287 => x"08",
          3288 => x"52",
          3289 => x"33",
          3290 => x"ec",
          3291 => x"c8",
          3292 => x"38",
          3293 => x"80",
          3294 => x"74",
          3295 => x"81",
          3296 => x"a8",
          3297 => x"81",
          3298 => x"55",
          3299 => x"91",
          3300 => x"fd",
          3301 => x"9c",
          3302 => x"17",
          3303 => x"06",
          3304 => x"31",
          3305 => x"76",
          3306 => x"78",
          3307 => x"94",
          3308 => x"ff",
          3309 => x"05",
          3310 => x"cb",
          3311 => x"76",
          3312 => x"17",
          3313 => x"1d",
          3314 => x"18",
          3315 => x"5d",
          3316 => x"b7",
          3317 => x"75",
          3318 => x"0c",
          3319 => x"04",
          3320 => x"7f",
          3321 => x"5f",
          3322 => x"80",
          3323 => x"3d",
          3324 => x"76",
          3325 => x"3f",
          3326 => x"08",
          3327 => x"c8",
          3328 => x"91",
          3329 => x"74",
          3330 => x"38",
          3331 => x"82",
          3332 => x"33",
          3333 => x"70",
          3334 => x"56",
          3335 => x"74",
          3336 => x"ee",
          3337 => x"82",
          3338 => x"34",
          3339 => x"e2",
          3340 => x"91",
          3341 => x"56",
          3342 => x"81",
          3343 => x"34",
          3344 => x"ce",
          3345 => x"91",
          3346 => x"56",
          3347 => x"81",
          3348 => x"34",
          3349 => x"ba",
          3350 => x"91",
          3351 => x"56",
          3352 => x"94",
          3353 => x"55",
          3354 => x"08",
          3355 => x"94",
          3356 => x"59",
          3357 => x"83",
          3358 => x"17",
          3359 => x"ff",
          3360 => x"74",
          3361 => x"7d",
          3362 => x"ff",
          3363 => x"2a",
          3364 => x"7a",
          3365 => x"75",
          3366 => x"17",
          3367 => x"a3",
          3368 => x"76",
          3369 => x"3f",
          3370 => x"08",
          3371 => x"98",
          3372 => x"76",
          3373 => x"3f",
          3374 => x"08",
          3375 => x"2e",
          3376 => x"74",
          3377 => x"df",
          3378 => x"2e",
          3379 => x"74",
          3380 => x"88",
          3381 => x"38",
          3382 => x"0c",
          3383 => x"70",
          3384 => x"58",
          3385 => x"a5",
          3386 => x"9c",
          3387 => x"a8",
          3388 => x"81",
          3389 => x"55",
          3390 => x"91",
          3391 => x"fe",
          3392 => x"17",
          3393 => x"06",
          3394 => x"18",
          3395 => x"08",
          3396 => x"cd",
          3397 => x"d3",
          3398 => x"2e",
          3399 => x"91",
          3400 => x"1b",
          3401 => x"5b",
          3402 => x"2e",
          3403 => x"79",
          3404 => x"11",
          3405 => x"56",
          3406 => x"85",
          3407 => x"31",
          3408 => x"77",
          3409 => x"7d",
          3410 => x"52",
          3411 => x"3f",
          3412 => x"08",
          3413 => x"9c",
          3414 => x"31",
          3415 => x"27",
          3416 => x"80",
          3417 => x"80",
          3418 => x"a8",
          3419 => x"b9",
          3420 => x"33",
          3421 => x"55",
          3422 => x"34",
          3423 => x"56",
          3424 => x"9c",
          3425 => x"2e",
          3426 => x"17",
          3427 => x"08",
          3428 => x"81",
          3429 => x"a8",
          3430 => x"81",
          3431 => x"55",
          3432 => x"91",
          3433 => x"fd",
          3434 => x"9c",
          3435 => x"17",
          3436 => x"06",
          3437 => x"31",
          3438 => x"76",
          3439 => x"78",
          3440 => x"7b",
          3441 => x"08",
          3442 => x"17",
          3443 => x"c7",
          3444 => x"17",
          3445 => x"07",
          3446 => x"18",
          3447 => x"31",
          3448 => x"7e",
          3449 => x"94",
          3450 => x"70",
          3451 => x"8c",
          3452 => x"58",
          3453 => x"76",
          3454 => x"75",
          3455 => x"18",
          3456 => x"f6",
          3457 => x"33",
          3458 => x"55",
          3459 => x"34",
          3460 => x"91",
          3461 => x"8f",
          3462 => x"f7",
          3463 => x"8c",
          3464 => x"53",
          3465 => x"f1",
          3466 => x"d3",
          3467 => x"91",
          3468 => x"81",
          3469 => x"18",
          3470 => x"2a",
          3471 => x"51",
          3472 => x"80",
          3473 => x"38",
          3474 => x"55",
          3475 => x"a7",
          3476 => x"9c",
          3477 => x"a8",
          3478 => x"81",
          3479 => x"55",
          3480 => x"81",
          3481 => x"c8",
          3482 => x"38",
          3483 => x"80",
          3484 => x"74",
          3485 => x"a0",
          3486 => x"79",
          3487 => x"3f",
          3488 => x"08",
          3489 => x"c8",
          3490 => x"38",
          3491 => x"8b",
          3492 => x"07",
          3493 => x"8b",
          3494 => x"18",
          3495 => x"52",
          3496 => x"d9",
          3497 => x"18",
          3498 => x"16",
          3499 => x"3f",
          3500 => x"0a",
          3501 => x"51",
          3502 => x"76",
          3503 => x"51",
          3504 => x"79",
          3505 => x"83",
          3506 => x"51",
          3507 => x"91",
          3508 => x"90",
          3509 => x"bf",
          3510 => x"74",
          3511 => x"76",
          3512 => x"d3",
          3513 => x"3d",
          3514 => x"3d",
          3515 => x"52",
          3516 => x"3f",
          3517 => x"08",
          3518 => x"c8",
          3519 => x"86",
          3520 => x"52",
          3521 => x"a1",
          3522 => x"c8",
          3523 => x"d3",
          3524 => x"38",
          3525 => x"08",
          3526 => x"91",
          3527 => x"86",
          3528 => x"fe",
          3529 => x"3d",
          3530 => x"3f",
          3531 => x"0b",
          3532 => x"08",
          3533 => x"91",
          3534 => x"91",
          3535 => x"80",
          3536 => x"d3",
          3537 => x"3d",
          3538 => x"3d",
          3539 => x"93",
          3540 => x"52",
          3541 => x"e7",
          3542 => x"d3",
          3543 => x"91",
          3544 => x"80",
          3545 => x"58",
          3546 => x"3d",
          3547 => x"e1",
          3548 => x"d3",
          3549 => x"91",
          3550 => x"be",
          3551 => x"c7",
          3552 => x"98",
          3553 => x"73",
          3554 => x"38",
          3555 => x"12",
          3556 => x"39",
          3557 => x"33",
          3558 => x"70",
          3559 => x"55",
          3560 => x"2e",
          3561 => x"7f",
          3562 => x"54",
          3563 => x"91",
          3564 => x"94",
          3565 => x"39",
          3566 => x"84",
          3567 => x"06",
          3568 => x"55",
          3569 => x"c8",
          3570 => x"0d",
          3571 => x"0d",
          3572 => x"a3",
          3573 => x"5c",
          3574 => x"80",
          3575 => x"ff",
          3576 => x"a2",
          3577 => x"f5",
          3578 => x"c8",
          3579 => x"d3",
          3580 => x"93",
          3581 => x"7b",
          3582 => x"08",
          3583 => x"56",
          3584 => x"2e",
          3585 => x"96",
          3586 => x"3d",
          3587 => x"a0",
          3588 => x"d1",
          3589 => x"d3",
          3590 => x"91",
          3591 => x"81",
          3592 => x"52",
          3593 => x"a0",
          3594 => x"c8",
          3595 => x"d3",
          3596 => x"cb",
          3597 => x"7e",
          3598 => x"3f",
          3599 => x"08",
          3600 => x"7a",
          3601 => x"3f",
          3602 => x"08",
          3603 => x"c8",
          3604 => x"38",
          3605 => x"52",
          3606 => x"f1",
          3607 => x"c8",
          3608 => x"d3",
          3609 => x"38",
          3610 => x"51",
          3611 => x"91",
          3612 => x"75",
          3613 => x"76",
          3614 => x"d2",
          3615 => x"d3",
          3616 => x"91",
          3617 => x"80",
          3618 => x"76",
          3619 => x"81",
          3620 => x"82",
          3621 => x"ef",
          3622 => x"ff",
          3623 => x"d4",
          3624 => x"ee",
          3625 => x"3d",
          3626 => x"81",
          3627 => x"52",
          3628 => x"73",
          3629 => x"38",
          3630 => x"16",
          3631 => x"51",
          3632 => x"f4",
          3633 => x"54",
          3634 => x"85",
          3635 => x"af",
          3636 => x"2e",
          3637 => x"58",
          3638 => x"3d",
          3639 => x"18",
          3640 => x"58",
          3641 => x"14",
          3642 => x"75",
          3643 => x"19",
          3644 => x"11",
          3645 => x"74",
          3646 => x"74",
          3647 => x"76",
          3648 => x"78",
          3649 => x"81",
          3650 => x"ff",
          3651 => x"08",
          3652 => x"af",
          3653 => x"70",
          3654 => x"33",
          3655 => x"91",
          3656 => x"70",
          3657 => x"52",
          3658 => x"57",
          3659 => x"2e",
          3660 => x"16",
          3661 => x"33",
          3662 => x"73",
          3663 => x"16",
          3664 => x"26",
          3665 => x"58",
          3666 => x"94",
          3667 => x"54",
          3668 => x"70",
          3669 => x"34",
          3670 => x"75",
          3671 => x"38",
          3672 => x"81",
          3673 => x"81",
          3674 => x"83",
          3675 => x"76",
          3676 => x"3d",
          3677 => x"1a",
          3678 => x"33",
          3679 => x"05",
          3680 => x"79",
          3681 => x"80",
          3682 => x"91",
          3683 => x"a1",
          3684 => x"f4",
          3685 => x"60",
          3686 => x"05",
          3687 => x"59",
          3688 => x"3f",
          3689 => x"08",
          3690 => x"c8",
          3691 => x"91",
          3692 => x"79",
          3693 => x"38",
          3694 => x"f9",
          3695 => x"08",
          3696 => x"38",
          3697 => x"70",
          3698 => x"81",
          3699 => x"56",
          3700 => x"8c",
          3701 => x"94",
          3702 => x"80",
          3703 => x"0c",
          3704 => x"2e",
          3705 => x"7c",
          3706 => x"70",
          3707 => x"51",
          3708 => x"2e",
          3709 => x"52",
          3710 => x"ff",
          3711 => x"91",
          3712 => x"ff",
          3713 => x"70",
          3714 => x"ff",
          3715 => x"91",
          3716 => x"75",
          3717 => x"78",
          3718 => x"94",
          3719 => x"94",
          3720 => x"98",
          3721 => x"58",
          3722 => x"88",
          3723 => x"75",
          3724 => x"52",
          3725 => x"a7",
          3726 => x"c8",
          3727 => x"d3",
          3728 => x"2e",
          3729 => x"8b",
          3730 => x"91",
          3731 => x"55",
          3732 => x"91",
          3733 => x"ff",
          3734 => x"06",
          3735 => x"0b",
          3736 => x"81",
          3737 => x"39",
          3738 => x"08",
          3739 => x"75",
          3740 => x"75",
          3741 => x"a1",
          3742 => x"27",
          3743 => x"77",
          3744 => x"18",
          3745 => x"19",
          3746 => x"33",
          3747 => x"70",
          3748 => x"57",
          3749 => x"80",
          3750 => x"75",
          3751 => x"c8",
          3752 => x"d3",
          3753 => x"91",
          3754 => x"94",
          3755 => x"c8",
          3756 => x"39",
          3757 => x"51",
          3758 => x"91",
          3759 => x"56",
          3760 => x"81",
          3761 => x"76",
          3762 => x"7c",
          3763 => x"08",
          3764 => x"38",
          3765 => x"18",
          3766 => x"81",
          3767 => x"98",
          3768 => x"79",
          3769 => x"38",
          3770 => x"18",
          3771 => x"77",
          3772 => x"55",
          3773 => x"a1",
          3774 => x"7c",
          3775 => x"3f",
          3776 => x"08",
          3777 => x"0b",
          3778 => x"82",
          3779 => x"39",
          3780 => x"91",
          3781 => x"05",
          3782 => x"08",
          3783 => x"27",
          3784 => x"17",
          3785 => x"0c",
          3786 => x"80",
          3787 => x"74",
          3788 => x"94",
          3789 => x"ff",
          3790 => x"80",
          3791 => x"38",
          3792 => x"7b",
          3793 => x"38",
          3794 => x"70",
          3795 => x"5c",
          3796 => x"b0",
          3797 => x"9c",
          3798 => x"a8",
          3799 => x"81",
          3800 => x"55",
          3801 => x"3f",
          3802 => x"08",
          3803 => x"38",
          3804 => x"18",
          3805 => x"bd",
          3806 => x"33",
          3807 => x"55",
          3808 => x"34",
          3809 => x"53",
          3810 => x"7c",
          3811 => x"52",
          3812 => x"eb",
          3813 => x"c8",
          3814 => x"93",
          3815 => x"91",
          3816 => x"55",
          3817 => x"0b",
          3818 => x"81",
          3819 => x"7a",
          3820 => x"79",
          3821 => x"d3",
          3822 => x"3d",
          3823 => x"3d",
          3824 => x"89",
          3825 => x"2e",
          3826 => x"80",
          3827 => x"fc",
          3828 => x"3d",
          3829 => x"de",
          3830 => x"d3",
          3831 => x"91",
          3832 => x"80",
          3833 => x"76",
          3834 => x"75",
          3835 => x"3f",
          3836 => x"08",
          3837 => x"c8",
          3838 => x"38",
          3839 => x"70",
          3840 => x"57",
          3841 => x"a6",
          3842 => x"33",
          3843 => x"70",
          3844 => x"55",
          3845 => x"2e",
          3846 => x"16",
          3847 => x"51",
          3848 => x"91",
          3849 => x"88",
          3850 => x"39",
          3851 => x"95",
          3852 => x"86",
          3853 => x"17",
          3854 => x"75",
          3855 => x"3f",
          3856 => x"08",
          3857 => x"2e",
          3858 => x"83",
          3859 => x"74",
          3860 => x"38",
          3861 => x"74",
          3862 => x"d3",
          3863 => x"3d",
          3864 => x"3d",
          3865 => x"3d",
          3866 => x"70",
          3867 => x"b9",
          3868 => x"c8",
          3869 => x"d3",
          3870 => x"38",
          3871 => x"08",
          3872 => x"91",
          3873 => x"86",
          3874 => x"fb",
          3875 => x"79",
          3876 => x"05",
          3877 => x"56",
          3878 => x"3f",
          3879 => x"08",
          3880 => x"c8",
          3881 => x"38",
          3882 => x"91",
          3883 => x"52",
          3884 => x"c5",
          3885 => x"c8",
          3886 => x"39",
          3887 => x"51",
          3888 => x"91",
          3889 => x"53",
          3890 => x"08",
          3891 => x"81",
          3892 => x"80",
          3893 => x"38",
          3894 => x"51",
          3895 => x"72",
          3896 => x"c9",
          3897 => x"d3",
          3898 => x"91",
          3899 => x"84",
          3900 => x"06",
          3901 => x"53",
          3902 => x"c8",
          3903 => x"0d",
          3904 => x"0d",
          3905 => x"53",
          3906 => x"53",
          3907 => x"54",
          3908 => x"91",
          3909 => x"55",
          3910 => x"08",
          3911 => x"52",
          3912 => x"e9",
          3913 => x"c8",
          3914 => x"d3",
          3915 => x"38",
          3916 => x"05",
          3917 => x"2b",
          3918 => x"80",
          3919 => x"86",
          3920 => x"75",
          3921 => x"38",
          3922 => x"3d",
          3923 => x"d0",
          3924 => x"91",
          3925 => x"93",
          3926 => x"f2",
          3927 => x"63",
          3928 => x"53",
          3929 => x"05",
          3930 => x"51",
          3931 => x"91",
          3932 => x"59",
          3933 => x"08",
          3934 => x"7a",
          3935 => x"08",
          3936 => x"fe",
          3937 => x"90",
          3938 => x"26",
          3939 => x"15",
          3940 => x"81",
          3941 => x"59",
          3942 => x"82",
          3943 => x"39",
          3944 => x"33",
          3945 => x"73",
          3946 => x"81",
          3947 => x"38",
          3948 => x"56",
          3949 => x"3d",
          3950 => x"ff",
          3951 => x"91",
          3952 => x"ff",
          3953 => x"91",
          3954 => x"81",
          3955 => x"91",
          3956 => x"30",
          3957 => x"c8",
          3958 => x"25",
          3959 => x"18",
          3960 => x"58",
          3961 => x"08",
          3962 => x"38",
          3963 => x"7a",
          3964 => x"a4",
          3965 => x"57",
          3966 => x"74",
          3967 => x"52",
          3968 => x"52",
          3969 => x"c0",
          3970 => x"c8",
          3971 => x"d3",
          3972 => x"d5",
          3973 => x"33",
          3974 => x"82",
          3975 => x"06",
          3976 => x"15",
          3977 => x"ff",
          3978 => x"91",
          3979 => x"83",
          3980 => x"70",
          3981 => x"25",
          3982 => x"58",
          3983 => x"9d",
          3984 => x"b4",
          3985 => x"b5",
          3986 => x"d3",
          3987 => x"0a",
          3988 => x"70",
          3989 => x"84",
          3990 => x"51",
          3991 => x"ff",
          3992 => x"57",
          3993 => x"93",
          3994 => x"0c",
          3995 => x"12",
          3996 => x"84",
          3997 => x"07",
          3998 => x"84",
          3999 => x"91",
          4000 => x"90",
          4001 => x"f8",
          4002 => x"8b",
          4003 => x"53",
          4004 => x"e0",
          4005 => x"d3",
          4006 => x"91",
          4007 => x"8a",
          4008 => x"33",
          4009 => x"2e",
          4010 => x"56",
          4011 => x"90",
          4012 => x"81",
          4013 => x"06",
          4014 => x"87",
          4015 => x"2e",
          4016 => x"94",
          4017 => x"19",
          4018 => x"bc",
          4019 => x"08",
          4020 => x"53",
          4021 => x"52",
          4022 => x"be",
          4023 => x"d3",
          4024 => x"80",
          4025 => x"0c",
          4026 => x"98",
          4027 => x"77",
          4028 => x"f4",
          4029 => x"c8",
          4030 => x"c8",
          4031 => x"70",
          4032 => x"07",
          4033 => x"57",
          4034 => x"d3",
          4035 => x"2e",
          4036 => x"83",
          4037 => x"76",
          4038 => x"55",
          4039 => x"08",
          4040 => x"98",
          4041 => x"75",
          4042 => x"ff",
          4043 => x"91",
          4044 => x"57",
          4045 => x"8c",
          4046 => x"18",
          4047 => x"07",
          4048 => x"19",
          4049 => x"38",
          4050 => x"55",
          4051 => x"ab",
          4052 => x"9c",
          4053 => x"a8",
          4054 => x"81",
          4055 => x"55",
          4056 => x"3f",
          4057 => x"08",
          4058 => x"38",
          4059 => x"39",
          4060 => x"80",
          4061 => x"74",
          4062 => x"76",
          4063 => x"38",
          4064 => x"34",
          4065 => x"39",
          4066 => x"91",
          4067 => x"8a",
          4068 => x"e3",
          4069 => x"bb",
          4070 => x"96",
          4071 => x"53",
          4072 => x"a4",
          4073 => x"3d",
          4074 => x"3f",
          4075 => x"08",
          4076 => x"c8",
          4077 => x"38",
          4078 => x"51",
          4079 => x"3f",
          4080 => x"52",
          4081 => x"05",
          4082 => x"3f",
          4083 => x"08",
          4084 => x"52",
          4085 => x"9a",
          4086 => x"ae",
          4087 => x"f7",
          4088 => x"85",
          4089 => x"06",
          4090 => x"73",
          4091 => x"38",
          4092 => x"82",
          4093 => x"bb",
          4094 => x"95",
          4095 => x"80",
          4096 => x"70",
          4097 => x"55",
          4098 => x"85",
          4099 => x"90",
          4100 => x"d2",
          4101 => x"06",
          4102 => x"2e",
          4103 => x"56",
          4104 => x"38",
          4105 => x"51",
          4106 => x"91",
          4107 => x"02",
          4108 => x"d2",
          4109 => x"84",
          4110 => x"06",
          4111 => x"57",
          4112 => x"80",
          4113 => x"bb",
          4114 => x"95",
          4115 => x"78",
          4116 => x"14",
          4117 => x"80",
          4118 => x"bb",
          4119 => x"95",
          4120 => x"59",
          4121 => x"bb",
          4122 => x"95",
          4123 => x"52",
          4124 => x"52",
          4125 => x"3f",
          4126 => x"08",
          4127 => x"c8",
          4128 => x"38",
          4129 => x"08",
          4130 => x"c6",
          4131 => x"d3",
          4132 => x"91",
          4133 => x"83",
          4134 => x"75",
          4135 => x"30",
          4136 => x"9f",
          4137 => x"58",
          4138 => x"80",
          4139 => x"bb",
          4140 => x"94",
          4141 => x"3d",
          4142 => x"c9",
          4143 => x"d3",
          4144 => x"d3",
          4145 => x"70",
          4146 => x"08",
          4147 => x"79",
          4148 => x"07",
          4149 => x"06",
          4150 => x"56",
          4151 => x"2e",
          4152 => x"bb",
          4153 => x"94",
          4154 => x"53",
          4155 => x"3d",
          4156 => x"ff",
          4157 => x"91",
          4158 => x"56",
          4159 => x"77",
          4160 => x"8b",
          4161 => x"c8",
          4162 => x"bb",
          4163 => x"93",
          4164 => x"91",
          4165 => x"9f",
          4166 => x"ea",
          4167 => x"53",
          4168 => x"05",
          4169 => x"51",
          4170 => x"91",
          4171 => x"55",
          4172 => x"08",
          4173 => x"77",
          4174 => x"98",
          4175 => x"51",
          4176 => x"91",
          4177 => x"55",
          4178 => x"08",
          4179 => x"55",
          4180 => x"09",
          4181 => x"93",
          4182 => x"db",
          4183 => x"85",
          4184 => x"06",
          4185 => x"73",
          4186 => x"38",
          4187 => x"84",
          4188 => x"06",
          4189 => x"77",
          4190 => x"98",
          4191 => x"51",
          4192 => x"3f",
          4193 => x"08",
          4194 => x"91",
          4195 => x"75",
          4196 => x"06",
          4197 => x"55",
          4198 => x"09",
          4199 => x"38",
          4200 => x"ff",
          4201 => x"06",
          4202 => x"55",
          4203 => x"0a",
          4204 => x"aa",
          4205 => x"77",
          4206 => x"c7",
          4207 => x"c8",
          4208 => x"d3",
          4209 => x"96",
          4210 => x"a0",
          4211 => x"51",
          4212 => x"3f",
          4213 => x"0b",
          4214 => x"77",
          4215 => x"bf",
          4216 => x"52",
          4217 => x"51",
          4218 => x"3f",
          4219 => x"18",
          4220 => x"c3",
          4221 => x"53",
          4222 => x"80",
          4223 => x"ff",
          4224 => x"77",
          4225 => x"80",
          4226 => x"7e",
          4227 => x"18",
          4228 => x"c3",
          4229 => x"54",
          4230 => x"15",
          4231 => x"d4",
          4232 => x"e7",
          4233 => x"c8",
          4234 => x"d3",
          4235 => x"38",
          4236 => x"96",
          4237 => x"ae",
          4238 => x"53",
          4239 => x"51",
          4240 => x"63",
          4241 => x"8b",
          4242 => x"54",
          4243 => x"15",
          4244 => x"ff",
          4245 => x"91",
          4246 => x"55",
          4247 => x"53",
          4248 => x"3d",
          4249 => x"ff",
          4250 => x"74",
          4251 => x"0c",
          4252 => x"04",
          4253 => x"a8",
          4254 => x"51",
          4255 => x"82",
          4256 => x"ff",
          4257 => x"a8",
          4258 => x"d1",
          4259 => x"c8",
          4260 => x"d3",
          4261 => x"d7",
          4262 => x"a8",
          4263 => x"a7",
          4264 => x"51",
          4265 => x"91",
          4266 => x"55",
          4267 => x"08",
          4268 => x"02",
          4269 => x"33",
          4270 => x"54",
          4271 => x"83",
          4272 => x"74",
          4273 => x"a0",
          4274 => x"08",
          4275 => x"ff",
          4276 => x"ff",
          4277 => x"ac",
          4278 => x"d4",
          4279 => x"3d",
          4280 => x"ff",
          4281 => x"a9",
          4282 => x"73",
          4283 => x"3f",
          4284 => x"08",
          4285 => x"c8",
          4286 => x"62",
          4287 => x"81",
          4288 => x"84",
          4289 => x"3d",
          4290 => x"38",
          4291 => x"84",
          4292 => x"06",
          4293 => x"a7",
          4294 => x"05",
          4295 => x"3f",
          4296 => x"08",
          4297 => x"c8",
          4298 => x"38",
          4299 => x"53",
          4300 => x"95",
          4301 => x"16",
          4302 => x"ed",
          4303 => x"05",
          4304 => x"34",
          4305 => x"70",
          4306 => x"81",
          4307 => x"57",
          4308 => x"76",
          4309 => x"73",
          4310 => x"77",
          4311 => x"83",
          4312 => x"16",
          4313 => x"2a",
          4314 => x"51",
          4315 => x"80",
          4316 => x"38",
          4317 => x"80",
          4318 => x"52",
          4319 => x"bf",
          4320 => x"d3",
          4321 => x"77",
          4322 => x"b2",
          4323 => x"91",
          4324 => x"80",
          4325 => x"91",
          4326 => x"52",
          4327 => x"ae",
          4328 => x"d3",
          4329 => x"d4",
          4330 => x"91",
          4331 => x"bf",
          4332 => x"33",
          4333 => x"2e",
          4334 => x"92",
          4335 => x"75",
          4336 => x"ff",
          4337 => x"77",
          4338 => x"83",
          4339 => x"9f",
          4340 => x"d4",
          4341 => x"89",
          4342 => x"c8",
          4343 => x"d3",
          4344 => x"38",
          4345 => x"ae",
          4346 => x"d3",
          4347 => x"74",
          4348 => x"0c",
          4349 => x"04",
          4350 => x"02",
          4351 => x"33",
          4352 => x"80",
          4353 => x"57",
          4354 => x"95",
          4355 => x"52",
          4356 => x"cd",
          4357 => x"d3",
          4358 => x"91",
          4359 => x"80",
          4360 => x"5a",
          4361 => x"3d",
          4362 => x"c7",
          4363 => x"d3",
          4364 => x"91",
          4365 => x"bd",
          4366 => x"cf",
          4367 => x"a0",
          4368 => x"80",
          4369 => x"86",
          4370 => x"38",
          4371 => x"61",
          4372 => x"12",
          4373 => x"7a",
          4374 => x"51",
          4375 => x"74",
          4376 => x"78",
          4377 => x"83",
          4378 => x"51",
          4379 => x"3f",
          4380 => x"08",
          4381 => x"d3",
          4382 => x"3d",
          4383 => x"3d",
          4384 => x"82",
          4385 => x"d0",
          4386 => x"3d",
          4387 => x"3f",
          4388 => x"08",
          4389 => x"c8",
          4390 => x"38",
          4391 => x"52",
          4392 => x"05",
          4393 => x"3f",
          4394 => x"08",
          4395 => x"c8",
          4396 => x"02",
          4397 => x"33",
          4398 => x"54",
          4399 => x"83",
          4400 => x"74",
          4401 => x"16",
          4402 => x"22",
          4403 => x"72",
          4404 => x"54",
          4405 => x"51",
          4406 => x"3f",
          4407 => x"0b",
          4408 => x"77",
          4409 => x"a7",
          4410 => x"c8",
          4411 => x"91",
          4412 => x"94",
          4413 => x"ea",
          4414 => x"6b",
          4415 => x"53",
          4416 => x"05",
          4417 => x"51",
          4418 => x"91",
          4419 => x"91",
          4420 => x"30",
          4421 => x"c8",
          4422 => x"25",
          4423 => x"7d",
          4424 => x"72",
          4425 => x"51",
          4426 => x"80",
          4427 => x"38",
          4428 => x"5f",
          4429 => x"3d",
          4430 => x"ff",
          4431 => x"91",
          4432 => x"56",
          4433 => x"08",
          4434 => x"81",
          4435 => x"ff",
          4436 => x"91",
          4437 => x"56",
          4438 => x"08",
          4439 => x"d3",
          4440 => x"d3",
          4441 => x"5c",
          4442 => x"17",
          4443 => x"1a",
          4444 => x"74",
          4445 => x"81",
          4446 => x"77",
          4447 => x"77",
          4448 => x"74",
          4449 => x"2e",
          4450 => x"18",
          4451 => x"33",
          4452 => x"73",
          4453 => x"38",
          4454 => x"09",
          4455 => x"38",
          4456 => x"80",
          4457 => x"70",
          4458 => x"25",
          4459 => x"7e",
          4460 => x"72",
          4461 => x"51",
          4462 => x"2e",
          4463 => x"a0",
          4464 => x"51",
          4465 => x"3f",
          4466 => x"08",
          4467 => x"c8",
          4468 => x"7b",
          4469 => x"54",
          4470 => x"73",
          4471 => x"38",
          4472 => x"73",
          4473 => x"38",
          4474 => x"18",
          4475 => x"ff",
          4476 => x"91",
          4477 => x"7b",
          4478 => x"d3",
          4479 => x"3d",
          4480 => x"3d",
          4481 => x"9a",
          4482 => x"05",
          4483 => x"51",
          4484 => x"91",
          4485 => x"55",
          4486 => x"08",
          4487 => x"8b",
          4488 => x"9a",
          4489 => x"05",
          4490 => x"a1",
          4491 => x"70",
          4492 => x"57",
          4493 => x"74",
          4494 => x"38",
          4495 => x"81",
          4496 => x"81",
          4497 => x"56",
          4498 => x"3f",
          4499 => x"08",
          4500 => x"38",
          4501 => x"70",
          4502 => x"ff",
          4503 => x"91",
          4504 => x"80",
          4505 => x"75",
          4506 => x"07",
          4507 => x"4c",
          4508 => x"80",
          4509 => x"16",
          4510 => x"26",
          4511 => x"16",
          4512 => x"ff",
          4513 => x"80",
          4514 => x"87",
          4515 => x"f8",
          4516 => x"75",
          4517 => x"38",
          4518 => x"bc",
          4519 => x"a6",
          4520 => x"d3",
          4521 => x"38",
          4522 => x"27",
          4523 => x"89",
          4524 => x"8b",
          4525 => x"27",
          4526 => x"55",
          4527 => x"81",
          4528 => x"93",
          4529 => x"77",
          4530 => x"05",
          4531 => x"55",
          4532 => x"34",
          4533 => x"9a",
          4534 => x"ff",
          4535 => x"75",
          4536 => x"17",
          4537 => x"56",
          4538 => x"9f",
          4539 => x"38",
          4540 => x"54",
          4541 => x"81",
          4542 => x"ea",
          4543 => x"2e",
          4544 => x"9f",
          4545 => x"12",
          4546 => x"52",
          4547 => x"a0",
          4548 => x"06",
          4549 => x"17",
          4550 => x"2e",
          4551 => x"15",
          4552 => x"54",
          4553 => x"ee",
          4554 => x"80",
          4555 => x"8f",
          4556 => x"55",
          4557 => x"3f",
          4558 => x"08",
          4559 => x"c8",
          4560 => x"38",
          4561 => x"51",
          4562 => x"3f",
          4563 => x"08",
          4564 => x"c8",
          4565 => x"76",
          4566 => x"38",
          4567 => x"3d",
          4568 => x"52",
          4569 => x"a4",
          4570 => x"39",
          4571 => x"74",
          4572 => x"81",
          4573 => x"34",
          4574 => x"a7",
          4575 => x"d3",
          4576 => x"80",
          4577 => x"d3",
          4578 => x"2e",
          4579 => x"80",
          4580 => x"54",
          4581 => x"80",
          4582 => x"52",
          4583 => x"05",
          4584 => x"b2",
          4585 => x"c8",
          4586 => x"d3",
          4587 => x"38",
          4588 => x"d3",
          4589 => x"65",
          4590 => x"91",
          4591 => x"88",
          4592 => x"34",
          4593 => x"3d",
          4594 => x"52",
          4595 => x"a3",
          4596 => x"54",
          4597 => x"15",
          4598 => x"ff",
          4599 => x"91",
          4600 => x"54",
          4601 => x"91",
          4602 => x"9a",
          4603 => x"f1",
          4604 => x"63",
          4605 => x"80",
          4606 => x"94",
          4607 => x"55",
          4608 => x"5c",
          4609 => x"3f",
          4610 => x"08",
          4611 => x"c8",
          4612 => x"91",
          4613 => x"76",
          4614 => x"38",
          4615 => x"b7",
          4616 => x"2e",
          4617 => x"18",
          4618 => x"90",
          4619 => x"81",
          4620 => x"06",
          4621 => x"73",
          4622 => x"54",
          4623 => x"82",
          4624 => x"39",
          4625 => x"84",
          4626 => x"11",
          4627 => x"2b",
          4628 => x"54",
          4629 => x"fe",
          4630 => x"ff",
          4631 => x"70",
          4632 => x"07",
          4633 => x"d3",
          4634 => x"62",
          4635 => x"5d",
          4636 => x"55",
          4637 => x"79",
          4638 => x"98",
          4639 => x"26",
          4640 => x"59",
          4641 => x"5d",
          4642 => x"52",
          4643 => x"a6",
          4644 => x"d3",
          4645 => x"16",
          4646 => x"56",
          4647 => x"75",
          4648 => x"82",
          4649 => x"2e",
          4650 => x"75",
          4651 => x"94",
          4652 => x"38",
          4653 => x"79",
          4654 => x"38",
          4655 => x"5d",
          4656 => x"79",
          4657 => x"06",
          4658 => x"57",
          4659 => x"38",
          4660 => x"b9",
          4661 => x"57",
          4662 => x"2e",
          4663 => x"15",
          4664 => x"2e",
          4665 => x"83",
          4666 => x"73",
          4667 => x"7f",
          4668 => x"f0",
          4669 => x"c8",
          4670 => x"d3",
          4671 => x"38",
          4672 => x"ff",
          4673 => x"5f",
          4674 => x"84",
          4675 => x"5f",
          4676 => x"38",
          4677 => x"12",
          4678 => x"80",
          4679 => x"7c",
          4680 => x"7a",
          4681 => x"90",
          4682 => x"c0",
          4683 => x"90",
          4684 => x"98",
          4685 => x"05",
          4686 => x"15",
          4687 => x"95",
          4688 => x"08",
          4689 => x"16",
          4690 => x"11",
          4691 => x"55",
          4692 => x"16",
          4693 => x"73",
          4694 => x"0c",
          4695 => x"04",
          4696 => x"6a",
          4697 => x"80",
          4698 => x"9b",
          4699 => x"58",
          4700 => x"3f",
          4701 => x"08",
          4702 => x"80",
          4703 => x"c8",
          4704 => x"d1",
          4705 => x"c8",
          4706 => x"91",
          4707 => x"55",
          4708 => x"2e",
          4709 => x"08",
          4710 => x"34",
          4711 => x"06",
          4712 => x"79",
          4713 => x"cb",
          4714 => x"c8",
          4715 => x"06",
          4716 => x"56",
          4717 => x"74",
          4718 => x"75",
          4719 => x"81",
          4720 => x"8a",
          4721 => x"8d",
          4722 => x"fc",
          4723 => x"52",
          4724 => x"9d",
          4725 => x"d3",
          4726 => x"38",
          4727 => x"93",
          4728 => x"80",
          4729 => x"38",
          4730 => x"67",
          4731 => x"80",
          4732 => x"81",
          4733 => x"5e",
          4734 => x"86",
          4735 => x"26",
          4736 => x"81",
          4737 => x"8b",
          4738 => x"78",
          4739 => x"80",
          4740 => x"93",
          4741 => x"39",
          4742 => x"51",
          4743 => x"3f",
          4744 => x"08",
          4745 => x"6e",
          4746 => x"fe",
          4747 => x"91",
          4748 => x"7e",
          4749 => x"08",
          4750 => x"70",
          4751 => x"25",
          4752 => x"08",
          4753 => x"d3",
          4754 => x"80",
          4755 => x"52",
          4756 => x"46",
          4757 => x"75",
          4758 => x"98",
          4759 => x"53",
          4760 => x"51",
          4761 => x"3f",
          4762 => x"d3",
          4763 => x"e5",
          4764 => x"2a",
          4765 => x"51",
          4766 => x"74",
          4767 => x"81",
          4768 => x"bf",
          4769 => x"63",
          4770 => x"c9",
          4771 => x"31",
          4772 => x"80",
          4773 => x"8a",
          4774 => x"57",
          4775 => x"26",
          4776 => x"7c",
          4777 => x"81",
          4778 => x"74",
          4779 => x"38",
          4780 => x"55",
          4781 => x"88",
          4782 => x"06",
          4783 => x"38",
          4784 => x"39",
          4785 => x"55",
          4786 => x"42",
          4787 => x"8a",
          4788 => x"59",
          4789 => x"09",
          4790 => x"f1",
          4791 => x"38",
          4792 => x"78",
          4793 => x"0b",
          4794 => x"70",
          4795 => x"58",
          4796 => x"80",
          4797 => x"74",
          4798 => x"38",
          4799 => x"10",
          4800 => x"70",
          4801 => x"5a",
          4802 => x"2e",
          4803 => x"75",
          4804 => x"78",
          4805 => x"fe",
          4806 => x"91",
          4807 => x"91",
          4808 => x"10",
          4809 => x"54",
          4810 => x"56",
          4811 => x"3f",
          4812 => x"08",
          4813 => x"80",
          4814 => x"8a",
          4815 => x"fd",
          4816 => x"75",
          4817 => x"38",
          4818 => x"89",
          4819 => x"38",
          4820 => x"78",
          4821 => x"0b",
          4822 => x"70",
          4823 => x"58",
          4824 => x"80",
          4825 => x"74",
          4826 => x"38",
          4827 => x"10",
          4828 => x"70",
          4829 => x"5a",
          4830 => x"2e",
          4831 => x"75",
          4832 => x"78",
          4833 => x"fe",
          4834 => x"91",
          4835 => x"10",
          4836 => x"91",
          4837 => x"9f",
          4838 => x"38",
          4839 => x"d3",
          4840 => x"29",
          4841 => x"2a",
          4842 => x"58",
          4843 => x"76",
          4844 => x"51",
          4845 => x"3f",
          4846 => x"08",
          4847 => x"53",
          4848 => x"80",
          4849 => x"ef",
          4850 => x"c8",
          4851 => x"ff",
          4852 => x"1b",
          4853 => x"05",
          4854 => x"05",
          4855 => x"72",
          4856 => x"52",
          4857 => x"40",
          4858 => x"09",
          4859 => x"38",
          4860 => x"18",
          4861 => x"39",
          4862 => x"78",
          4863 => x"70",
          4864 => x"55",
          4865 => x"87",
          4866 => x"7b",
          4867 => x"79",
          4868 => x"31",
          4869 => x"f2",
          4870 => x"d3",
          4871 => x"61",
          4872 => x"81",
          4873 => x"91",
          4874 => x"83",
          4875 => x"91",
          4876 => x"38",
          4877 => x"58",
          4878 => x"38",
          4879 => x"95",
          4880 => x"2e",
          4881 => x"80",
          4882 => x"ff",
          4883 => x"b4",
          4884 => x"38",
          4885 => x"74",
          4886 => x"86",
          4887 => x"fc",
          4888 => x"81",
          4889 => x"55",
          4890 => x"86",
          4891 => x"fc",
          4892 => x"8b",
          4893 => x"58",
          4894 => x"27",
          4895 => x"8e",
          4896 => x"39",
          4897 => x"26",
          4898 => x"8b",
          4899 => x"58",
          4900 => x"27",
          4901 => x"8e",
          4902 => x"39",
          4903 => x"81",
          4904 => x"06",
          4905 => x"55",
          4906 => x"26",
          4907 => x"8e",
          4908 => x"a1",
          4909 => x"80",
          4910 => x"ff",
          4911 => x"8b",
          4912 => x"b4",
          4913 => x"ff",
          4914 => x"7d",
          4915 => x"51",
          4916 => x"3f",
          4917 => x"05",
          4918 => x"ff",
          4919 => x"8e",
          4920 => x"98",
          4921 => x"7f",
          4922 => x"61",
          4923 => x"30",
          4924 => x"84",
          4925 => x"51",
          4926 => x"51",
          4927 => x"3f",
          4928 => x"ff",
          4929 => x"02",
          4930 => x"22",
          4931 => x"51",
          4932 => x"3f",
          4933 => x"52",
          4934 => x"ff",
          4935 => x"f8",
          4936 => x"34",
          4937 => x"1f",
          4938 => x"b0",
          4939 => x"52",
          4940 => x"ff",
          4941 => x"63",
          4942 => x"51",
          4943 => x"3f",
          4944 => x"09",
          4945 => x"cf",
          4946 => x"b2",
          4947 => x"c3",
          4948 => x"98",
          4949 => x"52",
          4950 => x"ff",
          4951 => x"82",
          4952 => x"51",
          4953 => x"3f",
          4954 => x"1f",
          4955 => x"ec",
          4956 => x"b2",
          4957 => x"97",
          4958 => x"80",
          4959 => x"05",
          4960 => x"80",
          4961 => x"93",
          4962 => x"c0",
          4963 => x"1f",
          4964 => x"95",
          4965 => x"82",
          4966 => x"52",
          4967 => x"ff",
          4968 => x"7b",
          4969 => x"06",
          4970 => x"51",
          4971 => x"3f",
          4972 => x"a4",
          4973 => x"7f",
          4974 => x"93",
          4975 => x"d4",
          4976 => x"51",
          4977 => x"3f",
          4978 => x"52",
          4979 => x"51",
          4980 => x"3f",
          4981 => x"53",
          4982 => x"51",
          4983 => x"3f",
          4984 => x"d3",
          4985 => x"ed",
          4986 => x"2e",
          4987 => x"80",
          4988 => x"54",
          4989 => x"53",
          4990 => x"51",
          4991 => x"3f",
          4992 => x"52",
          4993 => x"97",
          4994 => x"8b",
          4995 => x"52",
          4996 => x"96",
          4997 => x"8a",
          4998 => x"52",
          4999 => x"51",
          5000 => x"3f",
          5001 => x"83",
          5002 => x"ff",
          5003 => x"82",
          5004 => x"1f",
          5005 => x"c2",
          5006 => x"d5",
          5007 => x"1f",
          5008 => x"98",
          5009 => x"63",
          5010 => x"7e",
          5011 => x"ff",
          5012 => x"81",
          5013 => x"05",
          5014 => x"79",
          5015 => x"f8",
          5016 => x"80",
          5017 => x"ff",
          5018 => x"7f",
          5019 => x"61",
          5020 => x"81",
          5021 => x"f8",
          5022 => x"ff",
          5023 => x"ff",
          5024 => x"51",
          5025 => x"3f",
          5026 => x"88",
          5027 => x"95",
          5028 => x"39",
          5029 => x"f8",
          5030 => x"2e",
          5031 => x"55",
          5032 => x"51",
          5033 => x"3f",
          5034 => x"57",
          5035 => x"83",
          5036 => x"76",
          5037 => x"7e",
          5038 => x"ff",
          5039 => x"91",
          5040 => x"82",
          5041 => x"53",
          5042 => x"51",
          5043 => x"3f",
          5044 => x"78",
          5045 => x"74",
          5046 => x"1b",
          5047 => x"2e",
          5048 => x"78",
          5049 => x"2e",
          5050 => x"55",
          5051 => x"61",
          5052 => x"74",
          5053 => x"75",
          5054 => x"79",
          5055 => x"d8",
          5056 => x"c8",
          5057 => x"38",
          5058 => x"78",
          5059 => x"74",
          5060 => x"57",
          5061 => x"93",
          5062 => x"65",
          5063 => x"26",
          5064 => x"57",
          5065 => x"83",
          5066 => x"7c",
          5067 => x"06",
          5068 => x"ff",
          5069 => x"77",
          5070 => x"ff",
          5071 => x"82",
          5072 => x"83",
          5073 => x"ff",
          5074 => x"83",
          5075 => x"77",
          5076 => x"0b",
          5077 => x"81",
          5078 => x"34",
          5079 => x"34",
          5080 => x"34",
          5081 => x"57",
          5082 => x"52",
          5083 => x"eb",
          5084 => x"0b",
          5085 => x"91",
          5086 => x"82",
          5087 => x"55",
          5088 => x"34",
          5089 => x"08",
          5090 => x"63",
          5091 => x"1f",
          5092 => x"e6",
          5093 => x"83",
          5094 => x"ff",
          5095 => x"81",
          5096 => x"7e",
          5097 => x"ff",
          5098 => x"81",
          5099 => x"c8",
          5100 => x"80",
          5101 => x"79",
          5102 => x"f6",
          5103 => x"91",
          5104 => x"91",
          5105 => x"8e",
          5106 => x"81",
          5107 => x"81",
          5108 => x"80",
          5109 => x"d3",
          5110 => x"3d",
          5111 => x"3d",
          5112 => x"71",
          5113 => x"e2",
          5114 => x"10",
          5115 => x"05",
          5116 => x"04",
          5117 => x"51",
          5118 => x"3f",
          5119 => x"91",
          5120 => x"ff",
          5121 => x"81",
          5122 => x"c2",
          5123 => x"80",
          5124 => x"be",
          5125 => x"ac",
          5126 => x"88",
          5127 => x"39",
          5128 => x"51",
          5129 => x"3f",
          5130 => x"91",
          5131 => x"fe",
          5132 => x"81",
          5133 => x"c2",
          5134 => x"ff",
          5135 => x"92",
          5136 => x"f0",
          5137 => x"dc",
          5138 => x"39",
          5139 => x"51",
          5140 => x"3f",
          5141 => x"91",
          5142 => x"fe",
          5143 => x"80",
          5144 => x"c3",
          5145 => x"ff",
          5146 => x"e6",
          5147 => x"d4",
          5148 => x"b0",
          5149 => x"39",
          5150 => x"51",
          5151 => x"3f",
          5152 => x"91",
          5153 => x"fe",
          5154 => x"80",
          5155 => x"c4",
          5156 => x"ff",
          5157 => x"39",
          5158 => x"51",
          5159 => x"3f",
          5160 => x"c4",
          5161 => x"fe",
          5162 => x"39",
          5163 => x"51",
          5164 => x"3f",
          5165 => x"c5",
          5166 => x"fe",
          5167 => x"39",
          5168 => x"51",
          5169 => x"3f",
          5170 => x"c5",
          5171 => x"fe",
          5172 => x"3d",
          5173 => x"3d",
          5174 => x"56",
          5175 => x"e7",
          5176 => x"74",
          5177 => x"e8",
          5178 => x"e8",
          5179 => x"d3",
          5180 => x"9a",
          5181 => x"52",
          5182 => x"e8",
          5183 => x"d3",
          5184 => x"75",
          5185 => x"af",
          5186 => x"c8",
          5187 => x"54",
          5188 => x"52",
          5189 => x"51",
          5190 => x"3f",
          5191 => x"04",
          5192 => x"0d",
          5193 => x"08",
          5194 => x"08",
          5195 => x"84",
          5196 => x"71",
          5197 => x"75",
          5198 => x"87",
          5199 => x"07",
          5200 => x"5c",
          5201 => x"55",
          5202 => x"38",
          5203 => x"52",
          5204 => x"fb",
          5205 => x"ff",
          5206 => x"91",
          5207 => x"58",
          5208 => x"08",
          5209 => x"d3",
          5210 => x"c0",
          5211 => x"91",
          5212 => x"59",
          5213 => x"fb",
          5214 => x"55",
          5215 => x"76",
          5216 => x"15",
          5217 => x"3f",
          5218 => x"08",
          5219 => x"c8",
          5220 => x"7a",
          5221 => x"38",
          5222 => x"18",
          5223 => x"39",
          5224 => x"fb",
          5225 => x"ca",
          5226 => x"30",
          5227 => x"80",
          5228 => x"70",
          5229 => x"06",
          5230 => x"56",
          5231 => x"90",
          5232 => x"e4",
          5233 => x"98",
          5234 => x"78",
          5235 => x"3f",
          5236 => x"91",
          5237 => x"81",
          5238 => x"04",
          5239 => x"02",
          5240 => x"57",
          5241 => x"59",
          5242 => x"52",
          5243 => x"b0",
          5244 => x"c8",
          5245 => x"76",
          5246 => x"38",
          5247 => x"98",
          5248 => x"61",
          5249 => x"91",
          5250 => x"7f",
          5251 => x"75",
          5252 => x"c8",
          5253 => x"39",
          5254 => x"91",
          5255 => x"8a",
          5256 => x"fb",
          5257 => x"9f",
          5258 => x"c5",
          5259 => x"c5",
          5260 => x"ff",
          5261 => x"91",
          5262 => x"22",
          5263 => x"f9",
          5264 => x"c6",
          5265 => x"c6",
          5266 => x"15",
          5267 => x"c6",
          5268 => x"81",
          5269 => x"80",
          5270 => x"fe",
          5271 => x"87",
          5272 => x"fe",
          5273 => x"c0",
          5274 => x"53",
          5275 => x"3f",
          5276 => x"ee",
          5277 => x"c6",
          5278 => x"f0",
          5279 => x"51",
          5280 => x"3f",
          5281 => x"70",
          5282 => x"52",
          5283 => x"95",
          5284 => x"fe",
          5285 => x"91",
          5286 => x"fe",
          5287 => x"80",
          5288 => x"d0",
          5289 => x"2a",
          5290 => x"51",
          5291 => x"2e",
          5292 => x"51",
          5293 => x"3f",
          5294 => x"51",
          5295 => x"3f",
          5296 => x"ee",
          5297 => x"83",
          5298 => x"06",
          5299 => x"80",
          5300 => x"81",
          5301 => x"9c",
          5302 => x"f0",
          5303 => x"92",
          5304 => x"fe",
          5305 => x"72",
          5306 => x"81",
          5307 => x"71",
          5308 => x"38",
          5309 => x"ed",
          5310 => x"c7",
          5311 => x"ef",
          5312 => x"51",
          5313 => x"3f",
          5314 => x"70",
          5315 => x"52",
          5316 => x"95",
          5317 => x"fe",
          5318 => x"91",
          5319 => x"fe",
          5320 => x"80",
          5321 => x"cc",
          5322 => x"2a",
          5323 => x"51",
          5324 => x"2e",
          5325 => x"51",
          5326 => x"3f",
          5327 => x"51",
          5328 => x"3f",
          5329 => x"ed",
          5330 => x"87",
          5331 => x"06",
          5332 => x"80",
          5333 => x"81",
          5334 => x"98",
          5335 => x"c0",
          5336 => x"8e",
          5337 => x"fe",
          5338 => x"72",
          5339 => x"81",
          5340 => x"71",
          5341 => x"38",
          5342 => x"ec",
          5343 => x"c7",
          5344 => x"ee",
          5345 => x"51",
          5346 => x"3f",
          5347 => x"3f",
          5348 => x"04",
          5349 => x"78",
          5350 => x"55",
          5351 => x"80",
          5352 => x"38",
          5353 => x"77",
          5354 => x"33",
          5355 => x"39",
          5356 => x"80",
          5357 => x"54",
          5358 => x"83",
          5359 => x"72",
          5360 => x"2a",
          5361 => x"53",
          5362 => x"74",
          5363 => x"a0",
          5364 => x"06",
          5365 => x"75",
          5366 => x"57",
          5367 => x"75",
          5368 => x"cc",
          5369 => x"08",
          5370 => x"52",
          5371 => x"d0",
          5372 => x"c8",
          5373 => x"84",
          5374 => x"72",
          5375 => x"a6",
          5376 => x"70",
          5377 => x"57",
          5378 => x"27",
          5379 => x"53",
          5380 => x"c8",
          5381 => x"0d",
          5382 => x"0d",
          5383 => x"f6",
          5384 => x"0c",
          5385 => x"8c",
          5386 => x"7b",
          5387 => x"c3",
          5388 => x"c8",
          5389 => x"06",
          5390 => x"2e",
          5391 => x"9f",
          5392 => x"94",
          5393 => x"70",
          5394 => x"fd",
          5395 => x"53",
          5396 => x"b0",
          5397 => x"b5",
          5398 => x"d3",
          5399 => x"79",
          5400 => x"38",
          5401 => x"51",
          5402 => x"3f",
          5403 => x"70",
          5404 => x"c8",
          5405 => x"f7",
          5406 => x"3d",
          5407 => x"80",
          5408 => x"5a",
          5409 => x"51",
          5410 => x"3f",
          5411 => x"51",
          5412 => x"3f",
          5413 => x"f8",
          5414 => x"f8",
          5415 => x"c8",
          5416 => x"70",
          5417 => x"59",
          5418 => x"26",
          5419 => x"78",
          5420 => x"b2",
          5421 => x"78",
          5422 => x"3d",
          5423 => x"53",
          5424 => x"51",
          5425 => x"3f",
          5426 => x"08",
          5427 => x"c8",
          5428 => x"fc",
          5429 => x"9a",
          5430 => x"fe",
          5431 => x"fe",
          5432 => x"fe",
          5433 => x"91",
          5434 => x"80",
          5435 => x"81",
          5436 => x"38",
          5437 => x"bf",
          5438 => x"02",
          5439 => x"33",
          5440 => x"ef",
          5441 => x"c8",
          5442 => x"06",
          5443 => x"38",
          5444 => x"51",
          5445 => x"3f",
          5446 => x"d6",
          5447 => x"f4",
          5448 => x"80",
          5449 => x"39",
          5450 => x"f4",
          5451 => x"f8",
          5452 => x"fd",
          5453 => x"d3",
          5454 => x"2e",
          5455 => x"80",
          5456 => x"02",
          5457 => x"33",
          5458 => x"e6",
          5459 => x"c8",
          5460 => x"c9",
          5461 => x"fb",
          5462 => x"96",
          5463 => x"fe",
          5464 => x"fe",
          5465 => x"fe",
          5466 => x"91",
          5467 => x"80",
          5468 => x"60",
          5469 => x"fa",
          5470 => x"fe",
          5471 => x"fe",
          5472 => x"fe",
          5473 => x"91",
          5474 => x"86",
          5475 => x"c8",
          5476 => x"53",
          5477 => x"52",
          5478 => x"52",
          5479 => x"94",
          5480 => x"05",
          5481 => x"52",
          5482 => x"29",
          5483 => x"05",
          5484 => x"d0",
          5485 => x"c8",
          5486 => x"8c",
          5487 => x"c8",
          5488 => x"9a",
          5489 => x"39",
          5490 => x"51",
          5491 => x"3f",
          5492 => x"9e",
          5493 => x"fe",
          5494 => x"fe",
          5495 => x"91",
          5496 => x"b5",
          5497 => x"05",
          5498 => x"e4",
          5499 => x"53",
          5500 => x"08",
          5501 => x"f6",
          5502 => x"d3",
          5503 => x"2e",
          5504 => x"91",
          5505 => x"51",
          5506 => x"fc",
          5507 => x"3d",
          5508 => x"51",
          5509 => x"3f",
          5510 => x"08",
          5511 => x"f8",
          5512 => x"fe",
          5513 => x"91",
          5514 => x"b5",
          5515 => x"05",
          5516 => x"e4",
          5517 => x"d3",
          5518 => x"3d",
          5519 => x"52",
          5520 => x"a3",
          5521 => x"c4",
          5522 => x"fc",
          5523 => x"80",
          5524 => x"c8",
          5525 => x"06",
          5526 => x"79",
          5527 => x"f6",
          5528 => x"d3",
          5529 => x"2e",
          5530 => x"91",
          5531 => x"51",
          5532 => x"fb",
          5533 => x"c9",
          5534 => x"f3",
          5535 => x"51",
          5536 => x"3f",
          5537 => x"91",
          5538 => x"fe",
          5539 => x"a2",
          5540 => x"e2",
          5541 => x"39",
          5542 => x"0b",
          5543 => x"84",
          5544 => x"81",
          5545 => x"94",
          5546 => x"c9",
          5547 => x"f2",
          5548 => x"be",
          5549 => x"dc",
          5550 => x"e8",
          5551 => x"83",
          5552 => x"94",
          5553 => x"80",
          5554 => x"c0",
          5555 => x"fb",
          5556 => x"3d",
          5557 => x"53",
          5558 => x"51",
          5559 => x"3f",
          5560 => x"08",
          5561 => x"8a",
          5562 => x"91",
          5563 => x"fe",
          5564 => x"60",
          5565 => x"b4",
          5566 => x"11",
          5567 => x"05",
          5568 => x"a5",
          5569 => x"c8",
          5570 => x"fa",
          5571 => x"52",
          5572 => x"51",
          5573 => x"3f",
          5574 => x"2d",
          5575 => x"08",
          5576 => x"c8",
          5577 => x"fa",
          5578 => x"d3",
          5579 => x"91",
          5580 => x"fe",
          5581 => x"fa",
          5582 => x"ca",
          5583 => x"f1",
          5584 => x"d1",
          5585 => x"aa",
          5586 => x"e0",
          5587 => x"d4",
          5588 => x"ff",
          5589 => x"ed",
          5590 => x"96",
          5591 => x"33",
          5592 => x"80",
          5593 => x"38",
          5594 => x"59",
          5595 => x"80",
          5596 => x"3d",
          5597 => x"51",
          5598 => x"3f",
          5599 => x"56",
          5600 => x"08",
          5601 => x"f8",
          5602 => x"91",
          5603 => x"a0",
          5604 => x"59",
          5605 => x"3f",
          5606 => x"58",
          5607 => x"57",
          5608 => x"81",
          5609 => x"55",
          5610 => x"80",
          5611 => x"80",
          5612 => x"51",
          5613 => x"91",
          5614 => x"5e",
          5615 => x"7c",
          5616 => x"59",
          5617 => x"7d",
          5618 => x"81",
          5619 => x"38",
          5620 => x"51",
          5621 => x"3f",
          5622 => x"80",
          5623 => x"0b",
          5624 => x"34",
          5625 => x"e4",
          5626 => x"94",
          5627 => x"90",
          5628 => x"87",
          5629 => x"0c",
          5630 => x"0b",
          5631 => x"84",
          5632 => x"83",
          5633 => x"94",
          5634 => x"94",
          5635 => x"d3",
          5636 => x"97",
          5637 => x"d3",
          5638 => x"e8",
          5639 => x"ee",
          5640 => x"cb",
          5641 => x"e5",
          5642 => x"cb",
          5643 => x"ef",
          5644 => x"a4",
          5645 => x"ee",
          5646 => x"51",
          5647 => x"f7",
          5648 => x"04",
          5649 => x"0f",
          5650 => x"0f",
          5651 => x"0f",
          5652 => x"0f",
          5653 => x"0f",
          5654 => x"0f",
          5655 => x"11",
          5656 => x"11",
          5657 => x"11",
          5658 => x"11",
          5659 => x"11",
          5660 => x"11",
          5661 => x"11",
          5662 => x"11",
          5663 => x"11",
          5664 => x"11",
          5665 => x"11",
          5666 => x"11",
          5667 => x"11",
          5668 => x"11",
          5669 => x"11",
          5670 => x"11",
          5671 => x"11",
          5672 => x"11",
          5673 => x"11",
          5674 => x"11",
          5675 => x"11",
          5676 => x"11",
          5677 => x"11",
          5678 => x"50",
          5679 => x"4f",
          5680 => x"4f",
          5681 => x"50",
          5682 => x"50",
          5683 => x"50",
          5684 => x"50",
          5685 => x"50",
          5686 => x"50",
          5687 => x"50",
          5688 => x"50",
          5689 => x"50",
          5690 => x"50",
          5691 => x"50",
          5692 => x"50",
          5693 => x"50",
          5694 => x"50",
          5695 => x"50",
          5696 => x"50",
          5697 => x"50",
          5698 => x"54",
          5699 => x"57",
          5700 => x"54",
          5701 => x"57",
          5702 => x"55",
          5703 => x"57",
          5704 => x"57",
          5705 => x"57",
          5706 => x"57",
          5707 => x"57",
          5708 => x"57",
          5709 => x"57",
          5710 => x"57",
          5711 => x"57",
          5712 => x"57",
          5713 => x"57",
          5714 => x"57",
          5715 => x"57",
          5716 => x"57",
          5717 => x"57",
          5718 => x"55",
          5719 => x"57",
          5720 => x"57",
          5721 => x"57",
          5722 => x"57",
          5723 => x"57",
          5724 => x"57",
          5725 => x"57",
          5726 => x"57",
          5727 => x"57",
          5728 => x"57",
          5729 => x"57",
          5730 => x"57",
          5731 => x"57",
          5732 => x"57",
          5733 => x"57",
          5734 => x"57",
          5735 => x"57",
          5736 => x"57",
          5737 => x"57",
          5738 => x"57",
          5739 => x"57",
          5740 => x"57",
          5741 => x"55",
          5742 => x"57",
          5743 => x"57",
          5744 => x"57",
          5745 => x"57",
          5746 => x"56",
          5747 => x"57",
          5748 => x"57",
          5749 => x"57",
          5750 => x"57",
          5751 => x"57",
          5752 => x"57",
          5753 => x"57",
          5754 => x"57",
          5755 => x"57",
          5756 => x"57",
          5757 => x"57",
          5758 => x"57",
          5759 => x"57",
          5760 => x"57",
          5761 => x"57",
          5762 => x"57",
          5763 => x"57",
          5764 => x"57",
          5765 => x"57",
          5766 => x"57",
          5767 => x"57",
          5768 => x"57",
          5769 => x"57",
          5770 => x"57",
          5771 => x"57",
          5772 => x"57",
          5773 => x"57",
          5774 => x"57",
          5775 => x"57",
          5776 => x"57",
          5777 => x"57",
          5778 => x"56",
          5779 => x"56",
          5780 => x"57",
          5781 => x"57",
          5782 => x"56",
          5783 => x"56",
          5784 => x"57",
          5785 => x"57",
          5786 => x"57",
          5787 => x"57",
          5788 => x"57",
          5789 => x"57",
          5790 => x"57",
          5791 => x"57",
          5792 => x"57",
          5793 => x"57",
          5794 => x"57",
          5795 => x"57",
          5796 => x"57",
          5797 => x"57",
          5798 => x"57",
          5799 => x"57",
          5800 => x"57",
          5801 => x"57",
          5802 => x"57",
          5803 => x"57",
          5804 => x"57",
          5805 => x"57",
          5806 => x"57",
          5807 => x"57",
          5808 => x"57",
          5809 => x"57",
          5810 => x"57",
          5811 => x"57",
          5812 => x"57",
          5813 => x"57",
          5814 => x"57",
          5815 => x"57",
          5816 => x"57",
          5817 => x"57",
          5818 => x"56",
          5819 => x"56",
          5820 => x"57",
          5821 => x"57",
          5822 => x"57",
          5823 => x"57",
          5824 => x"57",
          5825 => x"57",
          5826 => x"57",
          5827 => x"57",
          5828 => x"57",
          5829 => x"57",
          5830 => x"57",
          5831 => x"57",
          5832 => x"57",
          5833 => x"54",
          5834 => x"2f",
          5835 => x"25",
          5836 => x"64",
          5837 => x"3a",
          5838 => x"25",
          5839 => x"0a",
          5840 => x"43",
          5841 => x"6e",
          5842 => x"75",
          5843 => x"69",
          5844 => x"00",
          5845 => x"66",
          5846 => x"20",
          5847 => x"20",
          5848 => x"66",
          5849 => x"00",
          5850 => x"44",
          5851 => x"63",
          5852 => x"69",
          5853 => x"65",
          5854 => x"74",
          5855 => x"0a",
          5856 => x"20",
          5857 => x"53",
          5858 => x"52",
          5859 => x"28",
          5860 => x"72",
          5861 => x"30",
          5862 => x"20",
          5863 => x"65",
          5864 => x"38",
          5865 => x"0a",
          5866 => x"20",
          5867 => x"41",
          5868 => x"53",
          5869 => x"74",
          5870 => x"38",
          5871 => x"53",
          5872 => x"3d",
          5873 => x"58",
          5874 => x"00",
          5875 => x"20",
          5876 => x"4d",
          5877 => x"74",
          5878 => x"3d",
          5879 => x"58",
          5880 => x"69",
          5881 => x"25",
          5882 => x"29",
          5883 => x"00",
          5884 => x"20",
          5885 => x"43",
          5886 => x"00",
          5887 => x"20",
          5888 => x"32",
          5889 => x"00",
          5890 => x"20",
          5891 => x"49",
          5892 => x"00",
          5893 => x"20",
          5894 => x"20",
          5895 => x"64",
          5896 => x"65",
          5897 => x"65",
          5898 => x"30",
          5899 => x"2e",
          5900 => x"00",
          5901 => x"20",
          5902 => x"54",
          5903 => x"55",
          5904 => x"43",
          5905 => x"52",
          5906 => x"45",
          5907 => x"00",
          5908 => x"20",
          5909 => x"4d",
          5910 => x"20",
          5911 => x"6d",
          5912 => x"3d",
          5913 => x"58",
          5914 => x"00",
          5915 => x"64",
          5916 => x"73",
          5917 => x"0a",
          5918 => x"20",
          5919 => x"55",
          5920 => x"73",
          5921 => x"56",
          5922 => x"6f",
          5923 => x"64",
          5924 => x"73",
          5925 => x"20",
          5926 => x"58",
          5927 => x"00",
          5928 => x"20",
          5929 => x"55",
          5930 => x"6d",
          5931 => x"20",
          5932 => x"72",
          5933 => x"64",
          5934 => x"73",
          5935 => x"20",
          5936 => x"58",
          5937 => x"00",
          5938 => x"20",
          5939 => x"61",
          5940 => x"53",
          5941 => x"74",
          5942 => x"64",
          5943 => x"73",
          5944 => x"20",
          5945 => x"20",
          5946 => x"58",
          5947 => x"00",
          5948 => x"20",
          5949 => x"55",
          5950 => x"20",
          5951 => x"20",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"20",
          5956 => x"58",
          5957 => x"00",
          5958 => x"20",
          5959 => x"73",
          5960 => x"20",
          5961 => x"63",
          5962 => x"72",
          5963 => x"20",
          5964 => x"20",
          5965 => x"20",
          5966 => x"58",
          5967 => x"00",
          5968 => x"61",
          5969 => x"00",
          5970 => x"64",
          5971 => x"00",
          5972 => x"65",
          5973 => x"00",
          5974 => x"4f",
          5975 => x"4f",
          5976 => x"00",
          5977 => x"6b",
          5978 => x"6e",
          5979 => x"00",
          5980 => x"2b",
          5981 => x"3c",
          5982 => x"5b",
          5983 => x"00",
          5984 => x"54",
          5985 => x"54",
          5986 => x"00",
          5987 => x"00",
          5988 => x"00",
          5989 => x"00",
          5990 => x"00",
          5991 => x"00",
          5992 => x"00",
          5993 => x"00",
          5994 => x"00",
          5995 => x"00",
          5996 => x"0a",
          5997 => x"90",
          5998 => x"4f",
          5999 => x"30",
          6000 => x"20",
          6001 => x"45",
          6002 => x"20",
          6003 => x"33",
          6004 => x"20",
          6005 => x"20",
          6006 => x"45",
          6007 => x"20",
          6008 => x"20",
          6009 => x"20",
          6010 => x"5d",
          6011 => x"00",
          6012 => x"00",
          6013 => x"00",
          6014 => x"45",
          6015 => x"8f",
          6016 => x"45",
          6017 => x"8e",
          6018 => x"92",
          6019 => x"55",
          6020 => x"9a",
          6021 => x"9e",
          6022 => x"4f",
          6023 => x"a6",
          6024 => x"aa",
          6025 => x"ae",
          6026 => x"b2",
          6027 => x"b6",
          6028 => x"ba",
          6029 => x"be",
          6030 => x"c2",
          6031 => x"c6",
          6032 => x"ca",
          6033 => x"ce",
          6034 => x"d2",
          6035 => x"d6",
          6036 => x"da",
          6037 => x"de",
          6038 => x"e2",
          6039 => x"e6",
          6040 => x"ea",
          6041 => x"ee",
          6042 => x"f2",
          6043 => x"f6",
          6044 => x"fa",
          6045 => x"fe",
          6046 => x"2c",
          6047 => x"5d",
          6048 => x"2a",
          6049 => x"3f",
          6050 => x"00",
          6051 => x"00",
          6052 => x"00",
          6053 => x"02",
          6054 => x"00",
          6055 => x"00",
          6056 => x"00",
          6057 => x"00",
          6058 => x"00",
          6059 => x"54",
          6060 => x"00",
          6061 => x"54",
          6062 => x"00",
          6063 => x"46",
          6064 => x"00",
          6065 => x"53",
          6066 => x"4f",
          6067 => x"4e",
          6068 => x"4c",
          6069 => x"00",
          6070 => x"53",
          6071 => x"55",
          6072 => x"52",
          6073 => x"4e",
          6074 => x"4c",
          6075 => x"00",
          6076 => x"4c",
          6077 => x"53",
          6078 => x"20",
          6079 => x"54",
          6080 => x"53",
          6081 => x"4d",
          6082 => x"00",
          6083 => x"52",
          6084 => x"52",
          6085 => x"00",
          6086 => x"53",
          6087 => x"47",
          6088 => x"45",
          6089 => x"49",
          6090 => x"00",
          6091 => x"53",
          6092 => x"4f",
          6093 => x"4e",
          6094 => x"00",
          6095 => x"75",
          6096 => x"00",
          6097 => x"6e",
          6098 => x"00",
          6099 => x"74",
          6100 => x"00",
          6101 => x"6f",
          6102 => x"00",
          6103 => x"75",
          6104 => x"00",
          6105 => x"64",
          6106 => x"00",
          6107 => x"65",
          6108 => x"00",
          6109 => x"72",
          6110 => x"00",
          6111 => x"69",
          6112 => x"00",
          6113 => x"65",
          6114 => x"00",
          6115 => x"6e",
          6116 => x"00",
          6117 => x"70",
          6118 => x"00",
          6119 => x"6c",
          6120 => x"00",
          6121 => x"65",
          6122 => x"00",
          6123 => x"65",
          6124 => x"00",
          6125 => x"6e",
          6126 => x"63",
          6127 => x"00",
          6128 => x"72",
          6129 => x"00",
          6130 => x"72",
          6131 => x"00",
          6132 => x"6c",
          6133 => x"00",
          6134 => x"74",
          6135 => x"00",
          6136 => x"69",
          6137 => x"00",
          6138 => x"65",
          6139 => x"65",
          6140 => x"65",
          6141 => x"00",
          6142 => x"6b",
          6143 => x"00",
          6144 => x"74",
          6145 => x"00",
          6146 => x"69",
          6147 => x"00",
          6148 => x"61",
          6149 => x"00",
          6150 => x"70",
          6151 => x"6f",
          6152 => x"74",
          6153 => x"74",
          6154 => x"74",
          6155 => x"6f",
          6156 => x"00",
          6157 => x"78",
          6158 => x"00",
          6159 => x"61",
          6160 => x"00",
          6161 => x"75",
          6162 => x"00",
          6163 => x"64",
          6164 => x"72",
          6165 => x"00",
          6166 => x"68",
          6167 => x"69",
          6168 => x"00",
          6169 => x"61",
          6170 => x"00",
          6171 => x"6b",
          6172 => x"00",
          6173 => x"6c",
          6174 => x"00",
          6175 => x"75",
          6176 => x"00",
          6177 => x"62",
          6178 => x"68",
          6179 => x"77",
          6180 => x"64",
          6181 => x"65",
          6182 => x"00",
          6183 => x"00",
          6184 => x"64",
          6185 => x"65",
          6186 => x"72",
          6187 => x"00",
          6188 => x"72",
          6189 => x"72",
          6190 => x"00",
          6191 => x"6c",
          6192 => x"00",
          6193 => x"70",
          6194 => x"73",
          6195 => x"74",
          6196 => x"73",
          6197 => x"00",
          6198 => x"6c",
          6199 => x"00",
          6200 => x"66",
          6201 => x"00",
          6202 => x"6d",
          6203 => x"00",
          6204 => x"73",
          6205 => x"00",
          6206 => x"73",
          6207 => x"72",
          6208 => x"0a",
          6209 => x"74",
          6210 => x"61",
          6211 => x"72",
          6212 => x"2e",
          6213 => x"00",
          6214 => x"73",
          6215 => x"6f",
          6216 => x"65",
          6217 => x"2e",
          6218 => x"00",
          6219 => x"20",
          6220 => x"65",
          6221 => x"75",
          6222 => x"0a",
          6223 => x"20",
          6224 => x"68",
          6225 => x"75",
          6226 => x"0a",
          6227 => x"76",
          6228 => x"64",
          6229 => x"6c",
          6230 => x"6d",
          6231 => x"00",
          6232 => x"63",
          6233 => x"20",
          6234 => x"69",
          6235 => x"0a",
          6236 => x"6c",
          6237 => x"6c",
          6238 => x"64",
          6239 => x"78",
          6240 => x"73",
          6241 => x"00",
          6242 => x"6c",
          6243 => x"61",
          6244 => x"65",
          6245 => x"76",
          6246 => x"64",
          6247 => x"00",
          6248 => x"20",
          6249 => x"77",
          6250 => x"65",
          6251 => x"6f",
          6252 => x"74",
          6253 => x"0a",
          6254 => x"69",
          6255 => x"6e",
          6256 => x"65",
          6257 => x"73",
          6258 => x"76",
          6259 => x"64",
          6260 => x"00",
          6261 => x"73",
          6262 => x"6f",
          6263 => x"6e",
          6264 => x"65",
          6265 => x"00",
          6266 => x"20",
          6267 => x"70",
          6268 => x"62",
          6269 => x"66",
          6270 => x"73",
          6271 => x"65",
          6272 => x"6f",
          6273 => x"20",
          6274 => x"64",
          6275 => x"2e",
          6276 => x"00",
          6277 => x"72",
          6278 => x"20",
          6279 => x"72",
          6280 => x"2e",
          6281 => x"00",
          6282 => x"6d",
          6283 => x"74",
          6284 => x"70",
          6285 => x"74",
          6286 => x"20",
          6287 => x"63",
          6288 => x"65",
          6289 => x"00",
          6290 => x"6c",
          6291 => x"73",
          6292 => x"63",
          6293 => x"2e",
          6294 => x"00",
          6295 => x"73",
          6296 => x"69",
          6297 => x"6e",
          6298 => x"65",
          6299 => x"79",
          6300 => x"00",
          6301 => x"6f",
          6302 => x"6e",
          6303 => x"70",
          6304 => x"66",
          6305 => x"73",
          6306 => x"00",
          6307 => x"72",
          6308 => x"74",
          6309 => x"20",
          6310 => x"6f",
          6311 => x"63",
          6312 => x"00",
          6313 => x"63",
          6314 => x"73",
          6315 => x"00",
          6316 => x"6b",
          6317 => x"6e",
          6318 => x"72",
          6319 => x"0a",
          6320 => x"6c",
          6321 => x"79",
          6322 => x"20",
          6323 => x"61",
          6324 => x"6c",
          6325 => x"79",
          6326 => x"2f",
          6327 => x"2e",
          6328 => x"00",
          6329 => x"61",
          6330 => x"00",
          6331 => x"55",
          6332 => x"00",
          6333 => x"2a",
          6334 => x"20",
          6335 => x"00",
          6336 => x"2f",
          6337 => x"32",
          6338 => x"00",
          6339 => x"2e",
          6340 => x"00",
          6341 => x"50",
          6342 => x"72",
          6343 => x"25",
          6344 => x"29",
          6345 => x"20",
          6346 => x"2a",
          6347 => x"00",
          6348 => x"55",
          6349 => x"49",
          6350 => x"72",
          6351 => x"74",
          6352 => x"6e",
          6353 => x"72",
          6354 => x"00",
          6355 => x"6d",
          6356 => x"69",
          6357 => x"72",
          6358 => x"74",
          6359 => x"00",
          6360 => x"32",
          6361 => x"74",
          6362 => x"75",
          6363 => x"00",
          6364 => x"43",
          6365 => x"52",
          6366 => x"6e",
          6367 => x"72",
          6368 => x"0a",
          6369 => x"43",
          6370 => x"57",
          6371 => x"6e",
          6372 => x"72",
          6373 => x"0a",
          6374 => x"52",
          6375 => x"52",
          6376 => x"6e",
          6377 => x"72",
          6378 => x"0a",
          6379 => x"52",
          6380 => x"54",
          6381 => x"6e",
          6382 => x"72",
          6383 => x"0a",
          6384 => x"52",
          6385 => x"52",
          6386 => x"6e",
          6387 => x"72",
          6388 => x"0a",
          6389 => x"52",
          6390 => x"54",
          6391 => x"6e",
          6392 => x"72",
          6393 => x"0a",
          6394 => x"74",
          6395 => x"67",
          6396 => x"20",
          6397 => x"65",
          6398 => x"2e",
          6399 => x"00",
          6400 => x"61",
          6401 => x"6e",
          6402 => x"69",
          6403 => x"2e",
          6404 => x"00",
          6405 => x"00",
          6406 => x"69",
          6407 => x"20",
          6408 => x"69",
          6409 => x"69",
          6410 => x"73",
          6411 => x"64",
          6412 => x"72",
          6413 => x"2c",
          6414 => x"65",
          6415 => x"20",
          6416 => x"74",
          6417 => x"6e",
          6418 => x"6c",
          6419 => x"00",
          6420 => x"00",
          6421 => x"64",
          6422 => x"73",
          6423 => x"64",
          6424 => x"00",
          6425 => x"69",
          6426 => x"6c",
          6427 => x"64",
          6428 => x"00",
          6429 => x"69",
          6430 => x"20",
          6431 => x"69",
          6432 => x"69",
          6433 => x"73",
          6434 => x"00",
          6435 => x"3d",
          6436 => x"00",
          6437 => x"3a",
          6438 => x"73",
          6439 => x"69",
          6440 => x"69",
          6441 => x"72",
          6442 => x"74",
          6443 => x"00",
          6444 => x"61",
          6445 => x"6e",
          6446 => x"6e",
          6447 => x"72",
          6448 => x"73",
          6449 => x"00",
          6450 => x"73",
          6451 => x"65",
          6452 => x"61",
          6453 => x"66",
          6454 => x"0a",
          6455 => x"61",
          6456 => x"6e",
          6457 => x"61",
          6458 => x"66",
          6459 => x"0a",
          6460 => x"65",
          6461 => x"69",
          6462 => x"63",
          6463 => x"20",
          6464 => x"30",
          6465 => x"2e",
          6466 => x"00",
          6467 => x"6c",
          6468 => x"67",
          6469 => x"64",
          6470 => x"20",
          6471 => x"78",
          6472 => x"2e",
          6473 => x"00",
          6474 => x"6c",
          6475 => x"65",
          6476 => x"6e",
          6477 => x"63",
          6478 => x"20",
          6479 => x"29",
          6480 => x"00",
          6481 => x"73",
          6482 => x"74",
          6483 => x"20",
          6484 => x"6c",
          6485 => x"74",
          6486 => x"2e",
          6487 => x"00",
          6488 => x"6c",
          6489 => x"65",
          6490 => x"74",
          6491 => x"2e",
          6492 => x"00",
          6493 => x"55",
          6494 => x"6e",
          6495 => x"3a",
          6496 => x"5c",
          6497 => x"25",
          6498 => x"00",
          6499 => x"64",
          6500 => x"6d",
          6501 => x"64",
          6502 => x"00",
          6503 => x"6e",
          6504 => x"67",
          6505 => x"0a",
          6506 => x"61",
          6507 => x"6e",
          6508 => x"6e",
          6509 => x"72",
          6510 => x"73",
          6511 => x"0a",
          6512 => x"00",
          6513 => x"00",
          6514 => x"7f",
          6515 => x"00",
          6516 => x"7f",
          6517 => x"00",
          6518 => x"7f",
          6519 => x"00",
          6520 => x"00",
          6521 => x"78",
          6522 => x"00",
          6523 => x"e1",
          6524 => x"01",
          6525 => x"01",
          6526 => x"01",
          6527 => x"00",
          6528 => x"00",
          6529 => x"00",
          6530 => x"5f",
          6531 => x"01",
          6532 => x"00",
          6533 => x"00",
          6534 => x"5f",
          6535 => x"01",
          6536 => x"00",
          6537 => x"00",
          6538 => x"5f",
          6539 => x"01",
          6540 => x"00",
          6541 => x"00",
          6542 => x"5f",
          6543 => x"01",
          6544 => x"00",
          6545 => x"00",
          6546 => x"5f",
          6547 => x"02",
          6548 => x"00",
          6549 => x"00",
          6550 => x"5f",
          6551 => x"02",
          6552 => x"00",
          6553 => x"00",
          6554 => x"5f",
          6555 => x"02",
          6556 => x"00",
          6557 => x"00",
          6558 => x"5f",
          6559 => x"02",
          6560 => x"00",
          6561 => x"00",
          6562 => x"5f",
          6563 => x"02",
          6564 => x"00",
          6565 => x"00",
          6566 => x"5f",
          6567 => x"02",
          6568 => x"00",
          6569 => x"00",
          6570 => x"5f",
          6571 => x"03",
          6572 => x"00",
          6573 => x"00",
          6574 => x"5f",
          6575 => x"03",
          6576 => x"00",
          6577 => x"00",
          6578 => x"5f",
          6579 => x"03",
          6580 => x"00",
          6581 => x"00",
          6582 => x"5f",
          6583 => x"03",
          6584 => x"00",
          6585 => x"00",
          6586 => x"5f",
          6587 => x"03",
          6588 => x"00",
          6589 => x"00",
          6590 => x"5f",
          6591 => x"03",
          6592 => x"00",
          6593 => x"00",
          6594 => x"5f",
          6595 => x"03",
          6596 => x"00",
          6597 => x"00",
          6598 => x"5f",
          6599 => x"03",
          6600 => x"00",
          6601 => x"00",
          6602 => x"5f",
          6603 => x"03",
          6604 => x"00",
          6605 => x"00",
          6606 => x"5f",
          6607 => x"03",
          6608 => x"00",
          6609 => x"00",
          6610 => x"5f",
          6611 => x"03",
          6612 => x"00",
          6613 => x"00",
          6614 => x"5f",
          6615 => x"03",
          6616 => x"00",
          6617 => x"00",
          6618 => x"5f",
          6619 => x"03",
          6620 => x"00",
          6621 => x"00",
          6622 => x"5f",
          6623 => x"03",
          6624 => x"00",
          6625 => x"00",
          6626 => x"60",
          6627 => x"03",
          6628 => x"00",
          6629 => x"00",
          6630 => x"60",
          6631 => x"03",
          6632 => x"00",
          6633 => x"00",
          6634 => x"60",
          6635 => x"03",
          6636 => x"00",
          6637 => x"00",
          6638 => x"60",
          6639 => x"03",
          6640 => x"00",
          6641 => x"00",
          6642 => x"60",
          6643 => x"03",
          6644 => x"00",
          6645 => x"00",
          6646 => x"60",
          6647 => x"03",
          6648 => x"00",
          6649 => x"00",
          6650 => x"60",
          6651 => x"03",
          6652 => x"00",
          6653 => x"00",
          6654 => x"60",
          6655 => x"03",
          6656 => x"00",
          6657 => x"00",
          6658 => x"60",
          6659 => x"03",
          6660 => x"00",
          6661 => x"00",
          6662 => x"60",
          6663 => x"03",
          6664 => x"00",
          6665 => x"00",
          6666 => x"60",
          6667 => x"03",
          6668 => x"00",
          6669 => x"00",
          6670 => x"60",
          6671 => x"03",
          6672 => x"00",
          6673 => x"00",
          6674 => x"60",
          6675 => x"03",
          6676 => x"00",
          6677 => x"00",
          6678 => x"60",
          6679 => x"03",
          6680 => x"00",
          6681 => x"00",
          6682 => x"60",
          6683 => x"03",
          6684 => x"00",
          6685 => x"00",
          6686 => x"60",
          6687 => x"04",
          6688 => x"00",
          6689 => x"00",
          6690 => x"60",
          6691 => x"04",
          6692 => x"00",
          6693 => x"00",
          6694 => x"60",
          6695 => x"04",
          6696 => x"00",
          6697 => x"00",
          6698 => x"60",
          6699 => x"04",
          6700 => x"00",
          6701 => x"00",
          6702 => x"60",
          6703 => x"04",
          6704 => x"00",
          6705 => x"00",
          6706 => x"60",
          6707 => x"05",
          6708 => x"00",
          6709 => x"00",
          6710 => x"60",
          6711 => x"05",
          6712 => x"00",
          6713 => x"00",
          6714 => x"60",
          6715 => x"05",
          6716 => x"00",
          6717 => x"00",
          6718 => x"60",
          6719 => x"05",
          6720 => x"00",
          6721 => x"00",
          6722 => x"60",
          6723 => x"05",
          6724 => x"00",
          6725 => x"00",
          6726 => x"60",
          6727 => x"05",
          6728 => x"00",
          6729 => x"00",
          6730 => x"60",
          6731 => x"06",
          6732 => x"00",
          6733 => x"00",
          6734 => x"60",
          6735 => x"06",
          6736 => x"00",
          6737 => x"00",
          6738 => x"60",
          6739 => x"07",
          6740 => x"00",
          6741 => x"00",
          6742 => x"60",
          6743 => x"07",
          6744 => x"00",
          6745 => x"00",
          6746 => x"60",
          6747 => x"08",
          6748 => x"00",
          6749 => x"00",
          6750 => x"60",
          6751 => x"08",
          6752 => x"00",
          6753 => x"00",
          6754 => x"60",
          6755 => x"08",
          6756 => x"00",
          6757 => x"00",
          6758 => x"60",
          6759 => x"08",
          6760 => x"00",
          6761 => x"00",
          6762 => x"60",
          6763 => x"08",
          6764 => x"00",
          6765 => x"00",
          6766 => x"60",
          6767 => x"08",
          6768 => x"00",
          6769 => x"00",
        others => X"00"
    );

    shared variable RAM2 : ramArray :=
    (
             0 => x"0b",
             1 => x"0b",
             2 => x"8a",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"04",
            10 => x"84",
            11 => x"0b",
            12 => x"04",
            13 => x"84",
            14 => x"0b",
            15 => x"04",
            16 => x"84",
            17 => x"0b",
            18 => x"04",
            19 => x"84",
            20 => x"0b",
            21 => x"04",
            22 => x"85",
            23 => x"0b",
            24 => x"04",
            25 => x"85",
            26 => x"0b",
            27 => x"04",
            28 => x"85",
            29 => x"0b",
            30 => x"04",
            31 => x"85",
            32 => x"0b",
            33 => x"04",
            34 => x"86",
            35 => x"0b",
            36 => x"04",
            37 => x"86",
            38 => x"0b",
            39 => x"04",
            40 => x"86",
            41 => x"0b",
            42 => x"04",
            43 => x"86",
            44 => x"0b",
            45 => x"04",
            46 => x"87",
            47 => x"0b",
            48 => x"04",
            49 => x"87",
            50 => x"0b",
            51 => x"04",
            52 => x"87",
            53 => x"0b",
            54 => x"04",
            55 => x"87",
            56 => x"0b",
            57 => x"04",
            58 => x"88",
            59 => x"0b",
            60 => x"04",
            61 => x"88",
            62 => x"0b",
            63 => x"04",
            64 => x"88",
            65 => x"0b",
            66 => x"04",
            67 => x"88",
            68 => x"0b",
            69 => x"04",
            70 => x"89",
            71 => x"0b",
            72 => x"04",
            73 => x"89",
            74 => x"0b",
            75 => x"04",
            76 => x"89",
            77 => x"0b",
            78 => x"04",
            79 => x"89",
            80 => x"0b",
            81 => x"04",
            82 => x"8a",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"90",
           129 => x"91",
           130 => x"90",
           131 => x"91",
           132 => x"83",
           133 => x"91",
           134 => x"90",
           135 => x"91",
           136 => x"83",
           137 => x"91",
           138 => x"90",
           139 => x"91",
           140 => x"83",
           141 => x"91",
           142 => x"90",
           143 => x"91",
           144 => x"83",
           145 => x"91",
           146 => x"90",
           147 => x"91",
           148 => x"83",
           149 => x"91",
           150 => x"90",
           151 => x"91",
           152 => x"83",
           153 => x"91",
           154 => x"90",
           155 => x"91",
           156 => x"83",
           157 => x"91",
           158 => x"90",
           159 => x"91",
           160 => x"83",
           161 => x"91",
           162 => x"90",
           163 => x"91",
           164 => x"83",
           165 => x"91",
           166 => x"90",
           167 => x"91",
           168 => x"83",
           169 => x"91",
           170 => x"90",
           171 => x"91",
           172 => x"83",
           173 => x"91",
           174 => x"90",
           175 => x"91",
           176 => x"83",
           177 => x"91",
           178 => x"90",
           179 => x"91",
           180 => x"83",
           181 => x"91",
           182 => x"90",
           183 => x"91",
           184 => x"83",
           185 => x"91",
           186 => x"90",
           187 => x"91",
           188 => x"83",
           189 => x"91",
           190 => x"90",
           191 => x"91",
           192 => x"83",
           193 => x"91",
           194 => x"90",
           195 => x"91",
           196 => x"83",
           197 => x"91",
           198 => x"90",
           199 => x"91",
           200 => x"83",
           201 => x"91",
           202 => x"90",
           203 => x"91",
           204 => x"83",
           205 => x"91",
           206 => x"90",
           207 => x"91",
           208 => x"83",
           209 => x"91",
           210 => x"90",
           211 => x"91",
           212 => x"83",
           213 => x"91",
           214 => x"90",
           215 => x"91",
           216 => x"83",
           217 => x"91",
           218 => x"90",
           219 => x"91",
           220 => x"83",
           221 => x"91",
           222 => x"90",
           223 => x"91",
           224 => x"83",
           225 => x"91",
           226 => x"90",
           227 => x"91",
           228 => x"83",
           229 => x"91",
           230 => x"90",
           231 => x"91",
           232 => x"83",
           233 => x"91",
           234 => x"90",
           235 => x"91",
           236 => x"83",
           237 => x"91",
           238 => x"91",
           239 => x"91",
           240 => x"83",
           241 => x"91",
           242 => x"90",
           243 => x"91",
           244 => x"83",
           245 => x"91",
           246 => x"91",
           247 => x"91",
           248 => x"83",
           249 => x"91",
           250 => x"90",
           251 => x"91",
           252 => x"83",
           253 => x"91",
           254 => x"91",
           255 => x"91",
           256 => x"83",
           257 => x"91",
           258 => x"91",
           259 => x"91",
           260 => x"83",
           261 => x"91",
           262 => x"90",
           263 => x"91",
           264 => x"83",
           265 => x"91",
           266 => x"90",
           267 => x"91",
           268 => x"83",
           269 => x"91",
           270 => x"90",
           271 => x"91",
           272 => x"83",
           273 => x"91",
           274 => x"90",
           275 => x"91",
           276 => x"83",
           277 => x"91",
           278 => x"91",
           279 => x"91",
           280 => x"83",
           281 => x"91",
           282 => x"91",
           283 => x"91",
           284 => x"83",
           285 => x"91",
           286 => x"91",
           287 => x"91",
           288 => x"83",
           289 => x"91",
           290 => x"90",
           291 => x"91",
           292 => x"83",
           293 => x"91",
           294 => x"91",
           295 => x"91",
           296 => x"83",
           297 => x"91",
           298 => x"90",
           299 => x"91",
           300 => x"83",
           301 => x"91",
           302 => x"90",
           303 => x"91",
           304 => x"83",
           305 => x"91",
           306 => x"90",
           307 => x"91",
           308 => x"83",
           309 => x"91",
           310 => x"90",
           311 => x"91",
           312 => x"83",
           313 => x"91",
           314 => x"90",
           315 => x"91",
           316 => x"83",
           317 => x"91",
           318 => x"90",
           319 => x"91",
           320 => x"83",
           321 => x"91",
           322 => x"91",
           323 => x"91",
           324 => x"83",
           325 => x"91",
           326 => x"91",
           327 => x"8e",
           328 => x"70",
           329 => x"0c",
           330 => x"8a",
           331 => x"84",
           332 => x"af",
           333 => x"04",
           334 => x"08",
           335 => x"d4",
           336 => x"0d",
           337 => x"d3",
           338 => x"05",
           339 => x"d3",
           340 => x"05",
           341 => x"c5",
           342 => x"c8",
           343 => x"d3",
           344 => x"85",
           345 => x"d3",
           346 => x"91",
           347 => x"02",
           348 => x"0c",
           349 => x"81",
           350 => x"d4",
           351 => x"08",
           352 => x"d4",
           353 => x"08",
           354 => x"91",
           355 => x"70",
           356 => x"0c",
           357 => x"0d",
           358 => x"0c",
           359 => x"d4",
           360 => x"d3",
           361 => x"3d",
           362 => x"91",
           363 => x"fc",
           364 => x"0b",
           365 => x"08",
           366 => x"91",
           367 => x"8c",
           368 => x"d3",
           369 => x"05",
           370 => x"38",
           371 => x"08",
           372 => x"80",
           373 => x"80",
           374 => x"d4",
           375 => x"08",
           376 => x"91",
           377 => x"8c",
           378 => x"91",
           379 => x"8c",
           380 => x"d3",
           381 => x"05",
           382 => x"d3",
           383 => x"05",
           384 => x"39",
           385 => x"08",
           386 => x"80",
           387 => x"38",
           388 => x"08",
           389 => x"91",
           390 => x"88",
           391 => x"ad",
           392 => x"d4",
           393 => x"08",
           394 => x"08",
           395 => x"31",
           396 => x"08",
           397 => x"91",
           398 => x"f8",
           399 => x"d3",
           400 => x"05",
           401 => x"d3",
           402 => x"05",
           403 => x"d4",
           404 => x"08",
           405 => x"d3",
           406 => x"05",
           407 => x"d4",
           408 => x"08",
           409 => x"d3",
           410 => x"05",
           411 => x"39",
           412 => x"08",
           413 => x"80",
           414 => x"91",
           415 => x"88",
           416 => x"91",
           417 => x"f4",
           418 => x"91",
           419 => x"d4",
           420 => x"08",
           421 => x"d4",
           422 => x"0c",
           423 => x"d4",
           424 => x"08",
           425 => x"0c",
           426 => x"91",
           427 => x"04",
           428 => x"76",
           429 => x"8c",
           430 => x"33",
           431 => x"55",
           432 => x"8a",
           433 => x"06",
           434 => x"2e",
           435 => x"12",
           436 => x"2e",
           437 => x"73",
           438 => x"55",
           439 => x"52",
           440 => x"09",
           441 => x"38",
           442 => x"c8",
           443 => x"0d",
           444 => x"88",
           445 => x"70",
           446 => x"07",
           447 => x"8f",
           448 => x"38",
           449 => x"84",
           450 => x"72",
           451 => x"05",
           452 => x"71",
           453 => x"53",
           454 => x"70",
           455 => x"0c",
           456 => x"71",
           457 => x"38",
           458 => x"90",
           459 => x"70",
           460 => x"0c",
           461 => x"71",
           462 => x"38",
           463 => x"8e",
           464 => x"0d",
           465 => x"72",
           466 => x"53",
           467 => x"93",
           468 => x"73",
           469 => x"54",
           470 => x"2e",
           471 => x"73",
           472 => x"71",
           473 => x"ff",
           474 => x"70",
           475 => x"38",
           476 => x"70",
           477 => x"81",
           478 => x"81",
           479 => x"71",
           480 => x"ff",
           481 => x"54",
           482 => x"38",
           483 => x"73",
           484 => x"75",
           485 => x"71",
           486 => x"d3",
           487 => x"52",
           488 => x"04",
           489 => x"f7",
           490 => x"14",
           491 => x"84",
           492 => x"06",
           493 => x"70",
           494 => x"14",
           495 => x"08",
           496 => x"71",
           497 => x"dc",
           498 => x"54",
           499 => x"39",
           500 => x"d3",
           501 => x"3d",
           502 => x"3d",
           503 => x"54",
           504 => x"2b",
           505 => x"3f",
           506 => x"08",
           507 => x"72",
           508 => x"54",
           509 => x"25",
           510 => x"91",
           511 => x"84",
           512 => x"fc",
           513 => x"70",
           514 => x"55",
           515 => x"2e",
           516 => x"73",
           517 => x"a0",
           518 => x"06",
           519 => x"14",
           520 => x"54",
           521 => x"f6",
           522 => x"84",
           523 => x"52",
           524 => x"52",
           525 => x"2e",
           526 => x"53",
           527 => x"9f",
           528 => x"51",
           529 => x"38",
           530 => x"70",
           531 => x"81",
           532 => x"80",
           533 => x"05",
           534 => x"75",
           535 => x"70",
           536 => x"0c",
           537 => x"04",
           538 => x"76",
           539 => x"80",
           540 => x"86",
           541 => x"52",
           542 => x"c4",
           543 => x"c8",
           544 => x"80",
           545 => x"74",
           546 => x"d3",
           547 => x"3d",
           548 => x"3d",
           549 => x"11",
           550 => x"5b",
           551 => x"79",
           552 => x"bf",
           553 => x"33",
           554 => x"82",
           555 => x"26",
           556 => x"84",
           557 => x"83",
           558 => x"26",
           559 => x"85",
           560 => x"84",
           561 => x"26",
           562 => x"86",
           563 => x"85",
           564 => x"26",
           565 => x"88",
           566 => x"86",
           567 => x"e7",
           568 => x"38",
           569 => x"5a",
           570 => x"87",
           571 => x"f3",
           572 => x"22",
           573 => x"22",
           574 => x"33",
           575 => x"33",
           576 => x"33",
           577 => x"33",
           578 => x"33",
           579 => x"52",
           580 => x"51",
           581 => x"87",
           582 => x"5b",
           583 => x"7b",
           584 => x"98",
           585 => x"1c",
           586 => x"98",
           587 => x"1c",
           588 => x"98",
           589 => x"1c",
           590 => x"98",
           591 => x"1c",
           592 => x"98",
           593 => x"1c",
           594 => x"98",
           595 => x"1c",
           596 => x"98",
           597 => x"1c",
           598 => x"98",
           599 => x"7b",
           600 => x"7a",
           601 => x"0c",
           602 => x"04",
           603 => x"7d",
           604 => x"98",
           605 => x"7c",
           606 => x"98",
           607 => x"7a",
           608 => x"c0",
           609 => x"5b",
           610 => x"34",
           611 => x"b4",
           612 => x"83",
           613 => x"c0",
           614 => x"5b",
           615 => x"34",
           616 => x"ac",
           617 => x"85",
           618 => x"c0",
           619 => x"5b",
           620 => x"34",
           621 => x"a4",
           622 => x"88",
           623 => x"c0",
           624 => x"5b",
           625 => x"23",
           626 => x"8a",
           627 => x"88",
           628 => x"86",
           629 => x"85",
           630 => x"84",
           631 => x"83",
           632 => x"82",
           633 => x"79",
           634 => x"b6",
           635 => x"af",
           636 => x"0d",
           637 => x"0d",
           638 => x"33",
           639 => x"9f",
           640 => x"51",
           641 => x"91",
           642 => x"82",
           643 => x"fd",
           644 => x"0b",
           645 => x"c0",
           646 => x"87",
           647 => x"51",
           648 => x"86",
           649 => x"94",
           650 => x"08",
           651 => x"70",
           652 => x"52",
           653 => x"2e",
           654 => x"91",
           655 => x"06",
           656 => x"d7",
           657 => x"2a",
           658 => x"81",
           659 => x"70",
           660 => x"38",
           661 => x"70",
           662 => x"51",
           663 => x"38",
           664 => x"cb",
           665 => x"87",
           666 => x"52",
           667 => x"86",
           668 => x"94",
           669 => x"72",
           670 => x"d3",
           671 => x"3d",
           672 => x"3d",
           673 => x"05",
           674 => x"91",
           675 => x"54",
           676 => x"94",
           677 => x"80",
           678 => x"87",
           679 => x"51",
           680 => x"96",
           681 => x"06",
           682 => x"70",
           683 => x"38",
           684 => x"70",
           685 => x"51",
           686 => x"71",
           687 => x"32",
           688 => x"51",
           689 => x"2e",
           690 => x"93",
           691 => x"06",
           692 => x"ff",
           693 => x"0b",
           694 => x"33",
           695 => x"94",
           696 => x"80",
           697 => x"87",
           698 => x"52",
           699 => x"85",
           700 => x"fb",
           701 => x"54",
           702 => x"52",
           703 => x"2e",
           704 => x"73",
           705 => x"55",
           706 => x"91",
           707 => x"54",
           708 => x"94",
           709 => x"80",
           710 => x"87",
           711 => x"51",
           712 => x"96",
           713 => x"06",
           714 => x"70",
           715 => x"38",
           716 => x"70",
           717 => x"51",
           718 => x"71",
           719 => x"32",
           720 => x"51",
           721 => x"2e",
           722 => x"93",
           723 => x"06",
           724 => x"ff",
           725 => x"0b",
           726 => x"33",
           727 => x"94",
           728 => x"80",
           729 => x"87",
           730 => x"52",
           731 => x"81",
           732 => x"52",
           733 => x"8b",
           734 => x"d3",
           735 => x"3d",
           736 => x"3d",
           737 => x"91",
           738 => x"52",
           739 => x"84",
           740 => x"2e",
           741 => x"c0",
           742 => x"70",
           743 => x"2a",
           744 => x"51",
           745 => x"80",
           746 => x"0b",
           747 => x"c0",
           748 => x"c0",
           749 => x"70",
           750 => x"38",
           751 => x"90",
           752 => x"70",
           753 => x"91",
           754 => x"51",
           755 => x"04",
           756 => x"0b",
           757 => x"c0",
           758 => x"c0",
           759 => x"70",
           760 => x"38",
           761 => x"94",
           762 => x"70",
           763 => x"81",
           764 => x"51",
           765 => x"80",
           766 => x"0b",
           767 => x"c0",
           768 => x"c0",
           769 => x"70",
           770 => x"38",
           771 => x"90",
           772 => x"70",
           773 => x"98",
           774 => x"51",
           775 => x"c8",
           776 => x"0d",
           777 => x"0d",
           778 => x"80",
           779 => x"9c",
           780 => x"51",
           781 => x"80",
           782 => x"38",
           783 => x"0b",
           784 => x"9c",
           785 => x"84",
           786 => x"9e",
           787 => x"0c",
           788 => x"87",
           789 => x"08",
           790 => x"8c",
           791 => x"9e",
           792 => x"0c",
           793 => x"87",
           794 => x"08",
           795 => x"94",
           796 => x"9e",
           797 => x"0c",
           798 => x"87",
           799 => x"08",
           800 => x"9c",
           801 => x"9e",
           802 => x"0c",
           803 => x"87",
           804 => x"08",
           805 => x"73",
           806 => x"70",
           807 => x"a8",
           808 => x"9e",
           809 => x"0c",
           810 => x"ac",
           811 => x"12",
           812 => x"87",
           813 => x"08",
           814 => x"06",
           815 => x"70",
           816 => x"38",
           817 => x"72",
           818 => x"87",
           819 => x"08",
           820 => x"80",
           821 => x"52",
           822 => x"83",
           823 => x"71",
           824 => x"34",
           825 => x"c0",
           826 => x"70",
           827 => x"06",
           828 => x"70",
           829 => x"38",
           830 => x"91",
           831 => x"80",
           832 => x"9e",
           833 => x"90",
           834 => x"52",
           835 => x"2e",
           836 => x"52",
           837 => x"f4",
           838 => x"87",
           839 => x"08",
           840 => x"06",
           841 => x"70",
           842 => x"38",
           843 => x"91",
           844 => x"80",
           845 => x"9e",
           846 => x"84",
           847 => x"52",
           848 => x"2e",
           849 => x"52",
           850 => x"f6",
           851 => x"87",
           852 => x"08",
           853 => x"06",
           854 => x"70",
           855 => x"38",
           856 => x"91",
           857 => x"80",
           858 => x"9e",
           859 => x"81",
           860 => x"52",
           861 => x"2e",
           862 => x"52",
           863 => x"f8",
           864 => x"f9",
           865 => x"9e",
           866 => x"70",
           867 => x"70",
           868 => x"51",
           869 => x"72",
           870 => x"54",
           871 => x"80",
           872 => x"90",
           873 => x"52",
           874 => x"83",
           875 => x"71",
           876 => x"0b",
           877 => x"88",
           878 => x"06",
           879 => x"70",
           880 => x"38",
           881 => x"91",
           882 => x"87",
           883 => x"08",
           884 => x"51",
           885 => x"cb",
           886 => x"3d",
           887 => x"3d",
           888 => x"c0",
           889 => x"3f",
           890 => x"33",
           891 => x"2e",
           892 => x"b6",
           893 => x"ad",
           894 => x"e8",
           895 => x"3f",
           896 => x"70",
           897 => x"73",
           898 => x"38",
           899 => x"53",
           900 => x"08",
           901 => x"80",
           902 => x"3f",
           903 => x"70",
           904 => x"73",
           905 => x"38",
           906 => x"53",
           907 => x"52",
           908 => x"51",
           909 => x"91",
           910 => x"33",
           911 => x"8a",
           912 => x"33",
           913 => x"2e",
           914 => x"cb",
           915 => x"54",
           916 => x"53",
           917 => x"cc",
           918 => x"3f",
           919 => x"33",
           920 => x"2e",
           921 => x"b7",
           922 => x"b9",
           923 => x"f6",
           924 => x"80",
           925 => x"91",
           926 => x"83",
           927 => x"cb",
           928 => x"73",
           929 => x"38",
           930 => x"51",
           931 => x"91",
           932 => x"33",
           933 => x"80",
           934 => x"81",
           935 => x"91",
           936 => x"88",
           937 => x"cb",
           938 => x"73",
           939 => x"38",
           940 => x"51",
           941 => x"91",
           942 => x"33",
           943 => x"80",
           944 => x"81",
           945 => x"91",
           946 => x"88",
           947 => x"b8",
           948 => x"d1",
           949 => x"dc",
           950 => x"84",
           951 => x"54",
           952 => x"53",
           953 => x"b7",
           954 => x"52",
           955 => x"51",
           956 => x"88",
           957 => x"91",
           958 => x"88",
           959 => x"15",
           960 => x"b9",
           961 => x"97",
           962 => x"08",
           963 => x"98",
           964 => x"3f",
           965 => x"04",
           966 => x"02",
           967 => x"52",
           968 => x"bb",
           969 => x"10",
           970 => x"b0",
           971 => x"71",
           972 => x"ba",
           973 => x"bb",
           974 => x"91",
           975 => x"f7",
           976 => x"39",
           977 => x"51",
           978 => x"9a",
           979 => x"d8",
           980 => x"3f",
           981 => x"ba",
           982 => x"97",
           983 => x"91",
           984 => x"f7",
           985 => x"3d",
           986 => x"88",
           987 => x"80",
           988 => x"96",
           989 => x"ff",
           990 => x"c0",
           991 => x"08",
           992 => x"72",
           993 => x"07",
           994 => x"80",
           995 => x"83",
           996 => x"ff",
           997 => x"c0",
           998 => x"08",
           999 => x"0c",
          1000 => x"0c",
          1001 => x"91",
          1002 => x"06",
          1003 => x"80",
          1004 => x"51",
          1005 => x"04",
          1006 => x"08",
          1007 => x"84",
          1008 => x"3d",
          1009 => x"05",
          1010 => x"8a",
          1011 => x"06",
          1012 => x"51",
          1013 => x"d3",
          1014 => x"2e",
          1015 => x"d3",
          1016 => x"72",
          1017 => x"d3",
          1018 => x"05",
          1019 => x"0c",
          1020 => x"d3",
          1021 => x"2e",
          1022 => x"51",
          1023 => x"08",
          1024 => x"84",
          1025 => x"fe",
          1026 => x"97",
          1027 => x"d3",
          1028 => x"91",
          1029 => x"54",
          1030 => x"3f",
          1031 => x"d8",
          1032 => x"0d",
          1033 => x"0d",
          1034 => x"53",
          1035 => x"2e",
          1036 => x"70",
          1037 => x"33",
          1038 => x"3f",
          1039 => x"71",
          1040 => x"3d",
          1041 => x"3d",
          1042 => x"d3",
          1043 => x"91",
          1044 => x"71",
          1045 => x"53",
          1046 => x"91",
          1047 => x"81",
          1048 => x"51",
          1049 => x"72",
          1050 => x"f1",
          1051 => x"d3",
          1052 => x"3d",
          1053 => x"3d",
          1054 => x"5d",
          1055 => x"81",
          1056 => x"56",
          1057 => x"85",
          1058 => x"a5",
          1059 => x"75",
          1060 => x"3f",
          1061 => x"70",
          1062 => x"05",
          1063 => x"5e",
          1064 => x"2e",
          1065 => x"8c",
          1066 => x"70",
          1067 => x"33",
          1068 => x"39",
          1069 => x"09",
          1070 => x"38",
          1071 => x"81",
          1072 => x"57",
          1073 => x"2e",
          1074 => x"92",
          1075 => x"1d",
          1076 => x"70",
          1077 => x"33",
          1078 => x"53",
          1079 => x"16",
          1080 => x"26",
          1081 => x"8a",
          1082 => x"05",
          1083 => x"05",
          1084 => x"11",
          1085 => x"89",
          1086 => x"38",
          1087 => x"32",
          1088 => x"72",
          1089 => x"78",
          1090 => x"70",
          1091 => x"07",
          1092 => x"07",
          1093 => x"52",
          1094 => x"80",
          1095 => x"7c",
          1096 => x"70",
          1097 => x"33",
          1098 => x"80",
          1099 => x"38",
          1100 => x"e0",
          1101 => x"38",
          1102 => x"81",
          1103 => x"53",
          1104 => x"53",
          1105 => x"81",
          1106 => x"10",
          1107 => x"dc",
          1108 => x"08",
          1109 => x"1d",
          1110 => x"5d",
          1111 => x"33",
          1112 => x"74",
          1113 => x"81",
          1114 => x"70",
          1115 => x"54",
          1116 => x"7c",
          1117 => x"81",
          1118 => x"72",
          1119 => x"81",
          1120 => x"72",
          1121 => x"38",
          1122 => x"81",
          1123 => x"51",
          1124 => x"75",
          1125 => x"81",
          1126 => x"79",
          1127 => x"38",
          1128 => x"81",
          1129 => x"15",
          1130 => x"7a",
          1131 => x"38",
          1132 => x"8e",
          1133 => x"15",
          1134 => x"73",
          1135 => x"fd",
          1136 => x"84",
          1137 => x"33",
          1138 => x"fb",
          1139 => x"ad",
          1140 => x"95",
          1141 => x"91",
          1142 => x"8d",
          1143 => x"89",
          1144 => x"fb",
          1145 => x"95",
          1146 => x"2a",
          1147 => x"51",
          1148 => x"2e",
          1149 => x"84",
          1150 => x"59",
          1151 => x"39",
          1152 => x"2e",
          1153 => x"8b",
          1154 => x"1d",
          1155 => x"5d",
          1156 => x"7b",
          1157 => x"08",
          1158 => x"74",
          1159 => x"70",
          1160 => x"07",
          1161 => x"80",
          1162 => x"51",
          1163 => x"72",
          1164 => x"38",
          1165 => x"90",
          1166 => x"80",
          1167 => x"76",
          1168 => x"3f",
          1169 => x"08",
          1170 => x"7b",
          1171 => x"55",
          1172 => x"91",
          1173 => x"57",
          1174 => x"99",
          1175 => x"16",
          1176 => x"06",
          1177 => x"75",
          1178 => x"89",
          1179 => x"70",
          1180 => x"56",
          1181 => x"78",
          1182 => x"b0",
          1183 => x"72",
          1184 => x"18",
          1185 => x"79",
          1186 => x"70",
          1187 => x"06",
          1188 => x"58",
          1189 => x"38",
          1190 => x"70",
          1191 => x"53",
          1192 => x"8e",
          1193 => x"78",
          1194 => x"53",
          1195 => x"81",
          1196 => x"7d",
          1197 => x"54",
          1198 => x"83",
          1199 => x"7c",
          1200 => x"81",
          1201 => x"72",
          1202 => x"81",
          1203 => x"72",
          1204 => x"38",
          1205 => x"81",
          1206 => x"51",
          1207 => x"75",
          1208 => x"81",
          1209 => x"79",
          1210 => x"38",
          1211 => x"3d",
          1212 => x"70",
          1213 => x"58",
          1214 => x"77",
          1215 => x"81",
          1216 => x"72",
          1217 => x"f5",
          1218 => x"f9",
          1219 => x"81",
          1220 => x"79",
          1221 => x"38",
          1222 => x"96",
          1223 => x"fd",
          1224 => x"3d",
          1225 => x"05",
          1226 => x"52",
          1227 => x"c6",
          1228 => x"0d",
          1229 => x"0d",
          1230 => x"e0",
          1231 => x"88",
          1232 => x"51",
          1233 => x"91",
          1234 => x"53",
          1235 => x"80",
          1236 => x"e0",
          1237 => x"0d",
          1238 => x"0d",
          1239 => x"08",
          1240 => x"d8",
          1241 => x"88",
          1242 => x"52",
          1243 => x"3f",
          1244 => x"d8",
          1245 => x"0d",
          1246 => x"0d",
          1247 => x"57",
          1248 => x"d3",
          1249 => x"2e",
          1250 => x"86",
          1251 => x"80",
          1252 => x"55",
          1253 => x"08",
          1254 => x"91",
          1255 => x"81",
          1256 => x"73",
          1257 => x"38",
          1258 => x"80",
          1259 => x"88",
          1260 => x"76",
          1261 => x"07",
          1262 => x"80",
          1263 => x"54",
          1264 => x"80",
          1265 => x"ff",
          1266 => x"ff",
          1267 => x"f7",
          1268 => x"39",
          1269 => x"ff",
          1270 => x"16",
          1271 => x"25",
          1272 => x"76",
          1273 => x"72",
          1274 => x"74",
          1275 => x"52",
          1276 => x"3f",
          1277 => x"74",
          1278 => x"72",
          1279 => x"f7",
          1280 => x"53",
          1281 => x"c8",
          1282 => x"0d",
          1283 => x"0d",
          1284 => x"08",
          1285 => x"dc",
          1286 => x"76",
          1287 => x"d9",
          1288 => x"d3",
          1289 => x"3d",
          1290 => x"3d",
          1291 => x"5a",
          1292 => x"7a",
          1293 => x"70",
          1294 => x"58",
          1295 => x"09",
          1296 => x"38",
          1297 => x"05",
          1298 => x"08",
          1299 => x"53",
          1300 => x"f0",
          1301 => x"2e",
          1302 => x"8e",
          1303 => x"08",
          1304 => x"75",
          1305 => x"56",
          1306 => x"b0",
          1307 => x"06",
          1308 => x"74",
          1309 => x"75",
          1310 => x"70",
          1311 => x"73",
          1312 => x"9a",
          1313 => x"f8",
          1314 => x"06",
          1315 => x"0b",
          1316 => x"0c",
          1317 => x"33",
          1318 => x"80",
          1319 => x"75",
          1320 => x"76",
          1321 => x"70",
          1322 => x"57",
          1323 => x"56",
          1324 => x"81",
          1325 => x"14",
          1326 => x"88",
          1327 => x"27",
          1328 => x"f3",
          1329 => x"53",
          1330 => x"89",
          1331 => x"38",
          1332 => x"56",
          1333 => x"80",
          1334 => x"39",
          1335 => x"56",
          1336 => x"80",
          1337 => x"e0",
          1338 => x"38",
          1339 => x"81",
          1340 => x"53",
          1341 => x"81",
          1342 => x"53",
          1343 => x"8e",
          1344 => x"70",
          1345 => x"55",
          1346 => x"27",
          1347 => x"77",
          1348 => x"76",
          1349 => x"75",
          1350 => x"76",
          1351 => x"70",
          1352 => x"56",
          1353 => x"ff",
          1354 => x"80",
          1355 => x"75",
          1356 => x"79",
          1357 => x"75",
          1358 => x"0c",
          1359 => x"04",
          1360 => x"7a",
          1361 => x"80",
          1362 => x"75",
          1363 => x"56",
          1364 => x"a0",
          1365 => x"06",
          1366 => x"08",
          1367 => x"0c",
          1368 => x"33",
          1369 => x"a0",
          1370 => x"73",
          1371 => x"81",
          1372 => x"81",
          1373 => x"76",
          1374 => x"70",
          1375 => x"58",
          1376 => x"09",
          1377 => x"d3",
          1378 => x"81",
          1379 => x"74",
          1380 => x"55",
          1381 => x"e2",
          1382 => x"73",
          1383 => x"09",
          1384 => x"38",
          1385 => x"14",
          1386 => x"08",
          1387 => x"54",
          1388 => x"39",
          1389 => x"81",
          1390 => x"75",
          1391 => x"56",
          1392 => x"39",
          1393 => x"74",
          1394 => x"38",
          1395 => x"80",
          1396 => x"89",
          1397 => x"38",
          1398 => x"d0",
          1399 => x"56",
          1400 => x"80",
          1401 => x"39",
          1402 => x"e1",
          1403 => x"80",
          1404 => x"57",
          1405 => x"74",
          1406 => x"38",
          1407 => x"27",
          1408 => x"14",
          1409 => x"06",
          1410 => x"14",
          1411 => x"06",
          1412 => x"74",
          1413 => x"f9",
          1414 => x"ff",
          1415 => x"89",
          1416 => x"38",
          1417 => x"c5",
          1418 => x"29",
          1419 => x"81",
          1420 => x"75",
          1421 => x"56",
          1422 => x"a0",
          1423 => x"38",
          1424 => x"84",
          1425 => x"56",
          1426 => x"81",
          1427 => x"d3",
          1428 => x"3d",
          1429 => x"3d",
          1430 => x"05",
          1431 => x"52",
          1432 => x"87",
          1433 => x"84",
          1434 => x"71",
          1435 => x"0c",
          1436 => x"04",
          1437 => x"02",
          1438 => x"02",
          1439 => x"05",
          1440 => x"83",
          1441 => x"26",
          1442 => x"72",
          1443 => x"c0",
          1444 => x"51",
          1445 => x"80",
          1446 => x"81",
          1447 => x"71",
          1448 => x"29",
          1449 => x"8c",
          1450 => x"71",
          1451 => x"87",
          1452 => x"0c",
          1453 => x"c0",
          1454 => x"71",
          1455 => x"06",
          1456 => x"80",
          1457 => x"73",
          1458 => x"ef",
          1459 => x"29",
          1460 => x"8c",
          1461 => x"fc",
          1462 => x"53",
          1463 => x"38",
          1464 => x"8c",
          1465 => x"80",
          1466 => x"71",
          1467 => x"14",
          1468 => x"84",
          1469 => x"70",
          1470 => x"0c",
          1471 => x"04",
          1472 => x"61",
          1473 => x"8c",
          1474 => x"05",
          1475 => x"5d",
          1476 => x"52",
          1477 => x"3f",
          1478 => x"08",
          1479 => x"55",
          1480 => x"ac",
          1481 => x"58",
          1482 => x"98",
          1483 => x"2b",
          1484 => x"8c",
          1485 => x"92",
          1486 => x"42",
          1487 => x"56",
          1488 => x"87",
          1489 => x"1a",
          1490 => x"52",
          1491 => x"74",
          1492 => x"2a",
          1493 => x"51",
          1494 => x"80",
          1495 => x"78",
          1496 => x"78",
          1497 => x"5a",
          1498 => x"57",
          1499 => x"52",
          1500 => x"87",
          1501 => x"52",
          1502 => x"75",
          1503 => x"80",
          1504 => x"76",
          1505 => x"99",
          1506 => x"0c",
          1507 => x"8c",
          1508 => x"08",
          1509 => x"51",
          1510 => x"38",
          1511 => x"8d",
          1512 => x"1c",
          1513 => x"81",
          1514 => x"53",
          1515 => x"2e",
          1516 => x"fc",
          1517 => x"52",
          1518 => x"7e",
          1519 => x"80",
          1520 => x"80",
          1521 => x"71",
          1522 => x"38",
          1523 => x"54",
          1524 => x"c8",
          1525 => x"0d",
          1526 => x"0d",
          1527 => x"02",
          1528 => x"05",
          1529 => x"5c",
          1530 => x"52",
          1531 => x"3f",
          1532 => x"08",
          1533 => x"55",
          1534 => x"ae",
          1535 => x"87",
          1536 => x"73",
          1537 => x"c0",
          1538 => x"87",
          1539 => x"12",
          1540 => x"57",
          1541 => x"76",
          1542 => x"92",
          1543 => x"71",
          1544 => x"75",
          1545 => x"74",
          1546 => x"2a",
          1547 => x"51",
          1548 => x"80",
          1549 => x"76",
          1550 => x"58",
          1551 => x"81",
          1552 => x"81",
          1553 => x"06",
          1554 => x"80",
          1555 => x"75",
          1556 => x"d3",
          1557 => x"52",
          1558 => x"87",
          1559 => x"80",
          1560 => x"81",
          1561 => x"c0",
          1562 => x"53",
          1563 => x"82",
          1564 => x"71",
          1565 => x"1a",
          1566 => x"81",
          1567 => x"ff",
          1568 => x"1d",
          1569 => x"79",
          1570 => x"38",
          1571 => x"80",
          1572 => x"87",
          1573 => x"26",
          1574 => x"73",
          1575 => x"06",
          1576 => x"2e",
          1577 => x"52",
          1578 => x"91",
          1579 => x"8f",
          1580 => x"f7",
          1581 => x"02",
          1582 => x"05",
          1583 => x"05",
          1584 => x"71",
          1585 => x"56",
          1586 => x"91",
          1587 => x"81",
          1588 => x"54",
          1589 => x"81",
          1590 => x"2e",
          1591 => x"74",
          1592 => x"72",
          1593 => x"38",
          1594 => x"83",
          1595 => x"a0",
          1596 => x"29",
          1597 => x"8c",
          1598 => x"51",
          1599 => x"88",
          1600 => x"0c",
          1601 => x"39",
          1602 => x"0c",
          1603 => x"39",
          1604 => x"91",
          1605 => x"8b",
          1606 => x"ff",
          1607 => x"70",
          1608 => x"33",
          1609 => x"72",
          1610 => x"c8",
          1611 => x"52",
          1612 => x"04",
          1613 => x"75",
          1614 => x"82",
          1615 => x"90",
          1616 => x"2b",
          1617 => x"33",
          1618 => x"33",
          1619 => x"07",
          1620 => x"0c",
          1621 => x"54",
          1622 => x"0d",
          1623 => x"0d",
          1624 => x"05",
          1625 => x"52",
          1626 => x"70",
          1627 => x"34",
          1628 => x"51",
          1629 => x"83",
          1630 => x"ff",
          1631 => x"75",
          1632 => x"72",
          1633 => x"54",
          1634 => x"2a",
          1635 => x"70",
          1636 => x"34",
          1637 => x"51",
          1638 => x"81",
          1639 => x"70",
          1640 => x"70",
          1641 => x"3d",
          1642 => x"3d",
          1643 => x"77",
          1644 => x"70",
          1645 => x"38",
          1646 => x"05",
          1647 => x"70",
          1648 => x"34",
          1649 => x"70",
          1650 => x"3d",
          1651 => x"3d",
          1652 => x"76",
          1653 => x"72",
          1654 => x"05",
          1655 => x"11",
          1656 => x"38",
          1657 => x"04",
          1658 => x"78",
          1659 => x"56",
          1660 => x"81",
          1661 => x"74",
          1662 => x"56",
          1663 => x"31",
          1664 => x"52",
          1665 => x"80",
          1666 => x"71",
          1667 => x"38",
          1668 => x"c8",
          1669 => x"0d",
          1670 => x"0d",
          1671 => x"33",
          1672 => x"70",
          1673 => x"38",
          1674 => x"94",
          1675 => x"70",
          1676 => x"70",
          1677 => x"38",
          1678 => x"09",
          1679 => x"38",
          1680 => x"d3",
          1681 => x"3d",
          1682 => x"0b",
          1683 => x"0c",
          1684 => x"91",
          1685 => x"04",
          1686 => x"79",
          1687 => x"83",
          1688 => x"58",
          1689 => x"80",
          1690 => x"54",
          1691 => x"53",
          1692 => x"53",
          1693 => x"52",
          1694 => x"3f",
          1695 => x"08",
          1696 => x"81",
          1697 => x"91",
          1698 => x"83",
          1699 => x"16",
          1700 => x"08",
          1701 => x"9c",
          1702 => x"a4",
          1703 => x"33",
          1704 => x"2e",
          1705 => x"98",
          1706 => x"b0",
          1707 => x"17",
          1708 => x"76",
          1709 => x"33",
          1710 => x"3f",
          1711 => x"58",
          1712 => x"c8",
          1713 => x"0d",
          1714 => x"0d",
          1715 => x"57",
          1716 => x"17",
          1717 => x"af",
          1718 => x"fe",
          1719 => x"d3",
          1720 => x"91",
          1721 => x"9f",
          1722 => x"74",
          1723 => x"52",
          1724 => x"51",
          1725 => x"91",
          1726 => x"80",
          1727 => x"ff",
          1728 => x"74",
          1729 => x"75",
          1730 => x"0c",
          1731 => x"04",
          1732 => x"7a",
          1733 => x"fe",
          1734 => x"d3",
          1735 => x"91",
          1736 => x"81",
          1737 => x"33",
          1738 => x"2e",
          1739 => x"80",
          1740 => x"17",
          1741 => x"81",
          1742 => x"06",
          1743 => x"84",
          1744 => x"d3",
          1745 => x"b4",
          1746 => x"56",
          1747 => x"82",
          1748 => x"84",
          1749 => x"fc",
          1750 => x"8b",
          1751 => x"52",
          1752 => x"97",
          1753 => x"85",
          1754 => x"84",
          1755 => x"fc",
          1756 => x"17",
          1757 => x"9c",
          1758 => x"ff",
          1759 => x"08",
          1760 => x"17",
          1761 => x"3f",
          1762 => x"81",
          1763 => x"19",
          1764 => x"53",
          1765 => x"17",
          1766 => x"bd",
          1767 => x"18",
          1768 => x"80",
          1769 => x"33",
          1770 => x"3f",
          1771 => x"08",
          1772 => x"38",
          1773 => x"91",
          1774 => x"8a",
          1775 => x"fb",
          1776 => x"fe",
          1777 => x"08",
          1778 => x"56",
          1779 => x"74",
          1780 => x"38",
          1781 => x"70",
          1782 => x"16",
          1783 => x"53",
          1784 => x"c8",
          1785 => x"0d",
          1786 => x"0d",
          1787 => x"08",
          1788 => x"81",
          1789 => x"38",
          1790 => x"75",
          1791 => x"81",
          1792 => x"39",
          1793 => x"54",
          1794 => x"2e",
          1795 => x"72",
          1796 => x"38",
          1797 => x"8d",
          1798 => x"39",
          1799 => x"81",
          1800 => x"b6",
          1801 => x"2a",
          1802 => x"2a",
          1803 => x"05",
          1804 => x"57",
          1805 => x"91",
          1806 => x"81",
          1807 => x"83",
          1808 => x"b4",
          1809 => x"19",
          1810 => x"a4",
          1811 => x"55",
          1812 => x"59",
          1813 => x"3f",
          1814 => x"08",
          1815 => x"76",
          1816 => x"14",
          1817 => x"70",
          1818 => x"07",
          1819 => x"71",
          1820 => x"52",
          1821 => x"72",
          1822 => x"77",
          1823 => x"56",
          1824 => x"74",
          1825 => x"15",
          1826 => x"73",
          1827 => x"3f",
          1828 => x"08",
          1829 => x"74",
          1830 => x"06",
          1831 => x"05",
          1832 => x"3f",
          1833 => x"08",
          1834 => x"06",
          1835 => x"74",
          1836 => x"15",
          1837 => x"73",
          1838 => x"3f",
          1839 => x"08",
          1840 => x"82",
          1841 => x"06",
          1842 => x"05",
          1843 => x"3f",
          1844 => x"08",
          1845 => x"56",
          1846 => x"56",
          1847 => x"c8",
          1848 => x"0d",
          1849 => x"0d",
          1850 => x"58",
          1851 => x"57",
          1852 => x"82",
          1853 => x"98",
          1854 => x"82",
          1855 => x"33",
          1856 => x"2e",
          1857 => x"72",
          1858 => x"38",
          1859 => x"8d",
          1860 => x"39",
          1861 => x"81",
          1862 => x"88",
          1863 => x"2a",
          1864 => x"2a",
          1865 => x"05",
          1866 => x"59",
          1867 => x"91",
          1868 => x"57",
          1869 => x"08",
          1870 => x"78",
          1871 => x"15",
          1872 => x"1b",
          1873 => x"56",
          1874 => x"75",
          1875 => x"2e",
          1876 => x"84",
          1877 => x"06",
          1878 => x"06",
          1879 => x"53",
          1880 => x"81",
          1881 => x"34",
          1882 => x"a4",
          1883 => x"52",
          1884 => x"d5",
          1885 => x"c8",
          1886 => x"d3",
          1887 => x"a4",
          1888 => x"ff",
          1889 => x"11",
          1890 => x"78",
          1891 => x"55",
          1892 => x"8f",
          1893 => x"2a",
          1894 => x"8f",
          1895 => x"f0",
          1896 => x"73",
          1897 => x"0b",
          1898 => x"80",
          1899 => x"88",
          1900 => x"08",
          1901 => x"51",
          1902 => x"91",
          1903 => x"57",
          1904 => x"08",
          1905 => x"75",
          1906 => x"06",
          1907 => x"83",
          1908 => x"05",
          1909 => x"f7",
          1910 => x"0b",
          1911 => x"80",
          1912 => x"87",
          1913 => x"08",
          1914 => x"51",
          1915 => x"91",
          1916 => x"57",
          1917 => x"08",
          1918 => x"f0",
          1919 => x"82",
          1920 => x"06",
          1921 => x"05",
          1922 => x"54",
          1923 => x"3f",
          1924 => x"08",
          1925 => x"76",
          1926 => x"51",
          1927 => x"81",
          1928 => x"34",
          1929 => x"c8",
          1930 => x"0d",
          1931 => x"0d",
          1932 => x"72",
          1933 => x"55",
          1934 => x"27",
          1935 => x"15",
          1936 => x"86",
          1937 => x"81",
          1938 => x"80",
          1939 => x"ff",
          1940 => x"74",
          1941 => x"3f",
          1942 => x"08",
          1943 => x"c8",
          1944 => x"38",
          1945 => x"56",
          1946 => x"81",
          1947 => x"39",
          1948 => x"08",
          1949 => x"39",
          1950 => x"51",
          1951 => x"91",
          1952 => x"56",
          1953 => x"08",
          1954 => x"c9",
          1955 => x"c8",
          1956 => x"d2",
          1957 => x"c8",
          1958 => x"cf",
          1959 => x"73",
          1960 => x"fc",
          1961 => x"d3",
          1962 => x"38",
          1963 => x"fe",
          1964 => x"15",
          1965 => x"93",
          1966 => x"08",
          1967 => x"16",
          1968 => x"33",
          1969 => x"73",
          1970 => x"75",
          1971 => x"08",
          1972 => x"a4",
          1973 => x"75",
          1974 => x"0c",
          1975 => x"04",
          1976 => x"7d",
          1977 => x"5b",
          1978 => x"95",
          1979 => x"08",
          1980 => x"2e",
          1981 => x"19",
          1982 => x"b7",
          1983 => x"b3",
          1984 => x"7b",
          1985 => x"3f",
          1986 => x"91",
          1987 => x"27",
          1988 => x"91",
          1989 => x"55",
          1990 => x"08",
          1991 => x"db",
          1992 => x"c8",
          1993 => x"19",
          1994 => x"c8",
          1995 => x"cb",
          1996 => x"80",
          1997 => x"08",
          1998 => x"bf",
          1999 => x"77",
          2000 => x"81",
          2001 => x"38",
          2002 => x"98",
          2003 => x"26",
          2004 => x"57",
          2005 => x"51",
          2006 => x"91",
          2007 => x"56",
          2008 => x"d3",
          2009 => x"2e",
          2010 => x"86",
          2011 => x"c8",
          2012 => x"ff",
          2013 => x"70",
          2014 => x"25",
          2015 => x"79",
          2016 => x"56",
          2017 => x"f3",
          2018 => x"2e",
          2019 => x"19",
          2020 => x"76",
          2021 => x"75",
          2022 => x"27",
          2023 => x"58",
          2024 => x"80",
          2025 => x"57",
          2026 => x"98",
          2027 => x"26",
          2028 => x"57",
          2029 => x"81",
          2030 => x"52",
          2031 => x"a9",
          2032 => x"c8",
          2033 => x"d3",
          2034 => x"2e",
          2035 => x"5a",
          2036 => x"08",
          2037 => x"81",
          2038 => x"91",
          2039 => x"5a",
          2040 => x"70",
          2041 => x"07",
          2042 => x"7d",
          2043 => x"56",
          2044 => x"ff",
          2045 => x"2e",
          2046 => x"ff",
          2047 => x"55",
          2048 => x"ff",
          2049 => x"78",
          2050 => x"3f",
          2051 => x"08",
          2052 => x"08",
          2053 => x"d3",
          2054 => x"80",
          2055 => x"70",
          2056 => x"2a",
          2057 => x"57",
          2058 => x"74",
          2059 => x"38",
          2060 => x"52",
          2061 => x"ad",
          2062 => x"c8",
          2063 => x"a6",
          2064 => x"1a",
          2065 => x"08",
          2066 => x"90",
          2067 => x"26",
          2068 => x"19",
          2069 => x"90",
          2070 => x"19",
          2071 => x"54",
          2072 => x"34",
          2073 => x"57",
          2074 => x"8d",
          2075 => x"80",
          2076 => x"75",
          2077 => x"81",
          2078 => x"74",
          2079 => x"0c",
          2080 => x"04",
          2081 => x"7b",
          2082 => x"f3",
          2083 => x"55",
          2084 => x"08",
          2085 => x"7c",
          2086 => x"f6",
          2087 => x"d3",
          2088 => x"d3",
          2089 => x"19",
          2090 => x"80",
          2091 => x"b4",
          2092 => x"55",
          2093 => x"74",
          2094 => x"80",
          2095 => x"77",
          2096 => x"17",
          2097 => x"75",
          2098 => x"77",
          2099 => x"53",
          2100 => x"17",
          2101 => x"81",
          2102 => x"c8",
          2103 => x"df",
          2104 => x"8a",
          2105 => x"58",
          2106 => x"83",
          2107 => x"77",
          2108 => x"d3",
          2109 => x"3d",
          2110 => x"3d",
          2111 => x"71",
          2112 => x"57",
          2113 => x"0a",
          2114 => x"74",
          2115 => x"72",
          2116 => x"38",
          2117 => x"ae",
          2118 => x"18",
          2119 => x"08",
          2120 => x"38",
          2121 => x"82",
          2122 => x"38",
          2123 => x"54",
          2124 => x"74",
          2125 => x"82",
          2126 => x"22",
          2127 => x"79",
          2128 => x"38",
          2129 => x"98",
          2130 => x"d1",
          2131 => x"22",
          2132 => x"54",
          2133 => x"26",
          2134 => x"52",
          2135 => x"89",
          2136 => x"c8",
          2137 => x"d3",
          2138 => x"2e",
          2139 => x"0b",
          2140 => x"08",
          2141 => x"98",
          2142 => x"d3",
          2143 => x"86",
          2144 => x"80",
          2145 => x"73",
          2146 => x"73",
          2147 => x"73",
          2148 => x"f4",
          2149 => x"d3",
          2150 => x"18",
          2151 => x"18",
          2152 => x"98",
          2153 => x"2e",
          2154 => x"39",
          2155 => x"39",
          2156 => x"98",
          2157 => x"98",
          2158 => x"83",
          2159 => x"b4",
          2160 => x"0c",
          2161 => x"91",
          2162 => x"8a",
          2163 => x"f9",
          2164 => x"7b",
          2165 => x"13",
          2166 => x"59",
          2167 => x"f0",
          2168 => x"27",
          2169 => x"0b",
          2170 => x"84",
          2171 => x"08",
          2172 => x"da",
          2173 => x"ff",
          2174 => x"81",
          2175 => x"15",
          2176 => x"98",
          2177 => x"15",
          2178 => x"75",
          2179 => x"18",
          2180 => x"77",
          2181 => x"a6",
          2182 => x"16",
          2183 => x"81",
          2184 => x"17",
          2185 => x"77",
          2186 => x"51",
          2187 => x"8e",
          2188 => x"08",
          2189 => x"f3",
          2190 => x"d3",
          2191 => x"82",
          2192 => x"91",
          2193 => x"27",
          2194 => x"81",
          2195 => x"c8",
          2196 => x"80",
          2197 => x"17",
          2198 => x"c8",
          2199 => x"cc",
          2200 => x"38",
          2201 => x"0c",
          2202 => x"e2",
          2203 => x"08",
          2204 => x"f8",
          2205 => x"d3",
          2206 => x"87",
          2207 => x"c8",
          2208 => x"80",
          2209 => x"53",
          2210 => x"08",
          2211 => x"38",
          2212 => x"d3",
          2213 => x"2e",
          2214 => x"d3",
          2215 => x"76",
          2216 => x"3f",
          2217 => x"d3",
          2218 => x"38",
          2219 => x"0c",
          2220 => x"51",
          2221 => x"91",
          2222 => x"98",
          2223 => x"90",
          2224 => x"83",
          2225 => x"b4",
          2226 => x"0c",
          2227 => x"91",
          2228 => x"89",
          2229 => x"f8",
          2230 => x"7c",
          2231 => x"5a",
          2232 => x"75",
          2233 => x"3f",
          2234 => x"08",
          2235 => x"c8",
          2236 => x"38",
          2237 => x"08",
          2238 => x"08",
          2239 => x"ef",
          2240 => x"d3",
          2241 => x"91",
          2242 => x"80",
          2243 => x"d3",
          2244 => x"17",
          2245 => x"51",
          2246 => x"81",
          2247 => x"81",
          2248 => x"81",
          2249 => x"70",
          2250 => x"07",
          2251 => x"80",
          2252 => x"81",
          2253 => x"79",
          2254 => x"83",
          2255 => x"81",
          2256 => x"fd",
          2257 => x"d3",
          2258 => x"91",
          2259 => x"80",
          2260 => x"38",
          2261 => x"09",
          2262 => x"38",
          2263 => x"91",
          2264 => x"8a",
          2265 => x"fd",
          2266 => x"9a",
          2267 => x"eb",
          2268 => x"d3",
          2269 => x"ff",
          2270 => x"70",
          2271 => x"53",
          2272 => x"09",
          2273 => x"38",
          2274 => x"eb",
          2275 => x"d3",
          2276 => x"2b",
          2277 => x"72",
          2278 => x"0c",
          2279 => x"04",
          2280 => x"77",
          2281 => x"ff",
          2282 => x"9a",
          2283 => x"55",
          2284 => x"76",
          2285 => x"53",
          2286 => x"09",
          2287 => x"38",
          2288 => x"52",
          2289 => x"eb",
          2290 => x"3d",
          2291 => x"3d",
          2292 => x"5b",
          2293 => x"08",
          2294 => x"16",
          2295 => x"81",
          2296 => x"16",
          2297 => x"51",
          2298 => x"91",
          2299 => x"58",
          2300 => x"08",
          2301 => x"9c",
          2302 => x"33",
          2303 => x"86",
          2304 => x"80",
          2305 => x"16",
          2306 => x"33",
          2307 => x"70",
          2308 => x"5a",
          2309 => x"72",
          2310 => x"74",
          2311 => x"70",
          2312 => x"32",
          2313 => x"73",
          2314 => x"53",
          2315 => x"54",
          2316 => x"9b",
          2317 => x"2e",
          2318 => x"77",
          2319 => x"54",
          2320 => x"09",
          2321 => x"38",
          2322 => x"7a",
          2323 => x"80",
          2324 => x"fa",
          2325 => x"d3",
          2326 => x"91",
          2327 => x"87",
          2328 => x"08",
          2329 => x"77",
          2330 => x"38",
          2331 => x"17",
          2332 => x"d3",
          2333 => x"3d",
          2334 => x"3d",
          2335 => x"08",
          2336 => x"52",
          2337 => x"f2",
          2338 => x"c8",
          2339 => x"d3",
          2340 => x"ef",
          2341 => x"84",
          2342 => x"39",
          2343 => x"52",
          2344 => x"a5",
          2345 => x"c8",
          2346 => x"d3",
          2347 => x"d1",
          2348 => x"08",
          2349 => x"54",
          2350 => x"db",
          2351 => x"08",
          2352 => x"bf",
          2353 => x"73",
          2354 => x"8b",
          2355 => x"83",
          2356 => x"06",
          2357 => x"73",
          2358 => x"53",
          2359 => x"74",
          2360 => x"3f",
          2361 => x"08",
          2362 => x"38",
          2363 => x"51",
          2364 => x"91",
          2365 => x"57",
          2366 => x"08",
          2367 => x"9c",
          2368 => x"73",
          2369 => x"0c",
          2370 => x"04",
          2371 => x"77",
          2372 => x"54",
          2373 => x"51",
          2374 => x"91",
          2375 => x"55",
          2376 => x"08",
          2377 => x"14",
          2378 => x"51",
          2379 => x"91",
          2380 => x"55",
          2381 => x"08",
          2382 => x"53",
          2383 => x"08",
          2384 => x"08",
          2385 => x"3f",
          2386 => x"14",
          2387 => x"08",
          2388 => x"3f",
          2389 => x"17",
          2390 => x"d3",
          2391 => x"3d",
          2392 => x"3d",
          2393 => x"08",
          2394 => x"54",
          2395 => x"53",
          2396 => x"91",
          2397 => x"54",
          2398 => x"08",
          2399 => x"13",
          2400 => x"73",
          2401 => x"83",
          2402 => x"91",
          2403 => x"86",
          2404 => x"fa",
          2405 => x"7a",
          2406 => x"0b",
          2407 => x"98",
          2408 => x"2e",
          2409 => x"80",
          2410 => x"9c",
          2411 => x"70",
          2412 => x"56",
          2413 => x"a0",
          2414 => x"72",
          2415 => x"81",
          2416 => x"81",
          2417 => x"89",
          2418 => x"06",
          2419 => x"15",
          2420 => x"ae",
          2421 => x"34",
          2422 => x"75",
          2423 => x"52",
          2424 => x"34",
          2425 => x"8a",
          2426 => x"38",
          2427 => x"05",
          2428 => x"81",
          2429 => x"17",
          2430 => x"12",
          2431 => x"34",
          2432 => x"9c",
          2433 => x"ac",
          2434 => x"c8",
          2435 => x"9c",
          2436 => x"05",
          2437 => x"3f",
          2438 => x"08",
          2439 => x"9c",
          2440 => x"05",
          2441 => x"3f",
          2442 => x"08",
          2443 => x"88",
          2444 => x"f5",
          2445 => x"70",
          2446 => x"05",
          2447 => x"8b",
          2448 => x"7a",
          2449 => x"3f",
          2450 => x"58",
          2451 => x"55",
          2452 => x"2e",
          2453 => x"80",
          2454 => x"17",
          2455 => x"19",
          2456 => x"70",
          2457 => x"2a",
          2458 => x"07",
          2459 => x"59",
          2460 => x"8c",
          2461 => x"54",
          2462 => x"81",
          2463 => x"39",
          2464 => x"70",
          2465 => x"dc",
          2466 => x"70",
          2467 => x"2a",
          2468 => x"51",
          2469 => x"2e",
          2470 => x"54",
          2471 => x"82",
          2472 => x"19",
          2473 => x"54",
          2474 => x"83",
          2475 => x"73",
          2476 => x"80",
          2477 => x"39",
          2478 => x"33",
          2479 => x"57",
          2480 => x"27",
          2481 => x"75",
          2482 => x"30",
          2483 => x"32",
          2484 => x"80",
          2485 => x"25",
          2486 => x"56",
          2487 => x"80",
          2488 => x"84",
          2489 => x"57",
          2490 => x"70",
          2491 => x"5a",
          2492 => x"09",
          2493 => x"38",
          2494 => x"77",
          2495 => x"51",
          2496 => x"80",
          2497 => x"81",
          2498 => x"81",
          2499 => x"07",
          2500 => x"38",
          2501 => x"75",
          2502 => x"30",
          2503 => x"7a",
          2504 => x"51",
          2505 => x"80",
          2506 => x"79",
          2507 => x"30",
          2508 => x"70",
          2509 => x"25",
          2510 => x"07",
          2511 => x"51",
          2512 => x"b1",
          2513 => x"8b",
          2514 => x"39",
          2515 => x"54",
          2516 => x"8c",
          2517 => x"ff",
          2518 => x"f8",
          2519 => x"54",
          2520 => x"e6",
          2521 => x"c8",
          2522 => x"b9",
          2523 => x"70",
          2524 => x"71",
          2525 => x"54",
          2526 => x"91",
          2527 => x"80",
          2528 => x"ff",
          2529 => x"78",
          2530 => x"86",
          2531 => x"39",
          2532 => x"75",
          2533 => x"18",
          2534 => x"58",
          2535 => x"81",
          2536 => x"94",
          2537 => x"91",
          2538 => x"e4",
          2539 => x"d3",
          2540 => x"c5",
          2541 => x"16",
          2542 => x"26",
          2543 => x"16",
          2544 => x"06",
          2545 => x"18",
          2546 => x"34",
          2547 => x"fd",
          2548 => x"19",
          2549 => x"54",
          2550 => x"a9",
          2551 => x"54",
          2552 => x"2e",
          2553 => x"84",
          2554 => x"34",
          2555 => x"76",
          2556 => x"89",
          2557 => x"8d",
          2558 => x"89",
          2559 => x"73",
          2560 => x"80",
          2561 => x"d3",
          2562 => x"3d",
          2563 => x"3d",
          2564 => x"08",
          2565 => x"7a",
          2566 => x"54",
          2567 => x"2e",
          2568 => x"55",
          2569 => x"33",
          2570 => x"72",
          2571 => x"83",
          2572 => x"74",
          2573 => x"72",
          2574 => x"38",
          2575 => x"88",
          2576 => x"39",
          2577 => x"80",
          2578 => x"51",
          2579 => x"af",
          2580 => x"06",
          2581 => x"55",
          2582 => x"33",
          2583 => x"72",
          2584 => x"09",
          2585 => x"38",
          2586 => x"74",
          2587 => x"d4",
          2588 => x"88",
          2589 => x"70",
          2590 => x"72",
          2591 => x"38",
          2592 => x"ab",
          2593 => x"52",
          2594 => x"ee",
          2595 => x"c8",
          2596 => x"aa",
          2597 => x"81",
          2598 => x"3d",
          2599 => x"75",
          2600 => x"3f",
          2601 => x"08",
          2602 => x"c8",
          2603 => x"38",
          2604 => x"c6",
          2605 => x"c8",
          2606 => x"33",
          2607 => x"d3",
          2608 => x"2e",
          2609 => x"91",
          2610 => x"84",
          2611 => x"06",
          2612 => x"73",
          2613 => x"81",
          2614 => x"72",
          2615 => x"38",
          2616 => x"70",
          2617 => x"53",
          2618 => x"ff",
          2619 => x"80",
          2620 => x"34",
          2621 => x"c6",
          2622 => x"2a",
          2623 => x"51",
          2624 => x"38",
          2625 => x"39",
          2626 => x"70",
          2627 => x"53",
          2628 => x"86",
          2629 => x"84",
          2630 => x"06",
          2631 => x"72",
          2632 => x"f1",
          2633 => x"08",
          2634 => x"17",
          2635 => x"76",
          2636 => x"3f",
          2637 => x"08",
          2638 => x"fe",
          2639 => x"91",
          2640 => x"88",
          2641 => x"f6",
          2642 => x"59",
          2643 => x"70",
          2644 => x"56",
          2645 => x"2e",
          2646 => x"76",
          2647 => x"58",
          2648 => x"32",
          2649 => x"a0",
          2650 => x"2a",
          2651 => x"52",
          2652 => x"38",
          2653 => x"09",
          2654 => x"a9",
          2655 => x"d0",
          2656 => x"70",
          2657 => x"38",
          2658 => x"81",
          2659 => x"11",
          2660 => x"70",
          2661 => x"ff",
          2662 => x"91",
          2663 => x"58",
          2664 => x"1b",
          2665 => x"08",
          2666 => x"75",
          2667 => x"57",
          2668 => x"81",
          2669 => x"ff",
          2670 => x"54",
          2671 => x"26",
          2672 => x"14",
          2673 => x"06",
          2674 => x"9f",
          2675 => x"99",
          2676 => x"e0",
          2677 => x"ff",
          2678 => x"73",
          2679 => x"32",
          2680 => x"72",
          2681 => x"73",
          2682 => x"53",
          2683 => x"70",
          2684 => x"73",
          2685 => x"32",
          2686 => x"72",
          2687 => x"73",
          2688 => x"53",
          2689 => x"70",
          2690 => x"38",
          2691 => x"83",
          2692 => x"8c",
          2693 => x"77",
          2694 => x"38",
          2695 => x"0c",
          2696 => x"86",
          2697 => x"f8",
          2698 => x"91",
          2699 => x"8c",
          2700 => x"fb",
          2701 => x"56",
          2702 => x"17",
          2703 => x"b0",
          2704 => x"52",
          2705 => x"81",
          2706 => x"91",
          2707 => x"81",
          2708 => x"b2",
          2709 => x"c3",
          2710 => x"c8",
          2711 => x"ff",
          2712 => x"55",
          2713 => x"d5",
          2714 => x"06",
          2715 => x"80",
          2716 => x"33",
          2717 => x"81",
          2718 => x"81",
          2719 => x"81",
          2720 => x"eb",
          2721 => x"70",
          2722 => x"07",
          2723 => x"73",
          2724 => x"16",
          2725 => x"81",
          2726 => x"81",
          2727 => x"83",
          2728 => x"80",
          2729 => x"16",
          2730 => x"3f",
          2731 => x"08",
          2732 => x"c8",
          2733 => x"9d",
          2734 => x"91",
          2735 => x"81",
          2736 => x"de",
          2737 => x"d3",
          2738 => x"91",
          2739 => x"80",
          2740 => x"82",
          2741 => x"d3",
          2742 => x"3d",
          2743 => x"3d",
          2744 => x"84",
          2745 => x"05",
          2746 => x"80",
          2747 => x"51",
          2748 => x"91",
          2749 => x"58",
          2750 => x"0b",
          2751 => x"08",
          2752 => x"38",
          2753 => x"08",
          2754 => x"d3",
          2755 => x"08",
          2756 => x"56",
          2757 => x"87",
          2758 => x"74",
          2759 => x"fe",
          2760 => x"54",
          2761 => x"2e",
          2762 => x"15",
          2763 => x"a6",
          2764 => x"c8",
          2765 => x"06",
          2766 => x"54",
          2767 => x"38",
          2768 => x"8f",
          2769 => x"2a",
          2770 => x"51",
          2771 => x"72",
          2772 => x"80",
          2773 => x"39",
          2774 => x"77",
          2775 => x"81",
          2776 => x"33",
          2777 => x"3f",
          2778 => x"08",
          2779 => x"70",
          2780 => x"54",
          2781 => x"86",
          2782 => x"80",
          2783 => x"73",
          2784 => x"81",
          2785 => x"8a",
          2786 => x"95",
          2787 => x"53",
          2788 => x"fd",
          2789 => x"d3",
          2790 => x"ff",
          2791 => x"82",
          2792 => x"06",
          2793 => x"79",
          2794 => x"29",
          2795 => x"75",
          2796 => x"f0",
          2797 => x"12",
          2798 => x"56",
          2799 => x"77",
          2800 => x"83",
          2801 => x"da",
          2802 => x"d3",
          2803 => x"76",
          2804 => x"14",
          2805 => x"27",
          2806 => x"54",
          2807 => x"10",
          2808 => x"11",
          2809 => x"83",
          2810 => x"2e",
          2811 => x"52",
          2812 => x"bf",
          2813 => x"c8",
          2814 => x"06",
          2815 => x"27",
          2816 => x"14",
          2817 => x"27",
          2818 => x"56",
          2819 => x"85",
          2820 => x"56",
          2821 => x"85",
          2822 => x"15",
          2823 => x"3f",
          2824 => x"08",
          2825 => x"06",
          2826 => x"72",
          2827 => x"09",
          2828 => x"ed",
          2829 => x"15",
          2830 => x"3f",
          2831 => x"08",
          2832 => x"06",
          2833 => x"38",
          2834 => x"51",
          2835 => x"91",
          2836 => x"54",
          2837 => x"0c",
          2838 => x"33",
          2839 => x"80",
          2840 => x"ff",
          2841 => x"56",
          2842 => x"84",
          2843 => x"15",
          2844 => x"29",
          2845 => x"33",
          2846 => x"72",
          2847 => x"72",
          2848 => x"06",
          2849 => x"2e",
          2850 => x"13",
          2851 => x"72",
          2852 => x"38",
          2853 => x"89",
          2854 => x"15",
          2855 => x"3f",
          2856 => x"08",
          2857 => x"91",
          2858 => x"83",
          2859 => x"8f",
          2860 => x"56",
          2861 => x"38",
          2862 => x"51",
          2863 => x"91",
          2864 => x"83",
          2865 => x"53",
          2866 => x"80",
          2867 => x"d8",
          2868 => x"d3",
          2869 => x"80",
          2870 => x"d8",
          2871 => x"d3",
          2872 => x"ff",
          2873 => x"8d",
          2874 => x"2e",
          2875 => x"88",
          2876 => x"1a",
          2877 => x"05",
          2878 => x"56",
          2879 => x"83",
          2880 => x"15",
          2881 => x"78",
          2882 => x"b0",
          2883 => x"d3",
          2884 => x"8d",
          2885 => x"c8",
          2886 => x"83",
          2887 => x"57",
          2888 => x"08",
          2889 => x"ff",
          2890 => x"38",
          2891 => x"83",
          2892 => x"83",
          2893 => x"72",
          2894 => x"83",
          2895 => x"8d",
          2896 => x"2e",
          2897 => x"82",
          2898 => x"0c",
          2899 => x"0c",
          2900 => x"16",
          2901 => x"ac",
          2902 => x"83",
          2903 => x"06",
          2904 => x"de",
          2905 => x"b3",
          2906 => x"c8",
          2907 => x"ff",
          2908 => x"56",
          2909 => x"38",
          2910 => x"53",
          2911 => x"82",
          2912 => x"e0",
          2913 => x"ac",
          2914 => x"c8",
          2915 => x"0c",
          2916 => x"82",
          2917 => x"39",
          2918 => x"53",
          2919 => x"80",
          2920 => x"38",
          2921 => x"14",
          2922 => x"76",
          2923 => x"81",
          2924 => x"98",
          2925 => x"53",
          2926 => x"15",
          2927 => x"16",
          2928 => x"81",
          2929 => x"08",
          2930 => x"51",
          2931 => x"13",
          2932 => x"8d",
          2933 => x"16",
          2934 => x"c5",
          2935 => x"90",
          2936 => x"0b",
          2937 => x"ff",
          2938 => x"16",
          2939 => x"2e",
          2940 => x"81",
          2941 => x"e4",
          2942 => x"9f",
          2943 => x"c8",
          2944 => x"ff",
          2945 => x"81",
          2946 => x"06",
          2947 => x"81",
          2948 => x"51",
          2949 => x"91",
          2950 => x"80",
          2951 => x"d3",
          2952 => x"16",
          2953 => x"15",
          2954 => x"3f",
          2955 => x"08",
          2956 => x"06",
          2957 => x"d4",
          2958 => x"81",
          2959 => x"38",
          2960 => x"d5",
          2961 => x"d3",
          2962 => x"8b",
          2963 => x"2e",
          2964 => x"b3",
          2965 => x"15",
          2966 => x"3f",
          2967 => x"08",
          2968 => x"e4",
          2969 => x"81",
          2970 => x"84",
          2971 => x"d5",
          2972 => x"d3",
          2973 => x"16",
          2974 => x"15",
          2975 => x"3f",
          2976 => x"08",
          2977 => x"76",
          2978 => x"d3",
          2979 => x"05",
          2980 => x"d3",
          2981 => x"86",
          2982 => x"0b",
          2983 => x"80",
          2984 => x"d3",
          2985 => x"3d",
          2986 => x"3d",
          2987 => x"89",
          2988 => x"2e",
          2989 => x"08",
          2990 => x"38",
          2991 => x"33",
          2992 => x"80",
          2993 => x"84",
          2994 => x"14",
          2995 => x"71",
          2996 => x"81",
          2997 => x"81",
          2998 => x"ce",
          2999 => x"d3",
          3000 => x"06",
          3001 => x"38",
          3002 => x"53",
          3003 => x"09",
          3004 => x"38",
          3005 => x"78",
          3006 => x"52",
          3007 => x"c8",
          3008 => x"0d",
          3009 => x"0d",
          3010 => x"33",
          3011 => x"3d",
          3012 => x"56",
          3013 => x"91",
          3014 => x"55",
          3015 => x"0b",
          3016 => x"08",
          3017 => x"38",
          3018 => x"08",
          3019 => x"d3",
          3020 => x"08",
          3021 => x"80",
          3022 => x"80",
          3023 => x"80",
          3024 => x"78",
          3025 => x"34",
          3026 => x"91",
          3027 => x"79",
          3028 => x"75",
          3029 => x"2e",
          3030 => x"53",
          3031 => x"53",
          3032 => x"f6",
          3033 => x"d3",
          3034 => x"73",
          3035 => x"0c",
          3036 => x"04",
          3037 => x"67",
          3038 => x"80",
          3039 => x"58",
          3040 => x"77",
          3041 => x"e9",
          3042 => x"06",
          3043 => x"3d",
          3044 => x"99",
          3045 => x"52",
          3046 => x"3f",
          3047 => x"08",
          3048 => x"c8",
          3049 => x"38",
          3050 => x"52",
          3051 => x"05",
          3052 => x"3f",
          3053 => x"08",
          3054 => x"c8",
          3055 => x"02",
          3056 => x"33",
          3057 => x"56",
          3058 => x"25",
          3059 => x"56",
          3060 => x"55",
          3061 => x"81",
          3062 => x"80",
          3063 => x"75",
          3064 => x"81",
          3065 => x"97",
          3066 => x"51",
          3067 => x"91",
          3068 => x"56",
          3069 => x"57",
          3070 => x"b2",
          3071 => x"06",
          3072 => x"2e",
          3073 => x"56",
          3074 => x"82",
          3075 => x"06",
          3076 => x"80",
          3077 => x"88",
          3078 => x"d0",
          3079 => x"2a",
          3080 => x"51",
          3081 => x"2e",
          3082 => x"62",
          3083 => x"e6",
          3084 => x"d3",
          3085 => x"82",
          3086 => x"52",
          3087 => x"51",
          3088 => x"62",
          3089 => x"8b",
          3090 => x"53",
          3091 => x"51",
          3092 => x"75",
          3093 => x"05",
          3094 => x"3f",
          3095 => x"0b",
          3096 => x"78",
          3097 => x"e9",
          3098 => x"11",
          3099 => x"7a",
          3100 => x"d4",
          3101 => x"55",
          3102 => x"91",
          3103 => x"56",
          3104 => x"08",
          3105 => x"74",
          3106 => x"d4",
          3107 => x"d3",
          3108 => x"ff",
          3109 => x"0c",
          3110 => x"39",
          3111 => x"38",
          3112 => x"33",
          3113 => x"70",
          3114 => x"56",
          3115 => x"2e",
          3116 => x"56",
          3117 => x"81",
          3118 => x"06",
          3119 => x"80",
          3120 => x"02",
          3121 => x"81",
          3122 => x"80",
          3123 => x"87",
          3124 => x"98",
          3125 => x"2a",
          3126 => x"51",
          3127 => x"2e",
          3128 => x"80",
          3129 => x"7a",
          3130 => x"a0",
          3131 => x"a4",
          3132 => x"75",
          3133 => x"62",
          3134 => x"e4",
          3135 => x"d3",
          3136 => x"19",
          3137 => x"05",
          3138 => x"3f",
          3139 => x"08",
          3140 => x"74",
          3141 => x"15",
          3142 => x"23",
          3143 => x"34",
          3144 => x"34",
          3145 => x"0c",
          3146 => x"0c",
          3147 => x"75",
          3148 => x"51",
          3149 => x"76",
          3150 => x"81",
          3151 => x"74",
          3152 => x"a3",
          3153 => x"08",
          3154 => x"9b",
          3155 => x"08",
          3156 => x"7a",
          3157 => x"70",
          3158 => x"1b",
          3159 => x"08",
          3160 => x"51",
          3161 => x"76",
          3162 => x"d4",
          3163 => x"d3",
          3164 => x"91",
          3165 => x"81",
          3166 => x"82",
          3167 => x"2e",
          3168 => x"83",
          3169 => x"78",
          3170 => x"75",
          3171 => x"07",
          3172 => x"7b",
          3173 => x"51",
          3174 => x"cb",
          3175 => x"19",
          3176 => x"c8",
          3177 => x"ff",
          3178 => x"80",
          3179 => x"76",
          3180 => x"d4",
          3181 => x"d3",
          3182 => x"38",
          3183 => x"39",
          3184 => x"91",
          3185 => x"05",
          3186 => x"0c",
          3187 => x"74",
          3188 => x"52",
          3189 => x"33",
          3190 => x"a4",
          3191 => x"c8",
          3192 => x"83",
          3193 => x"75",
          3194 => x"38",
          3195 => x"75",
          3196 => x"d3",
          3197 => x"3d",
          3198 => x"3d",
          3199 => x"64",
          3200 => x"5a",
          3201 => x"0c",
          3202 => x"05",
          3203 => x"f9",
          3204 => x"d3",
          3205 => x"91",
          3206 => x"8a",
          3207 => x"33",
          3208 => x"2e",
          3209 => x"56",
          3210 => x"90",
          3211 => x"06",
          3212 => x"74",
          3213 => x"a0",
          3214 => x"82",
          3215 => x"34",
          3216 => x"94",
          3217 => x"91",
          3218 => x"56",
          3219 => x"82",
          3220 => x"34",
          3221 => x"80",
          3222 => x"91",
          3223 => x"56",
          3224 => x"81",
          3225 => x"34",
          3226 => x"ec",
          3227 => x"91",
          3228 => x"56",
          3229 => x"8c",
          3230 => x"18",
          3231 => x"74",
          3232 => x"38",
          3233 => x"80",
          3234 => x"38",
          3235 => x"70",
          3236 => x"56",
          3237 => x"83",
          3238 => x"11",
          3239 => x"77",
          3240 => x"5c",
          3241 => x"38",
          3242 => x"88",
          3243 => x"8f",
          3244 => x"08",
          3245 => x"d2",
          3246 => x"d3",
          3247 => x"81",
          3248 => x"f7",
          3249 => x"2e",
          3250 => x"74",
          3251 => x"98",
          3252 => x"7d",
          3253 => x"3f",
          3254 => x"08",
          3255 => x"ef",
          3256 => x"c8",
          3257 => x"89",
          3258 => x"79",
          3259 => x"d7",
          3260 => x"7e",
          3261 => x"51",
          3262 => x"76",
          3263 => x"74",
          3264 => x"79",
          3265 => x"7b",
          3266 => x"11",
          3267 => x"c7",
          3268 => x"d3",
          3269 => x"c1",
          3270 => x"33",
          3271 => x"56",
          3272 => x"25",
          3273 => x"17",
          3274 => x"55",
          3275 => x"90",
          3276 => x"53",
          3277 => x"74",
          3278 => x"1c",
          3279 => x"3f",
          3280 => x"56",
          3281 => x"9c",
          3282 => x"2e",
          3283 => x"90",
          3284 => x"98",
          3285 => x"74",
          3286 => x"38",
          3287 => x"17",
          3288 => x"17",
          3289 => x"11",
          3290 => x"c8",
          3291 => x"d3",
          3292 => x"ef",
          3293 => x"33",
          3294 => x"55",
          3295 => x"34",
          3296 => x"53",
          3297 => x"7d",
          3298 => x"52",
          3299 => x"3f",
          3300 => x"08",
          3301 => x"77",
          3302 => x"94",
          3303 => x"ff",
          3304 => x"71",
          3305 => x"78",
          3306 => x"38",
          3307 => x"53",
          3308 => x"83",
          3309 => x"a8",
          3310 => x"51",
          3311 => x"78",
          3312 => x"08",
          3313 => x"76",
          3314 => x"08",
          3315 => x"0c",
          3316 => x"fd",
          3317 => x"56",
          3318 => x"c8",
          3319 => x"0d",
          3320 => x"0d",
          3321 => x"63",
          3322 => x"57",
          3323 => x"8f",
          3324 => x"52",
          3325 => x"b2",
          3326 => x"c8",
          3327 => x"d3",
          3328 => x"38",
          3329 => x"55",
          3330 => x"86",
          3331 => x"84",
          3332 => x"17",
          3333 => x"2a",
          3334 => x"51",
          3335 => x"56",
          3336 => x"83",
          3337 => x"39",
          3338 => x"18",
          3339 => x"83",
          3340 => x"0b",
          3341 => x"81",
          3342 => x"39",
          3343 => x"18",
          3344 => x"83",
          3345 => x"0b",
          3346 => x"82",
          3347 => x"39",
          3348 => x"18",
          3349 => x"83",
          3350 => x"0b",
          3351 => x"81",
          3352 => x"39",
          3353 => x"19",
          3354 => x"18",
          3355 => x"38",
          3356 => x"09",
          3357 => x"2e",
          3358 => x"94",
          3359 => x"83",
          3360 => x"56",
          3361 => x"38",
          3362 => x"22",
          3363 => x"89",
          3364 => x"55",
          3365 => x"38",
          3366 => x"88",
          3367 => x"74",
          3368 => x"52",
          3369 => x"b8",
          3370 => x"c8",
          3371 => x"39",
          3372 => x"52",
          3373 => x"a8",
          3374 => x"c8",
          3375 => x"80",
          3376 => x"38",
          3377 => x"fe",
          3378 => x"ff",
          3379 => x"38",
          3380 => x"0c",
          3381 => x"85",
          3382 => x"18",
          3383 => x"33",
          3384 => x"56",
          3385 => x"25",
          3386 => x"54",
          3387 => x"53",
          3388 => x"7d",
          3389 => x"52",
          3390 => x"3f",
          3391 => x"08",
          3392 => x"90",
          3393 => x"ff",
          3394 => x"90",
          3395 => x"17",
          3396 => x"51",
          3397 => x"91",
          3398 => x"80",
          3399 => x"38",
          3400 => x"08",
          3401 => x"2a",
          3402 => x"80",
          3403 => x"38",
          3404 => x"8a",
          3405 => x"56",
          3406 => x"27",
          3407 => x"7b",
          3408 => x"54",
          3409 => x"52",
          3410 => x"33",
          3411 => x"89",
          3412 => x"c8",
          3413 => x"38",
          3414 => x"78",
          3415 => x"7a",
          3416 => x"84",
          3417 => x"84",
          3418 => x"52",
          3419 => x"c8",
          3420 => x"17",
          3421 => x"06",
          3422 => x"18",
          3423 => x"2b",
          3424 => x"39",
          3425 => x"78",
          3426 => x"94",
          3427 => x"18",
          3428 => x"38",
          3429 => x"53",
          3430 => x"7d",
          3431 => x"52",
          3432 => x"3f",
          3433 => x"08",
          3434 => x"77",
          3435 => x"94",
          3436 => x"ff",
          3437 => x"71",
          3438 => x"78",
          3439 => x"38",
          3440 => x"53",
          3441 => x"17",
          3442 => x"06",
          3443 => x"51",
          3444 => x"90",
          3445 => x"80",
          3446 => x"90",
          3447 => x"76",
          3448 => x"17",
          3449 => x"1d",
          3450 => x"18",
          3451 => x"0c",
          3452 => x"58",
          3453 => x"74",
          3454 => x"38",
          3455 => x"8c",
          3456 => x"fc",
          3457 => x"17",
          3458 => x"07",
          3459 => x"18",
          3460 => x"75",
          3461 => x"0c",
          3462 => x"04",
          3463 => x"7b",
          3464 => x"05",
          3465 => x"58",
          3466 => x"91",
          3467 => x"57",
          3468 => x"08",
          3469 => x"90",
          3470 => x"86",
          3471 => x"06",
          3472 => x"74",
          3473 => x"98",
          3474 => x"2b",
          3475 => x"25",
          3476 => x"54",
          3477 => x"53",
          3478 => x"79",
          3479 => x"52",
          3480 => x"3f",
          3481 => x"d3",
          3482 => x"f6",
          3483 => x"33",
          3484 => x"55",
          3485 => x"34",
          3486 => x"52",
          3487 => x"c9",
          3488 => x"c8",
          3489 => x"d3",
          3490 => x"d4",
          3491 => x"08",
          3492 => x"a0",
          3493 => x"74",
          3494 => x"88",
          3495 => x"75",
          3496 => x"51",
          3497 => x"8c",
          3498 => x"9c",
          3499 => x"cb",
          3500 => x"b2",
          3501 => x"16",
          3502 => x"3f",
          3503 => x"16",
          3504 => x"3f",
          3505 => x"0b",
          3506 => x"79",
          3507 => x"3f",
          3508 => x"08",
          3509 => x"81",
          3510 => x"57",
          3511 => x"34",
          3512 => x"91",
          3513 => x"8b",
          3514 => x"fc",
          3515 => x"70",
          3516 => x"a8",
          3517 => x"c8",
          3518 => x"d3",
          3519 => x"38",
          3520 => x"05",
          3521 => x"ef",
          3522 => x"d3",
          3523 => x"91",
          3524 => x"87",
          3525 => x"c8",
          3526 => x"72",
          3527 => x"0c",
          3528 => x"04",
          3529 => x"85",
          3530 => x"9b",
          3531 => x"80",
          3532 => x"c8",
          3533 => x"38",
          3534 => x"08",
          3535 => x"34",
          3536 => x"91",
          3537 => x"84",
          3538 => x"ef",
          3539 => x"53",
          3540 => x"05",
          3541 => x"51",
          3542 => x"91",
          3543 => x"55",
          3544 => x"08",
          3545 => x"76",
          3546 => x"93",
          3547 => x"51",
          3548 => x"91",
          3549 => x"55",
          3550 => x"08",
          3551 => x"80",
          3552 => x"70",
          3553 => x"56",
          3554 => x"89",
          3555 => x"94",
          3556 => x"a7",
          3557 => x"05",
          3558 => x"2a",
          3559 => x"51",
          3560 => x"80",
          3561 => x"76",
          3562 => x"52",
          3563 => x"3f",
          3564 => x"08",
          3565 => x"83",
          3566 => x"74",
          3567 => x"81",
          3568 => x"85",
          3569 => x"d3",
          3570 => x"3d",
          3571 => x"3d",
          3572 => x"08",
          3573 => x"5b",
          3574 => x"34",
          3575 => x"3d",
          3576 => x"52",
          3577 => x"e5",
          3578 => x"d3",
          3579 => x"91",
          3580 => x"83",
          3581 => x"46",
          3582 => x"11",
          3583 => x"68",
          3584 => x"80",
          3585 => x"38",
          3586 => x"94",
          3587 => x"5b",
          3588 => x"51",
          3589 => x"91",
          3590 => x"57",
          3591 => x"08",
          3592 => x"6b",
          3593 => x"c5",
          3594 => x"d3",
          3595 => x"91",
          3596 => x"81",
          3597 => x"52",
          3598 => x"ab",
          3599 => x"c8",
          3600 => x"52",
          3601 => x"b2",
          3602 => x"c8",
          3603 => x"d3",
          3604 => x"ac",
          3605 => x"80",
          3606 => x"d6",
          3607 => x"d3",
          3608 => x"91",
          3609 => x"a4",
          3610 => x"7e",
          3611 => x"3f",
          3612 => x"08",
          3613 => x"38",
          3614 => x"51",
          3615 => x"91",
          3616 => x"57",
          3617 => x"08",
          3618 => x"38",
          3619 => x"09",
          3620 => x"38",
          3621 => x"81",
          3622 => x"3d",
          3623 => x"53",
          3624 => x"d9",
          3625 => x"93",
          3626 => x"12",
          3627 => x"51",
          3628 => x"56",
          3629 => x"8e",
          3630 => x"70",
          3631 => x"33",
          3632 => x"73",
          3633 => x"16",
          3634 => x"27",
          3635 => x"57",
          3636 => x"80",
          3637 => x"7d",
          3638 => x"a3",
          3639 => x"ff",
          3640 => x"57",
          3641 => x"81",
          3642 => x"34",
          3643 => x"ff",
          3644 => x"08",
          3645 => x"af",
          3646 => x"55",
          3647 => x"38",
          3648 => x"38",
          3649 => x"09",
          3650 => x"38",
          3651 => x"3d",
          3652 => x"59",
          3653 => x"80",
          3654 => x"f8",
          3655 => x"10",
          3656 => x"05",
          3657 => x"33",
          3658 => x"57",
          3659 => x"78",
          3660 => x"81",
          3661 => x"70",
          3662 => x"56",
          3663 => x"82",
          3664 => x"79",
          3665 => x"80",
          3666 => x"27",
          3667 => x"15",
          3668 => x"7a",
          3669 => x"5c",
          3670 => x"58",
          3671 => x"ee",
          3672 => x"70",
          3673 => x"34",
          3674 => x"77",
          3675 => x"57",
          3676 => x"a2",
          3677 => x"81",
          3678 => x"73",
          3679 => x"81",
          3680 => x"7b",
          3681 => x"38",
          3682 => x"76",
          3683 => x"0c",
          3684 => x"04",
          3685 => x"7e",
          3686 => x"fc",
          3687 => x"53",
          3688 => x"86",
          3689 => x"c8",
          3690 => x"d3",
          3691 => x"38",
          3692 => x"5a",
          3693 => x"86",
          3694 => x"83",
          3695 => x"17",
          3696 => x"94",
          3697 => x"33",
          3698 => x"70",
          3699 => x"56",
          3700 => x"38",
          3701 => x"58",
          3702 => x"56",
          3703 => x"19",
          3704 => x"7b",
          3705 => x"38",
          3706 => x"22",
          3707 => x"5b",
          3708 => x"7b",
          3709 => x"78",
          3710 => x"51",
          3711 => x"3f",
          3712 => x"08",
          3713 => x"54",
          3714 => x"55",
          3715 => x"3f",
          3716 => x"08",
          3717 => x"38",
          3718 => x"06",
          3719 => x"77",
          3720 => x"31",
          3721 => x"57",
          3722 => x"39",
          3723 => x"56",
          3724 => x"75",
          3725 => x"c9",
          3726 => x"d3",
          3727 => x"91",
          3728 => x"81",
          3729 => x"06",
          3730 => x"0b",
          3731 => x"82",
          3732 => x"39",
          3733 => x"08",
          3734 => x"81",
          3735 => x"81",
          3736 => x"34",
          3737 => x"ce",
          3738 => x"c8",
          3739 => x"0c",
          3740 => x"0c",
          3741 => x"81",
          3742 => x"78",
          3743 => x"38",
          3744 => x"94",
          3745 => x"94",
          3746 => x"18",
          3747 => x"2a",
          3748 => x"51",
          3749 => x"74",
          3750 => x"38",
          3751 => x"51",
          3752 => x"91",
          3753 => x"56",
          3754 => x"08",
          3755 => x"d3",
          3756 => x"b5",
          3757 => x"76",
          3758 => x"3f",
          3759 => x"08",
          3760 => x"2e",
          3761 => x"81",
          3762 => x"38",
          3763 => x"15",
          3764 => x"8b",
          3765 => x"91",
          3766 => x"55",
          3767 => x"75",
          3768 => x"77",
          3769 => x"98",
          3770 => x"08",
          3771 => x"0c",
          3772 => x"06",
          3773 => x"2e",
          3774 => x"52",
          3775 => x"bf",
          3776 => x"c8",
          3777 => x"82",
          3778 => x"34",
          3779 => x"a6",
          3780 => x"2a",
          3781 => x"08",
          3782 => x"17",
          3783 => x"08",
          3784 => x"94",
          3785 => x"18",
          3786 => x"33",
          3787 => x"55",
          3788 => x"34",
          3789 => x"83",
          3790 => x"74",
          3791 => x"f4",
          3792 => x"08",
          3793 => x"ec",
          3794 => x"33",
          3795 => x"56",
          3796 => x"25",
          3797 => x"54",
          3798 => x"53",
          3799 => x"7c",
          3800 => x"52",
          3801 => x"f1",
          3802 => x"c8",
          3803 => x"8a",
          3804 => x"91",
          3805 => x"55",
          3806 => x"17",
          3807 => x"06",
          3808 => x"18",
          3809 => x"7a",
          3810 => x"52",
          3811 => x"33",
          3812 => x"b6",
          3813 => x"d3",
          3814 => x"2e",
          3815 => x"0b",
          3816 => x"81",
          3817 => x"81",
          3818 => x"34",
          3819 => x"39",
          3820 => x"0c",
          3821 => x"91",
          3822 => x"8e",
          3823 => x"f9",
          3824 => x"56",
          3825 => x"80",
          3826 => x"38",
          3827 => x"3d",
          3828 => x"8a",
          3829 => x"51",
          3830 => x"91",
          3831 => x"55",
          3832 => x"08",
          3833 => x"77",
          3834 => x"52",
          3835 => x"9e",
          3836 => x"c8",
          3837 => x"d3",
          3838 => x"ca",
          3839 => x"33",
          3840 => x"55",
          3841 => x"24",
          3842 => x"16",
          3843 => x"2a",
          3844 => x"51",
          3845 => x"80",
          3846 => x"9c",
          3847 => x"77",
          3848 => x"3f",
          3849 => x"08",
          3850 => x"83",
          3851 => x"74",
          3852 => x"54",
          3853 => x"84",
          3854 => x"52",
          3855 => x"ba",
          3856 => x"c8",
          3857 => x"84",
          3858 => x"06",
          3859 => x"55",
          3860 => x"84",
          3861 => x"0c",
          3862 => x"91",
          3863 => x"89",
          3864 => x"fc",
          3865 => x"87",
          3866 => x"53",
          3867 => x"e4",
          3868 => x"d3",
          3869 => x"91",
          3870 => x"87",
          3871 => x"c8",
          3872 => x"72",
          3873 => x"0c",
          3874 => x"04",
          3875 => x"77",
          3876 => x"fc",
          3877 => x"53",
          3878 => x"8e",
          3879 => x"c8",
          3880 => x"d3",
          3881 => x"d1",
          3882 => x"38",
          3883 => x"08",
          3884 => x"c8",
          3885 => x"d3",
          3886 => x"bd",
          3887 => x"73",
          3888 => x"3f",
          3889 => x"08",
          3890 => x"c8",
          3891 => x"09",
          3892 => x"38",
          3893 => x"a1",
          3894 => x"73",
          3895 => x"3f",
          3896 => x"51",
          3897 => x"91",
          3898 => x"53",
          3899 => x"08",
          3900 => x"81",
          3901 => x"80",
          3902 => x"d3",
          3903 => x"3d",
          3904 => x"3d",
          3905 => x"80",
          3906 => x"70",
          3907 => x"52",
          3908 => x"3f",
          3909 => x"08",
          3910 => x"c8",
          3911 => x"63",
          3912 => x"d5",
          3913 => x"d3",
          3914 => x"91",
          3915 => x"a3",
          3916 => x"c7",
          3917 => x"98",
          3918 => x"73",
          3919 => x"38",
          3920 => x"39",
          3921 => x"8b",
          3922 => x"93",
          3923 => x"51",
          3924 => x"74",
          3925 => x"0c",
          3926 => x"04",
          3927 => x"61",
          3928 => x"80",
          3929 => x"ec",
          3930 => x"3d",
          3931 => x"3f",
          3932 => x"08",
          3933 => x"c8",
          3934 => x"38",
          3935 => x"73",
          3936 => x"08",
          3937 => x"55",
          3938 => x"74",
          3939 => x"90",
          3940 => x"0c",
          3941 => x"81",
          3942 => x"39",
          3943 => x"ca",
          3944 => x"70",
          3945 => x"57",
          3946 => x"09",
          3947 => x"c0",
          3948 => x"5d",
          3949 => x"90",
          3950 => x"51",
          3951 => x"3f",
          3952 => x"08",
          3953 => x"38",
          3954 => x"08",
          3955 => x"38",
          3956 => x"08",
          3957 => x"d3",
          3958 => x"80",
          3959 => x"81",
          3960 => x"58",
          3961 => x"14",
          3962 => x"c9",
          3963 => x"39",
          3964 => x"08",
          3965 => x"5a",
          3966 => x"55",
          3967 => x"77",
          3968 => x"7b",
          3969 => x"b9",
          3970 => x"d3",
          3971 => x"91",
          3972 => x"80",
          3973 => x"70",
          3974 => x"73",
          3975 => x"81",
          3976 => x"7a",
          3977 => x"51",
          3978 => x"3f",
          3979 => x"08",
          3980 => x"06",
          3981 => x"80",
          3982 => x"18",
          3983 => x"54",
          3984 => x"15",
          3985 => x"ff",
          3986 => x"91",
          3987 => x"f0",
          3988 => x"30",
          3989 => x"19",
          3990 => x"59",
          3991 => x"83",
          3992 => x"17",
          3993 => x"ff",
          3994 => x"7a",
          3995 => x"90",
          3996 => x"7a",
          3997 => x"81",
          3998 => x"73",
          3999 => x"78",
          4000 => x"0c",
          4001 => x"04",
          4002 => x"7a",
          4003 => x"05",
          4004 => x"58",
          4005 => x"91",
          4006 => x"57",
          4007 => x"08",
          4008 => x"18",
          4009 => x"80",
          4010 => x"76",
          4011 => x"39",
          4012 => x"70",
          4013 => x"81",
          4014 => x"56",
          4015 => x"80",
          4016 => x"38",
          4017 => x"8c",
          4018 => x"81",
          4019 => x"18",
          4020 => x"80",
          4021 => x"08",
          4022 => x"ff",
          4023 => x"91",
          4024 => x"57",
          4025 => x"19",
          4026 => x"39",
          4027 => x"52",
          4028 => x"b9",
          4029 => x"d3",
          4030 => x"d3",
          4031 => x"32",
          4032 => x"72",
          4033 => x"52",
          4034 => x"91",
          4035 => x"81",
          4036 => x"06",
          4037 => x"57",
          4038 => x"78",
          4039 => x"16",
          4040 => x"38",
          4041 => x"53",
          4042 => x"51",
          4043 => x"3f",
          4044 => x"08",
          4045 => x"08",
          4046 => x"90",
          4047 => x"c0",
          4048 => x"90",
          4049 => x"b9",
          4050 => x"2b",
          4051 => x"25",
          4052 => x"54",
          4053 => x"53",
          4054 => x"78",
          4055 => x"52",
          4056 => x"f5",
          4057 => x"c8",
          4058 => x"85",
          4059 => x"8c",
          4060 => x"33",
          4061 => x"55",
          4062 => x"34",
          4063 => x"89",
          4064 => x"19",
          4065 => x"83",
          4066 => x"75",
          4067 => x"0c",
          4068 => x"04",
          4069 => x"91",
          4070 => x"ff",
          4071 => x"82",
          4072 => x"ff",
          4073 => x"a0",
          4074 => x"b2",
          4075 => x"c8",
          4076 => x"d3",
          4077 => x"d3",
          4078 => x"90",
          4079 => x"b3",
          4080 => x"6f",
          4081 => x"d4",
          4082 => x"c2",
          4083 => x"c8",
          4084 => x"94",
          4085 => x"96",
          4086 => x"82",
          4087 => x"80",
          4088 => x"70",
          4089 => x"81",
          4090 => x"55",
          4091 => x"83",
          4092 => x"75",
          4093 => x"91",
          4094 => x"ff",
          4095 => x"02",
          4096 => x"33",
          4097 => x"55",
          4098 => x"25",
          4099 => x"56",
          4100 => x"80",
          4101 => x"81",
          4102 => x"80",
          4103 => x"87",
          4104 => x"e7",
          4105 => x"77",
          4106 => x"3f",
          4107 => x"08",
          4108 => x"80",
          4109 => x"70",
          4110 => x"81",
          4111 => x"56",
          4112 => x"2e",
          4113 => x"91",
          4114 => x"ff",
          4115 => x"87",
          4116 => x"94",
          4117 => x"2e",
          4118 => x"91",
          4119 => x"ff",
          4120 => x"77",
          4121 => x"91",
          4122 => x"ff",
          4123 => x"80",
          4124 => x"70",
          4125 => x"82",
          4126 => x"c8",
          4127 => x"d3",
          4128 => x"87",
          4129 => x"c8",
          4130 => x"51",
          4131 => x"91",
          4132 => x"56",
          4133 => x"08",
          4134 => x"56",
          4135 => x"70",
          4136 => x"07",
          4137 => x"06",
          4138 => x"75",
          4139 => x"91",
          4140 => x"ff",
          4141 => x"9f",
          4142 => x"51",
          4143 => x"91",
          4144 => x"91",
          4145 => x"30",
          4146 => x"c8",
          4147 => x"25",
          4148 => x"7b",
          4149 => x"72",
          4150 => x"51",
          4151 => x"80",
          4152 => x"91",
          4153 => x"ff",
          4154 => x"80",
          4155 => x"9f",
          4156 => x"51",
          4157 => x"3f",
          4158 => x"08",
          4159 => x"38",
          4160 => x"b4",
          4161 => x"d3",
          4162 => x"91",
          4163 => x"ff",
          4164 => x"75",
          4165 => x"0c",
          4166 => x"04",
          4167 => x"82",
          4168 => x"c0",
          4169 => x"3d",
          4170 => x"3f",
          4171 => x"08",
          4172 => x"c8",
          4173 => x"38",
          4174 => x"52",
          4175 => x"05",
          4176 => x"3f",
          4177 => x"08",
          4178 => x"c8",
          4179 => x"88",
          4180 => x"2e",
          4181 => x"82",
          4182 => x"80",
          4183 => x"70",
          4184 => x"81",
          4185 => x"56",
          4186 => x"83",
          4187 => x"74",
          4188 => x"81",
          4189 => x"38",
          4190 => x"52",
          4191 => x"05",
          4192 => x"dc",
          4193 => x"c8",
          4194 => x"55",
          4195 => x"08",
          4196 => x"81",
          4197 => x"87",
          4198 => x"2e",
          4199 => x"83",
          4200 => x"75",
          4201 => x"81",
          4202 => x"81",
          4203 => x"b2",
          4204 => x"81",
          4205 => x"52",
          4206 => x"bd",
          4207 => x"d3",
          4208 => x"91",
          4209 => x"81",
          4210 => x"53",
          4211 => x"18",
          4212 => x"fa",
          4213 => x"ae",
          4214 => x"34",
          4215 => x"0b",
          4216 => x"76",
          4217 => x"18",
          4218 => x"8f",
          4219 => x"b4",
          4220 => x"51",
          4221 => x"a0",
          4222 => x"52",
          4223 => x"51",
          4224 => x"3f",
          4225 => x"0b",
          4226 => x"34",
          4227 => x"d4",
          4228 => x"51",
          4229 => x"77",
          4230 => x"83",
          4231 => x"3d",
          4232 => x"c5",
          4233 => x"d3",
          4234 => x"91",
          4235 => x"af",
          4236 => x"63",
          4237 => x"ff",
          4238 => x"75",
          4239 => x"77",
          4240 => x"3f",
          4241 => x"0b",
          4242 => x"77",
          4243 => x"83",
          4244 => x"51",
          4245 => x"3f",
          4246 => x"08",
          4247 => x"80",
          4248 => x"98",
          4249 => x"51",
          4250 => x"3f",
          4251 => x"c8",
          4252 => x"0d",
          4253 => x"0d",
          4254 => x"05",
          4255 => x"3f",
          4256 => x"3d",
          4257 => x"52",
          4258 => x"d0",
          4259 => x"d3",
          4260 => x"91",
          4261 => x"82",
          4262 => x"4c",
          4263 => x"52",
          4264 => x"05",
          4265 => x"3f",
          4266 => x"08",
          4267 => x"c8",
          4268 => x"38",
          4269 => x"05",
          4270 => x"06",
          4271 => x"2e",
          4272 => x"55",
          4273 => x"38",
          4274 => x"3d",
          4275 => x"3d",
          4276 => x"51",
          4277 => x"3f",
          4278 => x"3d",
          4279 => x"91",
          4280 => x"54",
          4281 => x"3f",
          4282 => x"52",
          4283 => x"9e",
          4284 => x"c8",
          4285 => x"d3",
          4286 => x"38",
          4287 => x"09",
          4288 => x"38",
          4289 => x"a1",
          4290 => x"83",
          4291 => x"74",
          4292 => x"81",
          4293 => x"38",
          4294 => x"a8",
          4295 => x"ec",
          4296 => x"c8",
          4297 => x"d3",
          4298 => x"c4",
          4299 => x"93",
          4300 => x"ff",
          4301 => x"8d",
          4302 => x"ac",
          4303 => x"ab",
          4304 => x"17",
          4305 => x"33",
          4306 => x"70",
          4307 => x"55",
          4308 => x"38",
          4309 => x"54",
          4310 => x"34",
          4311 => x"0b",
          4312 => x"8b",
          4313 => x"84",
          4314 => x"06",
          4315 => x"73",
          4316 => x"db",
          4317 => x"2e",
          4318 => x"75",
          4319 => x"ff",
          4320 => x"91",
          4321 => x"52",
          4322 => x"b0",
          4323 => x"55",
          4324 => x"08",
          4325 => x"38",
          4326 => x"08",
          4327 => x"ff",
          4328 => x"91",
          4329 => x"80",
          4330 => x"55",
          4331 => x"08",
          4332 => x"16",
          4333 => x"ae",
          4334 => x"06",
          4335 => x"53",
          4336 => x"51",
          4337 => x"3f",
          4338 => x"0b",
          4339 => x"74",
          4340 => x"3d",
          4341 => x"c3",
          4342 => x"d3",
          4343 => x"91",
          4344 => x"8c",
          4345 => x"ff",
          4346 => x"91",
          4347 => x"55",
          4348 => x"c8",
          4349 => x"0d",
          4350 => x"0d",
          4351 => x"05",
          4352 => x"05",
          4353 => x"33",
          4354 => x"53",
          4355 => x"05",
          4356 => x"51",
          4357 => x"91",
          4358 => x"55",
          4359 => x"08",
          4360 => x"78",
          4361 => x"95",
          4362 => x"51",
          4363 => x"91",
          4364 => x"55",
          4365 => x"08",
          4366 => x"80",
          4367 => x"81",
          4368 => x"73",
          4369 => x"38",
          4370 => x"aa",
          4371 => x"06",
          4372 => x"8b",
          4373 => x"06",
          4374 => x"07",
          4375 => x"56",
          4376 => x"34",
          4377 => x"0b",
          4378 => x"78",
          4379 => x"a0",
          4380 => x"c8",
          4381 => x"91",
          4382 => x"95",
          4383 => x"ee",
          4384 => x"56",
          4385 => x"3d",
          4386 => x"95",
          4387 => x"ce",
          4388 => x"c8",
          4389 => x"d3",
          4390 => x"d3",
          4391 => x"64",
          4392 => x"d4",
          4393 => x"e6",
          4394 => x"c8",
          4395 => x"d3",
          4396 => x"38",
          4397 => x"05",
          4398 => x"06",
          4399 => x"2e",
          4400 => x"55",
          4401 => x"86",
          4402 => x"17",
          4403 => x"2b",
          4404 => x"57",
          4405 => x"05",
          4406 => x"9f",
          4407 => x"81",
          4408 => x"34",
          4409 => x"ac",
          4410 => x"d3",
          4411 => x"74",
          4412 => x"0c",
          4413 => x"04",
          4414 => x"69",
          4415 => x"80",
          4416 => x"d0",
          4417 => x"3d",
          4418 => x"3f",
          4419 => x"08",
          4420 => x"08",
          4421 => x"d3",
          4422 => x"80",
          4423 => x"70",
          4424 => x"2a",
          4425 => x"57",
          4426 => x"74",
          4427 => x"f6",
          4428 => x"80",
          4429 => x"8d",
          4430 => x"54",
          4431 => x"3f",
          4432 => x"08",
          4433 => x"c8",
          4434 => x"38",
          4435 => x"51",
          4436 => x"3f",
          4437 => x"08",
          4438 => x"c8",
          4439 => x"91",
          4440 => x"91",
          4441 => x"65",
          4442 => x"79",
          4443 => x"7a",
          4444 => x"55",
          4445 => x"34",
          4446 => x"8a",
          4447 => x"38",
          4448 => x"80",
          4449 => x"80",
          4450 => x"ff",
          4451 => x"70",
          4452 => x"58",
          4453 => x"e8",
          4454 => x"2e",
          4455 => x"86",
          4456 => x"34",
          4457 => x"30",
          4458 => x"80",
          4459 => x"70",
          4460 => x"2a",
          4461 => x"56",
          4462 => x"80",
          4463 => x"7b",
          4464 => x"53",
          4465 => x"81",
          4466 => x"c8",
          4467 => x"d3",
          4468 => x"38",
          4469 => x"51",
          4470 => x"58",
          4471 => x"8b",
          4472 => x"58",
          4473 => x"83",
          4474 => x"7b",
          4475 => x"51",
          4476 => x"3f",
          4477 => x"08",
          4478 => x"91",
          4479 => x"98",
          4480 => x"e8",
          4481 => x"53",
          4482 => x"b8",
          4483 => x"3d",
          4484 => x"3f",
          4485 => x"08",
          4486 => x"c8",
          4487 => x"38",
          4488 => x"52",
          4489 => x"bc",
          4490 => x"a7",
          4491 => x"6b",
          4492 => x"52",
          4493 => x"9f",
          4494 => x"b5",
          4495 => x"6b",
          4496 => x"70",
          4497 => x"52",
          4498 => x"fe",
          4499 => x"c8",
          4500 => x"a2",
          4501 => x"33",
          4502 => x"54",
          4503 => x"3f",
          4504 => x"08",
          4505 => x"38",
          4506 => x"74",
          4507 => x"05",
          4508 => x"39",
          4509 => x"9f",
          4510 => x"99",
          4511 => x"e0",
          4512 => x"ff",
          4513 => x"54",
          4514 => x"27",
          4515 => x"ba",
          4516 => x"56",
          4517 => x"a3",
          4518 => x"91",
          4519 => x"ff",
          4520 => x"91",
          4521 => x"93",
          4522 => x"76",
          4523 => x"76",
          4524 => x"38",
          4525 => x"77",
          4526 => x"86",
          4527 => x"39",
          4528 => x"27",
          4529 => x"3d",
          4530 => x"bc",
          4531 => x"2a",
          4532 => x"75",
          4533 => x"57",
          4534 => x"05",
          4535 => x"54",
          4536 => x"81",
          4537 => x"33",
          4538 => x"73",
          4539 => x"cd",
          4540 => x"33",
          4541 => x"73",
          4542 => x"81",
          4543 => x"80",
          4544 => x"02",
          4545 => x"78",
          4546 => x"51",
          4547 => x"73",
          4548 => x"81",
          4549 => x"ff",
          4550 => x"80",
          4551 => x"76",
          4552 => x"51",
          4553 => x"2e",
          4554 => x"5f",
          4555 => x"52",
          4556 => x"52",
          4557 => x"c2",
          4558 => x"c8",
          4559 => x"d3",
          4560 => x"a1",
          4561 => x"74",
          4562 => x"82",
          4563 => x"c8",
          4564 => x"d3",
          4565 => x"38",
          4566 => x"91",
          4567 => x"9a",
          4568 => x"05",
          4569 => x"ff",
          4570 => x"86",
          4571 => x"e5",
          4572 => x"54",
          4573 => x"15",
          4574 => x"ff",
          4575 => x"91",
          4576 => x"54",
          4577 => x"91",
          4578 => x"84",
          4579 => x"06",
          4580 => x"80",
          4581 => x"2e",
          4582 => x"81",
          4583 => x"d4",
          4584 => x"b6",
          4585 => x"d3",
          4586 => x"91",
          4587 => x"b5",
          4588 => x"91",
          4589 => x"52",
          4590 => x"a4",
          4591 => x"54",
          4592 => x"15",
          4593 => x"9a",
          4594 => x"05",
          4595 => x"ff",
          4596 => x"77",
          4597 => x"83",
          4598 => x"51",
          4599 => x"3f",
          4600 => x"08",
          4601 => x"74",
          4602 => x"0c",
          4603 => x"04",
          4604 => x"61",
          4605 => x"05",
          4606 => x"33",
          4607 => x"05",
          4608 => x"5e",
          4609 => x"a2",
          4610 => x"c8",
          4611 => x"d3",
          4612 => x"38",
          4613 => x"57",
          4614 => x"86",
          4615 => x"82",
          4616 => x"80",
          4617 => x"8c",
          4618 => x"38",
          4619 => x"70",
          4620 => x"81",
          4621 => x"55",
          4622 => x"87",
          4623 => x"39",
          4624 => x"89",
          4625 => x"81",
          4626 => x"8a",
          4627 => x"89",
          4628 => x"7d",
          4629 => x"54",
          4630 => x"3f",
          4631 => x"06",
          4632 => x"72",
          4633 => x"91",
          4634 => x"05",
          4635 => x"08",
          4636 => x"55",
          4637 => x"81",
          4638 => x"38",
          4639 => x"79",
          4640 => x"82",
          4641 => x"56",
          4642 => x"74",
          4643 => x"ff",
          4644 => x"91",
          4645 => x"81",
          4646 => x"56",
          4647 => x"08",
          4648 => x"38",
          4649 => x"81",
          4650 => x"38",
          4651 => x"ff",
          4652 => x"8b",
          4653 => x"5a",
          4654 => x"91",
          4655 => x"74",
          4656 => x"74",
          4657 => x"81",
          4658 => x"87",
          4659 => x"86",
          4660 => x"2e",
          4661 => x"7e",
          4662 => x"80",
          4663 => x"81",
          4664 => x"81",
          4665 => x"06",
          4666 => x"54",
          4667 => x"52",
          4668 => x"a7",
          4669 => x"d3",
          4670 => x"91",
          4671 => x"91",
          4672 => x"16",
          4673 => x"56",
          4674 => x"38",
          4675 => x"1d",
          4676 => x"c2",
          4677 => x"8c",
          4678 => x"7b",
          4679 => x"38",
          4680 => x"0c",
          4681 => x"0c",
          4682 => x"80",
          4683 => x"73",
          4684 => x"7f",
          4685 => x"fe",
          4686 => x"90",
          4687 => x"26",
          4688 => x"15",
          4689 => x"90",
          4690 => x"84",
          4691 => x"07",
          4692 => x"84",
          4693 => x"54",
          4694 => x"c8",
          4695 => x"0d",
          4696 => x"0d",
          4697 => x"05",
          4698 => x"33",
          4699 => x"5e",
          4700 => x"d3",
          4701 => x"c8",
          4702 => x"57",
          4703 => x"d3",
          4704 => x"8c",
          4705 => x"d3",
          4706 => x"10",
          4707 => x"05",
          4708 => x"80",
          4709 => x"74",
          4710 => x"75",
          4711 => x"ff",
          4712 => x"52",
          4713 => x"99",
          4714 => x"d3",
          4715 => x"ff",
          4716 => x"06",
          4717 => x"57",
          4718 => x"38",
          4719 => x"70",
          4720 => x"55",
          4721 => x"8c",
          4722 => x"3d",
          4723 => x"83",
          4724 => x"ff",
          4725 => x"91",
          4726 => x"98",
          4727 => x"2e",
          4728 => x"82",
          4729 => x"8c",
          4730 => x"05",
          4731 => x"74",
          4732 => x"38",
          4733 => x"80",
          4734 => x"2e",
          4735 => x"78",
          4736 => x"77",
          4737 => x"26",
          4738 => x"18",
          4739 => x"74",
          4740 => x"38",
          4741 => x"be",
          4742 => x"77",
          4743 => x"98",
          4744 => x"c8",
          4745 => x"54",
          4746 => x"58",
          4747 => x"3f",
          4748 => x"08",
          4749 => x"c8",
          4750 => x"30",
          4751 => x"80",
          4752 => x"c8",
          4753 => x"91",
          4754 => x"07",
          4755 => x"07",
          4756 => x"58",
          4757 => x"57",
          4758 => x"38",
          4759 => x"05",
          4760 => x"79",
          4761 => x"cb",
          4762 => x"91",
          4763 => x"8a",
          4764 => x"83",
          4765 => x"06",
          4766 => x"44",
          4767 => x"09",
          4768 => x"38",
          4769 => x"57",
          4770 => x"8a",
          4771 => x"64",
          4772 => x"57",
          4773 => x"27",
          4774 => x"93",
          4775 => x"80",
          4776 => x"38",
          4777 => x"70",
          4778 => x"55",
          4779 => x"95",
          4780 => x"06",
          4781 => x"2e",
          4782 => x"81",
          4783 => x"85",
          4784 => x"8f",
          4785 => x"06",
          4786 => x"82",
          4787 => x"2e",
          4788 => x"77",
          4789 => x"2e",
          4790 => x"80",
          4791 => x"b4",
          4792 => x"2a",
          4793 => x"81",
          4794 => x"9c",
          4795 => x"52",
          4796 => x"74",
          4797 => x"38",
          4798 => x"98",
          4799 => x"79",
          4800 => x"18",
          4801 => x"57",
          4802 => x"80",
          4803 => x"76",
          4804 => x"38",
          4805 => x"51",
          4806 => x"3f",
          4807 => x"08",
          4808 => x"08",
          4809 => x"7f",
          4810 => x"52",
          4811 => x"88",
          4812 => x"c8",
          4813 => x"5b",
          4814 => x"80",
          4815 => x"43",
          4816 => x"0a",
          4817 => x"8b",
          4818 => x"89",
          4819 => x"b4",
          4820 => x"2a",
          4821 => x"81",
          4822 => x"8c",
          4823 => x"52",
          4824 => x"74",
          4825 => x"38",
          4826 => x"98",
          4827 => x"79",
          4828 => x"18",
          4829 => x"57",
          4830 => x"80",
          4831 => x"76",
          4832 => x"38",
          4833 => x"51",
          4834 => x"3f",
          4835 => x"08",
          4836 => x"57",
          4837 => x"08",
          4838 => x"92",
          4839 => x"91",
          4840 => x"83",
          4841 => x"72",
          4842 => x"51",
          4843 => x"52",
          4844 => x"05",
          4845 => x"80",
          4846 => x"c8",
          4847 => x"7e",
          4848 => x"80",
          4849 => x"f2",
          4850 => x"d3",
          4851 => x"ff",
          4852 => x"63",
          4853 => x"64",
          4854 => x"ff",
          4855 => x"70",
          4856 => x"31",
          4857 => x"57",
          4858 => x"2e",
          4859 => x"89",
          4860 => x"60",
          4861 => x"84",
          4862 => x"5c",
          4863 => x"16",
          4864 => x"51",
          4865 => x"26",
          4866 => x"65",
          4867 => x"31",
          4868 => x"64",
          4869 => x"fe",
          4870 => x"91",
          4871 => x"56",
          4872 => x"09",
          4873 => x"38",
          4874 => x"08",
          4875 => x"26",
          4876 => x"89",
          4877 => x"2a",
          4878 => x"97",
          4879 => x"87",
          4880 => x"82",
          4881 => x"06",
          4882 => x"83",
          4883 => x"27",
          4884 => x"8f",
          4885 => x"55",
          4886 => x"26",
          4887 => x"58",
          4888 => x"7c",
          4889 => x"06",
          4890 => x"2e",
          4891 => x"42",
          4892 => x"77",
          4893 => x"19",
          4894 => x"78",
          4895 => x"38",
          4896 => x"d2",
          4897 => x"f5",
          4898 => x"77",
          4899 => x"19",
          4900 => x"78",
          4901 => x"38",
          4902 => x"ba",
          4903 => x"61",
          4904 => x"81",
          4905 => x"61",
          4906 => x"f5",
          4907 => x"55",
          4908 => x"86",
          4909 => x"53",
          4910 => x"51",
          4911 => x"3f",
          4912 => x"bb",
          4913 => x"51",
          4914 => x"3f",
          4915 => x"1f",
          4916 => x"89",
          4917 => x"8d",
          4918 => x"83",
          4919 => x"52",
          4920 => x"ff",
          4921 => x"81",
          4922 => x"34",
          4923 => x"70",
          4924 => x"2a",
          4925 => x"54",
          4926 => x"1f",
          4927 => x"dd",
          4928 => x"ff",
          4929 => x"38",
          4930 => x"05",
          4931 => x"1f",
          4932 => x"c9",
          4933 => x"65",
          4934 => x"51",
          4935 => x"3f",
          4936 => x"05",
          4937 => x"98",
          4938 => x"98",
          4939 => x"ff",
          4940 => x"51",
          4941 => x"3f",
          4942 => x"1f",
          4943 => x"bb",
          4944 => x"2e",
          4945 => x"80",
          4946 => x"88",
          4947 => x"80",
          4948 => x"ff",
          4949 => x"7b",
          4950 => x"51",
          4951 => x"3f",
          4952 => x"1f",
          4953 => x"93",
          4954 => x"b0",
          4955 => x"97",
          4956 => x"52",
          4957 => x"ff",
          4958 => x"ff",
          4959 => x"c0",
          4960 => x"7f",
          4961 => x"34",
          4962 => x"bb",
          4963 => x"c7",
          4964 => x"98",
          4965 => x"39",
          4966 => x"0a",
          4967 => x"51",
          4968 => x"3f",
          4969 => x"ff",
          4970 => x"1f",
          4971 => x"ad",
          4972 => x"7f",
          4973 => x"a9",
          4974 => x"34",
          4975 => x"bb",
          4976 => x"1f",
          4977 => x"e2",
          4978 => x"d5",
          4979 => x"1f",
          4980 => x"89",
          4981 => x"63",
          4982 => x"79",
          4983 => x"f9",
          4984 => x"91",
          4985 => x"83",
          4986 => x"83",
          4987 => x"06",
          4988 => x"81",
          4989 => x"05",
          4990 => x"79",
          4991 => x"d9",
          4992 => x"80",
          4993 => x"ff",
          4994 => x"84",
          4995 => x"d2",
          4996 => x"ff",
          4997 => x"86",
          4998 => x"f2",
          4999 => x"1f",
          5000 => x"d7",
          5001 => x"52",
          5002 => x"51",
          5003 => x"3f",
          5004 => x"ec",
          5005 => x"96",
          5006 => x"d4",
          5007 => x"fe",
          5008 => x"96",
          5009 => x"54",
          5010 => x"53",
          5011 => x"51",
          5012 => x"3f",
          5013 => x"81",
          5014 => x"52",
          5015 => x"92",
          5016 => x"53",
          5017 => x"51",
          5018 => x"3f",
          5019 => x"5b",
          5020 => x"09",
          5021 => x"38",
          5022 => x"51",
          5023 => x"3f",
          5024 => x"1f",
          5025 => x"f3",
          5026 => x"52",
          5027 => x"ff",
          5028 => x"95",
          5029 => x"ff",
          5030 => x"81",
          5031 => x"f8",
          5032 => x"7e",
          5033 => x"d3",
          5034 => x"60",
          5035 => x"26",
          5036 => x"57",
          5037 => x"53",
          5038 => x"51",
          5039 => x"3f",
          5040 => x"08",
          5041 => x"7d",
          5042 => x"7e",
          5043 => x"fe",
          5044 => x"75",
          5045 => x"56",
          5046 => x"81",
          5047 => x"80",
          5048 => x"38",
          5049 => x"83",
          5050 => x"62",
          5051 => x"74",
          5052 => x"38",
          5053 => x"54",
          5054 => x"52",
          5055 => x"91",
          5056 => x"d3",
          5057 => x"c8",
          5058 => x"75",
          5059 => x"56",
          5060 => x"8c",
          5061 => x"2e",
          5062 => x"57",
          5063 => x"ff",
          5064 => x"84",
          5065 => x"2e",
          5066 => x"57",
          5067 => x"81",
          5068 => x"80",
          5069 => x"53",
          5070 => x"51",
          5071 => x"3f",
          5072 => x"52",
          5073 => x"51",
          5074 => x"3f",
          5075 => x"56",
          5076 => x"81",
          5077 => x"34",
          5078 => x"17",
          5079 => x"17",
          5080 => x"17",
          5081 => x"05",
          5082 => x"c1",
          5083 => x"fe",
          5084 => x"fe",
          5085 => x"34",
          5086 => x"08",
          5087 => x"07",
          5088 => x"17",
          5089 => x"c8",
          5090 => x"34",
          5091 => x"c6",
          5092 => x"93",
          5093 => x"52",
          5094 => x"51",
          5095 => x"3f",
          5096 => x"53",
          5097 => x"51",
          5098 => x"3f",
          5099 => x"d3",
          5100 => x"38",
          5101 => x"52",
          5102 => x"91",
          5103 => x"57",
          5104 => x"08",
          5105 => x"39",
          5106 => x"39",
          5107 => x"39",
          5108 => x"39",
          5109 => x"91",
          5110 => x"98",
          5111 => x"ff",
          5112 => x"52",
          5113 => x"81",
          5114 => x"10",
          5115 => x"b8",
          5116 => x"08",
          5117 => x"f8",
          5118 => x"a9",
          5119 => x"39",
          5120 => x"51",
          5121 => x"3f",
          5122 => x"91",
          5123 => x"ff",
          5124 => x"81",
          5125 => x"c2",
          5126 => x"80",
          5127 => x"b3",
          5128 => x"bc",
          5129 => x"fd",
          5130 => x"39",
          5131 => x"51",
          5132 => x"3f",
          5133 => x"91",
          5134 => x"fe",
          5135 => x"81",
          5136 => x"c2",
          5137 => x"ff",
          5138 => x"87",
          5139 => x"88",
          5140 => x"d1",
          5141 => x"39",
          5142 => x"51",
          5143 => x"3f",
          5144 => x"91",
          5145 => x"fe",
          5146 => x"80",
          5147 => x"c3",
          5148 => x"ff",
          5149 => x"db",
          5150 => x"e8",
          5151 => x"a5",
          5152 => x"39",
          5153 => x"51",
          5154 => x"3f",
          5155 => x"91",
          5156 => x"fe",
          5157 => x"bb",
          5158 => x"c8",
          5159 => x"85",
          5160 => x"91",
          5161 => x"fe",
          5162 => x"a7",
          5163 => x"f4",
          5164 => x"f1",
          5165 => x"91",
          5166 => x"fe",
          5167 => x"93",
          5168 => x"a4",
          5169 => x"dd",
          5170 => x"91",
          5171 => x"fe",
          5172 => x"83",
          5173 => x"fb",
          5174 => x"79",
          5175 => x"87",
          5176 => x"38",
          5177 => x"87",
          5178 => x"fe",
          5179 => x"91",
          5180 => x"55",
          5181 => x"e8",
          5182 => x"fe",
          5183 => x"91",
          5184 => x"52",
          5185 => x"e8",
          5186 => x"d3",
          5187 => x"74",
          5188 => x"75",
          5189 => x"c0",
          5190 => x"83",
          5191 => x"0d",
          5192 => x"3d",
          5193 => x"3d",
          5194 => x"3d",
          5195 => x"05",
          5196 => x"33",
          5197 => x"70",
          5198 => x"25",
          5199 => x"27",
          5200 => x"5a",
          5201 => x"93",
          5202 => x"87",
          5203 => x"77",
          5204 => x"3d",
          5205 => x"51",
          5206 => x"3f",
          5207 => x"08",
          5208 => x"c8",
          5209 => x"91",
          5210 => x"87",
          5211 => x"0c",
          5212 => x"08",
          5213 => x"3d",
          5214 => x"55",
          5215 => x"53",
          5216 => x"d8",
          5217 => x"f2",
          5218 => x"c8",
          5219 => x"d3",
          5220 => x"38",
          5221 => x"89",
          5222 => x"7b",
          5223 => x"d5",
          5224 => x"3d",
          5225 => x"51",
          5226 => x"77",
          5227 => x"07",
          5228 => x"30",
          5229 => x"72",
          5230 => x"51",
          5231 => x"2e",
          5232 => x"c5",
          5233 => x"c0",
          5234 => x"52",
          5235 => x"87",
          5236 => x"74",
          5237 => x"0c",
          5238 => x"0d",
          5239 => x"0d",
          5240 => x"33",
          5241 => x"57",
          5242 => x"7b",
          5243 => x"fe",
          5244 => x"d3",
          5245 => x"38",
          5246 => x"88",
          5247 => x"2e",
          5248 => x"39",
          5249 => x"54",
          5250 => x"53",
          5251 => x"51",
          5252 => x"d3",
          5253 => x"83",
          5254 => x"78",
          5255 => x"0c",
          5256 => x"04",
          5257 => x"02",
          5258 => x"91",
          5259 => x"91",
          5260 => x"56",
          5261 => x"3f",
          5262 => x"70",
          5263 => x"fe",
          5264 => x"91",
          5265 => x"91",
          5266 => x"81",
          5267 => x"91",
          5268 => x"ff",
          5269 => x"75",
          5270 => x"38",
          5271 => x"3f",
          5272 => x"04",
          5273 => x"87",
          5274 => x"08",
          5275 => x"ff",
          5276 => x"fe",
          5277 => x"91",
          5278 => x"fe",
          5279 => x"80",
          5280 => x"f1",
          5281 => x"2a",
          5282 => x"51",
          5283 => x"2e",
          5284 => x"51",
          5285 => x"3f",
          5286 => x"51",
          5287 => x"3f",
          5288 => x"ee",
          5289 => x"82",
          5290 => x"06",
          5291 => x"80",
          5292 => x"81",
          5293 => x"bd",
          5294 => x"e0",
          5295 => x"b3",
          5296 => x"fe",
          5297 => x"72",
          5298 => x"81",
          5299 => x"71",
          5300 => x"38",
          5301 => x"ee",
          5302 => x"c6",
          5303 => x"f0",
          5304 => x"51",
          5305 => x"3f",
          5306 => x"70",
          5307 => x"52",
          5308 => x"95",
          5309 => x"fe",
          5310 => x"91",
          5311 => x"fe",
          5312 => x"80",
          5313 => x"ed",
          5314 => x"2a",
          5315 => x"51",
          5316 => x"2e",
          5317 => x"51",
          5318 => x"3f",
          5319 => x"51",
          5320 => x"3f",
          5321 => x"ed",
          5322 => x"86",
          5323 => x"06",
          5324 => x"80",
          5325 => x"81",
          5326 => x"b9",
          5327 => x"ac",
          5328 => x"af",
          5329 => x"fe",
          5330 => x"72",
          5331 => x"81",
          5332 => x"71",
          5333 => x"38",
          5334 => x"ed",
          5335 => x"c7",
          5336 => x"ef",
          5337 => x"51",
          5338 => x"3f",
          5339 => x"70",
          5340 => x"52",
          5341 => x"95",
          5342 => x"fe",
          5343 => x"91",
          5344 => x"fe",
          5345 => x"80",
          5346 => x"e9",
          5347 => x"a8",
          5348 => x"0d",
          5349 => x"0d",
          5350 => x"70",
          5351 => x"74",
          5352 => x"ed",
          5353 => x"74",
          5354 => x"14",
          5355 => x"e1",
          5356 => x"55",
          5357 => x"54",
          5358 => x"2e",
          5359 => x"54",
          5360 => x"9f",
          5361 => x"51",
          5362 => x"38",
          5363 => x"72",
          5364 => x"81",
          5365 => x"80",
          5366 => x"05",
          5367 => x"56",
          5368 => x"91",
          5369 => x"77",
          5370 => x"08",
          5371 => x"e6",
          5372 => x"d3",
          5373 => x"38",
          5374 => x"53",
          5375 => x"ff",
          5376 => x"16",
          5377 => x"06",
          5378 => x"76",
          5379 => x"ff",
          5380 => x"d3",
          5381 => x"3d",
          5382 => x"3d",
          5383 => x"91",
          5384 => x"71",
          5385 => x"5c",
          5386 => x"52",
          5387 => x"84",
          5388 => x"d3",
          5389 => x"ff",
          5390 => x"7c",
          5391 => x"06",
          5392 => x"c8",
          5393 => x"3d",
          5394 => x"fe",
          5395 => x"7b",
          5396 => x"ea",
          5397 => x"ff",
          5398 => x"91",
          5399 => x"5a",
          5400 => x"8b",
          5401 => x"98",
          5402 => x"b3",
          5403 => x"81",
          5404 => x"91",
          5405 => x"fe",
          5406 => x"96",
          5407 => x"59",
          5408 => x"54",
          5409 => x"78",
          5410 => x"a4",
          5411 => x"61",
          5412 => x"e5",
          5413 => x"fe",
          5414 => x"fd",
          5415 => x"d3",
          5416 => x"2b",
          5417 => x"51",
          5418 => x"87",
          5419 => x"38",
          5420 => x"91",
          5421 => x"59",
          5422 => x"b4",
          5423 => x"11",
          5424 => x"05",
          5425 => x"e2",
          5426 => x"c8",
          5427 => x"91",
          5428 => x"fe",
          5429 => x"ff",
          5430 => x"3d",
          5431 => x"53",
          5432 => x"51",
          5433 => x"3f",
          5434 => x"08",
          5435 => x"38",
          5436 => x"83",
          5437 => x"02",
          5438 => x"52",
          5439 => x"05",
          5440 => x"82",
          5441 => x"d3",
          5442 => x"ff",
          5443 => x"8e",
          5444 => x"e4",
          5445 => x"8d",
          5446 => x"fe",
          5447 => x"c8",
          5448 => x"f6",
          5449 => x"cb",
          5450 => x"fe",
          5451 => x"fe",
          5452 => x"fe",
          5453 => x"91",
          5454 => x"80",
          5455 => x"38",
          5456 => x"52",
          5457 => x"05",
          5458 => x"86",
          5459 => x"d3",
          5460 => x"91",
          5461 => x"fe",
          5462 => x"fe",
          5463 => x"3d",
          5464 => x"53",
          5465 => x"51",
          5466 => x"3f",
          5467 => x"08",
          5468 => x"38",
          5469 => x"fd",
          5470 => x"3d",
          5471 => x"53",
          5472 => x"51",
          5473 => x"3f",
          5474 => x"08",
          5475 => x"d3",
          5476 => x"60",
          5477 => x"94",
          5478 => x"70",
          5479 => x"fb",
          5480 => x"bf",
          5481 => x"78",
          5482 => x"b4",
          5483 => x"f8",
          5484 => x"b2",
          5485 => x"d3",
          5486 => x"2e",
          5487 => x"d3",
          5488 => x"f4",
          5489 => x"ab",
          5490 => x"e4",
          5491 => x"d5",
          5492 => x"fd",
          5493 => x"3d",
          5494 => x"51",
          5495 => x"3f",
          5496 => x"08",
          5497 => x"f8",
          5498 => x"fe",
          5499 => x"81",
          5500 => x"c8",
          5501 => x"51",
          5502 => x"91",
          5503 => x"80",
          5504 => x"38",
          5505 => x"08",
          5506 => x"3f",
          5507 => x"b4",
          5508 => x"05",
          5509 => x"eb",
          5510 => x"c8",
          5511 => x"fe",
          5512 => x"5b",
          5513 => x"3f",
          5514 => x"08",
          5515 => x"f8",
          5516 => x"fe",
          5517 => x"91",
          5518 => x"b5",
          5519 => x"05",
          5520 => x"e4",
          5521 => x"cb",
          5522 => x"d3",
          5523 => x"56",
          5524 => x"d3",
          5525 => x"ff",
          5526 => x"53",
          5527 => x"51",
          5528 => x"91",
          5529 => x"80",
          5530 => x"38",
          5531 => x"08",
          5532 => x"3f",
          5533 => x"91",
          5534 => x"fe",
          5535 => x"82",
          5536 => x"8f",
          5537 => x"39",
          5538 => x"51",
          5539 => x"3f",
          5540 => x"f1",
          5541 => x"db",
          5542 => x"81",
          5543 => x"94",
          5544 => x"80",
          5545 => x"c0",
          5546 => x"91",
          5547 => x"fe",
          5548 => x"fb",
          5549 => x"c9",
          5550 => x"f2",
          5551 => x"80",
          5552 => x"c0",
          5553 => x"8c",
          5554 => x"87",
          5555 => x"0c",
          5556 => x"b4",
          5557 => x"11",
          5558 => x"05",
          5559 => x"ca",
          5560 => x"c8",
          5561 => x"fb",
          5562 => x"52",
          5563 => x"51",
          5564 => x"3f",
          5565 => x"04",
          5566 => x"f4",
          5567 => x"f8",
          5568 => x"fa",
          5569 => x"d3",
          5570 => x"2e",
          5571 => x"60",
          5572 => x"8c",
          5573 => x"87",
          5574 => x"78",
          5575 => x"c8",
          5576 => x"d3",
          5577 => x"2e",
          5578 => x"91",
          5579 => x"52",
          5580 => x"51",
          5581 => x"3f",
          5582 => x"91",
          5583 => x"fe",
          5584 => x"fe",
          5585 => x"fa",
          5586 => x"ca",
          5587 => x"f1",
          5588 => x"59",
          5589 => x"fe",
          5590 => x"fa",
          5591 => x"70",
          5592 => x"78",
          5593 => x"8b",
          5594 => x"06",
          5595 => x"2e",
          5596 => x"b4",
          5597 => x"05",
          5598 => x"87",
          5599 => x"f4",
          5600 => x"c8",
          5601 => x"ca",
          5602 => x"53",
          5603 => x"52",
          5604 => x"52",
          5605 => x"9d",
          5606 => x"c4",
          5607 => x"fc",
          5608 => x"61",
          5609 => x"61",
          5610 => x"83",
          5611 => x"83",
          5612 => x"78",
          5613 => x"3f",
          5614 => x"08",
          5615 => x"32",
          5616 => x"07",
          5617 => x"38",
          5618 => x"09",
          5619 => x"a3",
          5620 => x"8c",
          5621 => x"c7",
          5622 => x"39",
          5623 => x"80",
          5624 => x"fc",
          5625 => x"86",
          5626 => x"c0",
          5627 => x"9b",
          5628 => x"0b",
          5629 => x"9c",
          5630 => x"83",
          5631 => x"94",
          5632 => x"80",
          5633 => x"c0",
          5634 => x"90",
          5635 => x"91",
          5636 => x"90",
          5637 => x"91",
          5638 => x"fe",
          5639 => x"fe",
          5640 => x"91",
          5641 => x"fe",
          5642 => x"91",
          5643 => x"fe",
          5644 => x"91",
          5645 => x"fe",
          5646 => x"81",
          5647 => x"3f",
          5648 => x"80",
          5649 => x"04",
          5650 => x"04",
          5651 => x"04",
          5652 => x"04",
          5653 => x"04",
          5654 => x"04",
          5655 => x"04",
          5656 => x"04",
          5657 => x"04",
          5658 => x"04",
          5659 => x"04",
          5660 => x"04",
          5661 => x"04",
          5662 => x"04",
          5663 => x"04",
          5664 => x"04",
          5665 => x"04",
          5666 => x"04",
          5667 => x"04",
          5668 => x"04",
          5669 => x"04",
          5670 => x"04",
          5671 => x"04",
          5672 => x"04",
          5673 => x"04",
          5674 => x"04",
          5675 => x"04",
          5676 => x"04",
          5677 => x"04",
          5678 => x"04",
          5679 => x"04",
          5680 => x"04",
          5681 => x"04",
          5682 => x"04",
          5683 => x"04",
          5684 => x"04",
          5685 => x"04",
          5686 => x"04",
          5687 => x"04",
          5688 => x"04",
          5689 => x"04",
          5690 => x"04",
          5691 => x"04",
          5692 => x"04",
          5693 => x"04",
          5694 => x"04",
          5695 => x"04",
          5696 => x"04",
          5697 => x"04",
          5698 => x"04",
          5699 => x"04",
          5700 => x"04",
          5701 => x"04",
          5702 => x"04",
          5703 => x"04",
          5704 => x"04",
          5705 => x"04",
          5706 => x"04",
          5707 => x"04",
          5708 => x"04",
          5709 => x"04",
          5710 => x"04",
          5711 => x"04",
          5712 => x"04",
          5713 => x"04",
          5714 => x"04",
          5715 => x"04",
          5716 => x"04",
          5717 => x"04",
          5718 => x"04",
          5719 => x"04",
          5720 => x"04",
          5721 => x"04",
          5722 => x"04",
          5723 => x"04",
          5724 => x"04",
          5725 => x"04",
          5726 => x"04",
          5727 => x"04",
          5728 => x"04",
          5729 => x"04",
          5730 => x"04",
          5731 => x"04",
          5732 => x"04",
          5733 => x"04",
          5734 => x"04",
          5735 => x"04",
          5736 => x"04",
          5737 => x"04",
          5738 => x"04",
          5739 => x"04",
          5740 => x"04",
          5741 => x"04",
          5742 => x"04",
          5743 => x"04",
          5744 => x"04",
          5745 => x"04",
          5746 => x"04",
          5747 => x"04",
          5748 => x"04",
          5749 => x"04",
          5750 => x"04",
          5751 => x"04",
          5752 => x"04",
          5753 => x"04",
          5754 => x"04",
          5755 => x"04",
          5756 => x"04",
          5757 => x"04",
          5758 => x"04",
          5759 => x"04",
          5760 => x"04",
          5761 => x"04",
          5762 => x"04",
          5763 => x"04",
          5764 => x"04",
          5765 => x"04",
          5766 => x"04",
          5767 => x"04",
          5768 => x"04",
          5769 => x"04",
          5770 => x"04",
          5771 => x"04",
          5772 => x"04",
          5773 => x"04",
          5774 => x"04",
          5775 => x"04",
          5776 => x"04",
          5777 => x"04",
          5778 => x"04",
          5779 => x"04",
          5780 => x"04",
          5781 => x"04",
          5782 => x"04",
          5783 => x"04",
          5784 => x"04",
          5785 => x"04",
          5786 => x"04",
          5787 => x"04",
          5788 => x"04",
          5789 => x"04",
          5790 => x"04",
          5791 => x"04",
          5792 => x"04",
          5793 => x"04",
          5794 => x"04",
          5795 => x"04",
          5796 => x"04",
          5797 => x"04",
          5798 => x"04",
          5799 => x"04",
          5800 => x"04",
          5801 => x"04",
          5802 => x"04",
          5803 => x"04",
          5804 => x"04",
          5805 => x"04",
          5806 => x"04",
          5807 => x"04",
          5808 => x"04",
          5809 => x"04",
          5810 => x"04",
          5811 => x"04",
          5812 => x"04",
          5813 => x"04",
          5814 => x"04",
          5815 => x"04",
          5816 => x"04",
          5817 => x"04",
          5818 => x"04",
          5819 => x"04",
          5820 => x"04",
          5821 => x"04",
          5822 => x"04",
          5823 => x"04",
          5824 => x"04",
          5825 => x"04",
          5826 => x"04",
          5827 => x"04",
          5828 => x"04",
          5829 => x"04",
          5830 => x"04",
          5831 => x"04",
          5832 => x"04",
          5833 => x"04",
          5834 => x"64",
          5835 => x"2f",
          5836 => x"25",
          5837 => x"64",
          5838 => x"2e",
          5839 => x"64",
          5840 => x"6f",
          5841 => x"6f",
          5842 => x"67",
          5843 => x"74",
          5844 => x"00",
          5845 => x"28",
          5846 => x"6d",
          5847 => x"43",
          5848 => x"6e",
          5849 => x"29",
          5850 => x"0a",
          5851 => x"69",
          5852 => x"20",
          5853 => x"6c",
          5854 => x"6e",
          5855 => x"3a",
          5856 => x"20",
          5857 => x"4e",
          5858 => x"42",
          5859 => x"20",
          5860 => x"61",
          5861 => x"25",
          5862 => x"2c",
          5863 => x"7a",
          5864 => x"30",
          5865 => x"2e",
          5866 => x"20",
          5867 => x"52",
          5868 => x"28",
          5869 => x"72",
          5870 => x"30",
          5871 => x"20",
          5872 => x"65",
          5873 => x"38",
          5874 => x"0a",
          5875 => x"20",
          5876 => x"41",
          5877 => x"53",
          5878 => x"74",
          5879 => x"38",
          5880 => x"53",
          5881 => x"3d",
          5882 => x"58",
          5883 => x"00",
          5884 => x"20",
          5885 => x"4f",
          5886 => x"0a",
          5887 => x"20",
          5888 => x"53",
          5889 => x"00",
          5890 => x"20",
          5891 => x"50",
          5892 => x"00",
          5893 => x"20",
          5894 => x"44",
          5895 => x"72",
          5896 => x"44",
          5897 => x"63",
          5898 => x"25",
          5899 => x"29",
          5900 => x"00",
          5901 => x"20",
          5902 => x"4e",
          5903 => x"52",
          5904 => x"20",
          5905 => x"54",
          5906 => x"4c",
          5907 => x"00",
          5908 => x"20",
          5909 => x"49",
          5910 => x"31",
          5911 => x"69",
          5912 => x"73",
          5913 => x"31",
          5914 => x"0a",
          5915 => x"64",
          5916 => x"73",
          5917 => x"3a",
          5918 => x"20",
          5919 => x"50",
          5920 => x"65",
          5921 => x"20",
          5922 => x"74",
          5923 => x"41",
          5924 => x"65",
          5925 => x"3d",
          5926 => x"38",
          5927 => x"00",
          5928 => x"20",
          5929 => x"50",
          5930 => x"65",
          5931 => x"79",
          5932 => x"61",
          5933 => x"41",
          5934 => x"65",
          5935 => x"3d",
          5936 => x"38",
          5937 => x"00",
          5938 => x"20",
          5939 => x"74",
          5940 => x"20",
          5941 => x"72",
          5942 => x"64",
          5943 => x"73",
          5944 => x"20",
          5945 => x"3d",
          5946 => x"38",
          5947 => x"00",
          5948 => x"20",
          5949 => x"50",
          5950 => x"64",
          5951 => x"20",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"3d",
          5956 => x"38",
          5957 => x"00",
          5958 => x"20",
          5959 => x"79",
          5960 => x"6d",
          5961 => x"6f",
          5962 => x"46",
          5963 => x"20",
          5964 => x"20",
          5965 => x"3d",
          5966 => x"38",
          5967 => x"00",
          5968 => x"6d",
          5969 => x"00",
          5970 => x"65",
          5971 => x"6d",
          5972 => x"6c",
          5973 => x"00",
          5974 => x"56",
          5975 => x"56",
          5976 => x"6e",
          5977 => x"6e",
          5978 => x"77",
          5979 => x"44",
          5980 => x"2a",
          5981 => x"3b",
          5982 => x"3f",
          5983 => x"7f",
          5984 => x"41",
          5985 => x"41",
          5986 => x"00",
          5987 => x"0a",
          5988 => x"0a",
          5989 => x"0a",
          5990 => x"0a",
          5991 => x"0a",
          5992 => x"0a",
          5993 => x"0a",
          5994 => x"0a",
          5995 => x"0a",
          5996 => x"30",
          5997 => x"fe",
          5998 => x"44",
          5999 => x"2e",
          6000 => x"4f",
          6001 => x"4d",
          6002 => x"20",
          6003 => x"54",
          6004 => x"20",
          6005 => x"4f",
          6006 => x"4d",
          6007 => x"20",
          6008 => x"54",
          6009 => x"20",
          6010 => x"04",
          6011 => x"00",
          6012 => x"00",
          6013 => x"00",
          6014 => x"9a",
          6015 => x"41",
          6016 => x"45",
          6017 => x"49",
          6018 => x"92",
          6019 => x"4f",
          6020 => x"99",
          6021 => x"9d",
          6022 => x"49",
          6023 => x"a5",
          6024 => x"a9",
          6025 => x"ad",
          6026 => x"b1",
          6027 => x"b5",
          6028 => x"b9",
          6029 => x"bd",
          6030 => x"c1",
          6031 => x"c5",
          6032 => x"c9",
          6033 => x"cd",
          6034 => x"d1",
          6035 => x"d5",
          6036 => x"d9",
          6037 => x"dd",
          6038 => x"e1",
          6039 => x"e5",
          6040 => x"e9",
          6041 => x"ed",
          6042 => x"f1",
          6043 => x"f5",
          6044 => x"f9",
          6045 => x"fd",
          6046 => x"2e",
          6047 => x"5b",
          6048 => x"22",
          6049 => x"3e",
          6050 => x"00",
          6051 => x"01",
          6052 => x"10",
          6053 => x"00",
          6054 => x"00",
          6055 => x"01",
          6056 => x"04",
          6057 => x"10",
          6058 => x"00",
          6059 => x"41",
          6060 => x"00",
          6061 => x"41",
          6062 => x"00",
          6063 => x"78",
          6064 => x"00",
          6065 => x"49",
          6066 => x"49",
          6067 => x"4f",
          6068 => x"4f",
          6069 => x"00",
          6070 => x"49",
          6071 => x"42",
          6072 => x"45",
          6073 => x"4f",
          6074 => x"4f",
          6075 => x"00",
          6076 => x"49",
          6077 => x"59",
          6078 => x"4d",
          6079 => x"4e",
          6080 => x"4c",
          6081 => x"45",
          6082 => x"59",
          6083 => x"41",
          6084 => x"41",
          6085 => x"00",
          6086 => x"45",
          6087 => x"4e",
          6088 => x"58",
          6089 => x"54",
          6090 => x"00",
          6091 => x"49",
          6092 => x"43",
          6093 => x"41",
          6094 => x"00",
          6095 => x"64",
          6096 => x"00",
          6097 => x"69",
          6098 => x"00",
          6099 => x"73",
          6100 => x"00",
          6101 => x"69",
          6102 => x"6c",
          6103 => x"64",
          6104 => x"00",
          6105 => x"65",
          6106 => x"00",
          6107 => x"72",
          6108 => x"00",
          6109 => x"77",
          6110 => x"65",
          6111 => x"66",
          6112 => x"00",
          6113 => x"6c",
          6114 => x"00",
          6115 => x"69",
          6116 => x"00",
          6117 => x"6f",
          6118 => x"00",
          6119 => x"63",
          6120 => x"65",
          6121 => x"73",
          6122 => x"00",
          6123 => x"72",
          6124 => x"00",
          6125 => x"69",
          6126 => x"65",
          6127 => x"00",
          6128 => x"77",
          6129 => x"65",
          6130 => x"74",
          6131 => x"63",
          6132 => x"61",
          6133 => x"63",
          6134 => x"61",
          6135 => x"00",
          6136 => x"74",
          6137 => x"00",
          6138 => x"72",
          6139 => x"6d",
          6140 => x"64",
          6141 => x"00",
          6142 => x"6d",
          6143 => x"72",
          6144 => x"73",
          6145 => x"00",
          6146 => x"64",
          6147 => x"00",
          6148 => x"63",
          6149 => x"00",
          6150 => x"63",
          6151 => x"63",
          6152 => x"61",
          6153 => x"78",
          6154 => x"63",
          6155 => x"6c",
          6156 => x"00",
          6157 => x"65",
          6158 => x"00",
          6159 => x"73",
          6160 => x"00",
          6161 => x"64",
          6162 => x"00",
          6163 => x"63",
          6164 => x"64",
          6165 => x"65",
          6166 => x"73",
          6167 => x"64",
          6168 => x"00",
          6169 => x"6c",
          6170 => x"6c",
          6171 => x"6d",
          6172 => x"00",
          6173 => x"63",
          6174 => x"00",
          6175 => x"64",
          6176 => x"00",
          6177 => x"65",
          6178 => x"65",
          6179 => x"65",
          6180 => x"69",
          6181 => x"69",
          6182 => x"72",
          6183 => x"74",
          6184 => x"66",
          6185 => x"66",
          6186 => x"68",
          6187 => x"00",
          6188 => x"6f",
          6189 => x"61",
          6190 => x"00",
          6191 => x"61",
          6192 => x"00",
          6193 => x"6d",
          6194 => x"65",
          6195 => x"72",
          6196 => x"65",
          6197 => x"00",
          6198 => x"65",
          6199 => x"00",
          6200 => x"6e",
          6201 => x"00",
          6202 => x"69",
          6203 => x"00",
          6204 => x"65",
          6205 => x"00",
          6206 => x"69",
          6207 => x"45",
          6208 => x"72",
          6209 => x"6e",
          6210 => x"6e",
          6211 => x"65",
          6212 => x"72",
          6213 => x"00",
          6214 => x"69",
          6215 => x"6e",
          6216 => x"72",
          6217 => x"79",
          6218 => x"00",
          6219 => x"6f",
          6220 => x"6c",
          6221 => x"6f",
          6222 => x"2e",
          6223 => x"6f",
          6224 => x"74",
          6225 => x"6f",
          6226 => x"2e",
          6227 => x"6e",
          6228 => x"69",
          6229 => x"69",
          6230 => x"61",
          6231 => x"0a",
          6232 => x"63",
          6233 => x"73",
          6234 => x"6e",
          6235 => x"2e",
          6236 => x"69",
          6237 => x"61",
          6238 => x"61",
          6239 => x"65",
          6240 => x"74",
          6241 => x"00",
          6242 => x"69",
          6243 => x"68",
          6244 => x"6c",
          6245 => x"6e",
          6246 => x"69",
          6247 => x"00",
          6248 => x"44",
          6249 => x"20",
          6250 => x"74",
          6251 => x"72",
          6252 => x"63",
          6253 => x"2e",
          6254 => x"72",
          6255 => x"20",
          6256 => x"62",
          6257 => x"69",
          6258 => x"6e",
          6259 => x"69",
          6260 => x"00",
          6261 => x"69",
          6262 => x"6e",
          6263 => x"65",
          6264 => x"6c",
          6265 => x"0a",
          6266 => x"6f",
          6267 => x"6d",
          6268 => x"69",
          6269 => x"20",
          6270 => x"65",
          6271 => x"74",
          6272 => x"66",
          6273 => x"64",
          6274 => x"20",
          6275 => x"6b",
          6276 => x"00",
          6277 => x"6f",
          6278 => x"74",
          6279 => x"6f",
          6280 => x"64",
          6281 => x"00",
          6282 => x"69",
          6283 => x"75",
          6284 => x"6f",
          6285 => x"61",
          6286 => x"6e",
          6287 => x"6e",
          6288 => x"6c",
          6289 => x"0a",
          6290 => x"69",
          6291 => x"69",
          6292 => x"6f",
          6293 => x"64",
          6294 => x"00",
          6295 => x"6e",
          6296 => x"66",
          6297 => x"65",
          6298 => x"6d",
          6299 => x"72",
          6300 => x"00",
          6301 => x"6f",
          6302 => x"61",
          6303 => x"6f",
          6304 => x"20",
          6305 => x"65",
          6306 => x"00",
          6307 => x"61",
          6308 => x"65",
          6309 => x"73",
          6310 => x"63",
          6311 => x"65",
          6312 => x"0a",
          6313 => x"75",
          6314 => x"73",
          6315 => x"00",
          6316 => x"6e",
          6317 => x"77",
          6318 => x"72",
          6319 => x"2e",
          6320 => x"25",
          6321 => x"62",
          6322 => x"73",
          6323 => x"20",
          6324 => x"25",
          6325 => x"62",
          6326 => x"73",
          6327 => x"63",
          6328 => x"00",
          6329 => x"65",
          6330 => x"00",
          6331 => x"50",
          6332 => x"00",
          6333 => x"2a",
          6334 => x"73",
          6335 => x"00",
          6336 => x"38",
          6337 => x"2f",
          6338 => x"39",
          6339 => x"31",
          6340 => x"00",
          6341 => x"5a",
          6342 => x"20",
          6343 => x"20",
          6344 => x"78",
          6345 => x"73",
          6346 => x"20",
          6347 => x"0a",
          6348 => x"50",
          6349 => x"20",
          6350 => x"65",
          6351 => x"70",
          6352 => x"61",
          6353 => x"65",
          6354 => x"00",
          6355 => x"69",
          6356 => x"20",
          6357 => x"65",
          6358 => x"70",
          6359 => x"00",
          6360 => x"53",
          6361 => x"6e",
          6362 => x"72",
          6363 => x"0a",
          6364 => x"4f",
          6365 => x"20",
          6366 => x"69",
          6367 => x"72",
          6368 => x"74",
          6369 => x"4f",
          6370 => x"20",
          6371 => x"69",
          6372 => x"72",
          6373 => x"74",
          6374 => x"41",
          6375 => x"20",
          6376 => x"69",
          6377 => x"72",
          6378 => x"74",
          6379 => x"41",
          6380 => x"20",
          6381 => x"69",
          6382 => x"72",
          6383 => x"74",
          6384 => x"41",
          6385 => x"20",
          6386 => x"69",
          6387 => x"72",
          6388 => x"74",
          6389 => x"41",
          6390 => x"20",
          6391 => x"69",
          6392 => x"72",
          6393 => x"74",
          6394 => x"65",
          6395 => x"6e",
          6396 => x"70",
          6397 => x"6d",
          6398 => x"2e",
          6399 => x"00",
          6400 => x"6e",
          6401 => x"69",
          6402 => x"74",
          6403 => x"72",
          6404 => x"0a",
          6405 => x"3a",
          6406 => x"61",
          6407 => x"64",
          6408 => x"20",
          6409 => x"74",
          6410 => x"69",
          6411 => x"73",
          6412 => x"61",
          6413 => x"30",
          6414 => x"6c",
          6415 => x"65",
          6416 => x"69",
          6417 => x"61",
          6418 => x"6c",
          6419 => x"0a",
          6420 => x"20",
          6421 => x"61",
          6422 => x"69",
          6423 => x"69",
          6424 => x"00",
          6425 => x"6e",
          6426 => x"61",
          6427 => x"65",
          6428 => x"00",
          6429 => x"61",
          6430 => x"64",
          6431 => x"20",
          6432 => x"74",
          6433 => x"69",
          6434 => x"0a",
          6435 => x"63",
          6436 => x"0a",
          6437 => x"75",
          6438 => x"69",
          6439 => x"6c",
          6440 => x"20",
          6441 => x"65",
          6442 => x"70",
          6443 => x"00",
          6444 => x"6e",
          6445 => x"69",
          6446 => x"69",
          6447 => x"72",
          6448 => x"74",
          6449 => x"00",
          6450 => x"69",
          6451 => x"6c",
          6452 => x"75",
          6453 => x"20",
          6454 => x"6f",
          6455 => x"6e",
          6456 => x"69",
          6457 => x"75",
          6458 => x"20",
          6459 => x"6f",
          6460 => x"78",
          6461 => x"74",
          6462 => x"20",
          6463 => x"65",
          6464 => x"25",
          6465 => x"20",
          6466 => x"0a",
          6467 => x"61",
          6468 => x"6e",
          6469 => x"6f",
          6470 => x"40",
          6471 => x"38",
          6472 => x"2e",
          6473 => x"00",
          6474 => x"61",
          6475 => x"72",
          6476 => x"72",
          6477 => x"20",
          6478 => x"65",
          6479 => x"64",
          6480 => x"00",
          6481 => x"65",
          6482 => x"72",
          6483 => x"67",
          6484 => x"70",
          6485 => x"61",
          6486 => x"6e",
          6487 => x"0a",
          6488 => x"6f",
          6489 => x"72",
          6490 => x"6f",
          6491 => x"67",
          6492 => x"0a",
          6493 => x"50",
          6494 => x"69",
          6495 => x"64",
          6496 => x"73",
          6497 => x"2e",
          6498 => x"00",
          6499 => x"61",
          6500 => x"6f",
          6501 => x"6e",
          6502 => x"00",
          6503 => x"75",
          6504 => x"6e",
          6505 => x"2e",
          6506 => x"6e",
          6507 => x"69",
          6508 => x"69",
          6509 => x"72",
          6510 => x"74",
          6511 => x"2e",
          6512 => x"00",
          6513 => x"00",
          6514 => x"00",
          6515 => x"00",
          6516 => x"00",
          6517 => x"01",
          6518 => x"00",
          6519 => x"00",
          6520 => x"00",
          6521 => x"00",
          6522 => x"00",
          6523 => x"f5",
          6524 => x"01",
          6525 => x"01",
          6526 => x"01",
          6527 => x"00",
          6528 => x"00",
          6529 => x"00",
          6530 => x"04",
          6531 => x"01",
          6532 => x"00",
          6533 => x"00",
          6534 => x"04",
          6535 => x"02",
          6536 => x"00",
          6537 => x"00",
          6538 => x"04",
          6539 => x"03",
          6540 => x"00",
          6541 => x"00",
          6542 => x"04",
          6543 => x"04",
          6544 => x"00",
          6545 => x"00",
          6546 => x"04",
          6547 => x"0a",
          6548 => x"00",
          6549 => x"00",
          6550 => x"04",
          6551 => x"0b",
          6552 => x"00",
          6553 => x"00",
          6554 => x"04",
          6555 => x"0c",
          6556 => x"00",
          6557 => x"00",
          6558 => x"04",
          6559 => x"0d",
          6560 => x"00",
          6561 => x"00",
          6562 => x"04",
          6563 => x"0e",
          6564 => x"00",
          6565 => x"00",
          6566 => x"04",
          6567 => x"0f",
          6568 => x"00",
          6569 => x"00",
          6570 => x"04",
          6571 => x"14",
          6572 => x"00",
          6573 => x"00",
          6574 => x"04",
          6575 => x"17",
          6576 => x"00",
          6577 => x"00",
          6578 => x"04",
          6579 => x"18",
          6580 => x"00",
          6581 => x"00",
          6582 => x"04",
          6583 => x"19",
          6584 => x"00",
          6585 => x"00",
          6586 => x"04",
          6587 => x"1a",
          6588 => x"00",
          6589 => x"00",
          6590 => x"04",
          6591 => x"1c",
          6592 => x"00",
          6593 => x"00",
          6594 => x"04",
          6595 => x"1d",
          6596 => x"00",
          6597 => x"00",
          6598 => x"04",
          6599 => x"1e",
          6600 => x"00",
          6601 => x"00",
          6602 => x"04",
          6603 => x"22",
          6604 => x"00",
          6605 => x"00",
          6606 => x"04",
          6607 => x"23",
          6608 => x"00",
          6609 => x"00",
          6610 => x"04",
          6611 => x"24",
          6612 => x"00",
          6613 => x"00",
          6614 => x"04",
          6615 => x"1f",
          6616 => x"00",
          6617 => x"00",
          6618 => x"04",
          6619 => x"20",
          6620 => x"00",
          6621 => x"00",
          6622 => x"04",
          6623 => x"21",
          6624 => x"00",
          6625 => x"00",
          6626 => x"04",
          6627 => x"15",
          6628 => x"00",
          6629 => x"00",
          6630 => x"04",
          6631 => x"16",
          6632 => x"00",
          6633 => x"00",
          6634 => x"04",
          6635 => x"1b",
          6636 => x"00",
          6637 => x"00",
          6638 => x"04",
          6639 => x"25",
          6640 => x"00",
          6641 => x"00",
          6642 => x"04",
          6643 => x"2d",
          6644 => x"00",
          6645 => x"00",
          6646 => x"04",
          6647 => x"2e",
          6648 => x"00",
          6649 => x"00",
          6650 => x"04",
          6651 => x"2b",
          6652 => x"00",
          6653 => x"00",
          6654 => x"04",
          6655 => x"30",
          6656 => x"00",
          6657 => x"00",
          6658 => x"04",
          6659 => x"2f",
          6660 => x"00",
          6661 => x"00",
          6662 => x"04",
          6663 => x"2c",
          6664 => x"00",
          6665 => x"00",
          6666 => x"04",
          6667 => x"26",
          6668 => x"00",
          6669 => x"00",
          6670 => x"04",
          6671 => x"27",
          6672 => x"00",
          6673 => x"00",
          6674 => x"04",
          6675 => x"28",
          6676 => x"00",
          6677 => x"00",
          6678 => x"04",
          6679 => x"29",
          6680 => x"00",
          6681 => x"00",
          6682 => x"04",
          6683 => x"2a",
          6684 => x"00",
          6685 => x"00",
          6686 => x"04",
          6687 => x"3c",
          6688 => x"00",
          6689 => x"00",
          6690 => x"04",
          6691 => x"3d",
          6692 => x"00",
          6693 => x"00",
          6694 => x"04",
          6695 => x"3e",
          6696 => x"00",
          6697 => x"00",
          6698 => x"04",
          6699 => x"3f",
          6700 => x"00",
          6701 => x"00",
          6702 => x"04",
          6703 => x"40",
          6704 => x"00",
          6705 => x"00",
          6706 => x"04",
          6707 => x"50",
          6708 => x"00",
          6709 => x"00",
          6710 => x"04",
          6711 => x"51",
          6712 => x"00",
          6713 => x"00",
          6714 => x"04",
          6715 => x"52",
          6716 => x"00",
          6717 => x"00",
          6718 => x"04",
          6719 => x"53",
          6720 => x"00",
          6721 => x"00",
          6722 => x"04",
          6723 => x"54",
          6724 => x"00",
          6725 => x"00",
          6726 => x"04",
          6727 => x"55",
          6728 => x"00",
          6729 => x"00",
          6730 => x"04",
          6731 => x"64",
          6732 => x"00",
          6733 => x"00",
          6734 => x"04",
          6735 => x"65",
          6736 => x"00",
          6737 => x"00",
          6738 => x"04",
          6739 => x"79",
          6740 => x"00",
          6741 => x"00",
          6742 => x"04",
          6743 => x"78",
          6744 => x"00",
          6745 => x"00",
          6746 => x"04",
          6747 => x"82",
          6748 => x"00",
          6749 => x"00",
          6750 => x"04",
          6751 => x"83",
          6752 => x"00",
          6753 => x"00",
          6754 => x"04",
          6755 => x"84",
          6756 => x"00",
          6757 => x"00",
          6758 => x"04",
          6759 => x"85",
          6760 => x"00",
          6761 => x"00",
          6762 => x"04",
          6763 => x"86",
          6764 => x"00",
          6765 => x"00",
          6766 => x"04",
          6767 => x"87",
          6768 => x"00",
          6769 => x"00",
        others => X"00"
    );

    shared variable RAM3 : ramArray :=
    (
             0 => x"0b",
             1 => x"80",
             2 => x"90",
             3 => x"ff",
             4 => x"ff",
             5 => x"ff",
             6 => x"ff",
             7 => x"ff",
             8 => x"0b",
             9 => x"80",
            10 => x"90",
            11 => x"0b",
            12 => x"95",
            13 => x"90",
            14 => x"0b",
            15 => x"b5",
            16 => x"90",
            17 => x"0b",
            18 => x"d5",
            19 => x"90",
            20 => x"0b",
            21 => x"f5",
            22 => x"90",
            23 => x"0b",
            24 => x"95",
            25 => x"90",
            26 => x"0b",
            27 => x"b5",
            28 => x"90",
            29 => x"0b",
            30 => x"d5",
            31 => x"90",
            32 => x"0b",
            33 => x"f5",
            34 => x"90",
            35 => x"0b",
            36 => x"95",
            37 => x"90",
            38 => x"0b",
            39 => x"b5",
            40 => x"90",
            41 => x"0b",
            42 => x"d5",
            43 => x"90",
            44 => x"0b",
            45 => x"f5",
            46 => x"90",
            47 => x"0b",
            48 => x"95",
            49 => x"90",
            50 => x"0b",
            51 => x"b5",
            52 => x"90",
            53 => x"0b",
            54 => x"d5",
            55 => x"90",
            56 => x"0b",
            57 => x"f5",
            58 => x"90",
            59 => x"0b",
            60 => x"95",
            61 => x"90",
            62 => x"0b",
            63 => x"b5",
            64 => x"90",
            65 => x"0b",
            66 => x"d5",
            67 => x"90",
            68 => x"0b",
            69 => x"f5",
            70 => x"90",
            71 => x"0b",
            72 => x"95",
            73 => x"90",
            74 => x"0b",
            75 => x"b5",
            76 => x"90",
            77 => x"0b",
            78 => x"d5",
            79 => x"90",
            80 => x"0b",
            81 => x"f5",
            82 => x"90",
            83 => x"00",
            84 => x"00",
            85 => x"00",
            86 => x"00",
            87 => x"00",
            88 => x"00",
            89 => x"00",
            90 => x"00",
            91 => x"00",
            92 => x"00",
            93 => x"00",
            94 => x"00",
            95 => x"00",
            96 => x"00",
            97 => x"00",
            98 => x"00",
            99 => x"00",
           100 => x"00",
           101 => x"00",
           102 => x"00",
           103 => x"00",
           104 => x"00",
           105 => x"00",
           106 => x"00",
           107 => x"00",
           108 => x"00",
           109 => x"00",
           110 => x"00",
           111 => x"00",
           112 => x"00",
           113 => x"00",
           114 => x"00",
           115 => x"00",
           116 => x"00",
           117 => x"00",
           118 => x"00",
           119 => x"00",
           120 => x"00",
           121 => x"00",
           122 => x"00",
           123 => x"00",
           124 => x"00",
           125 => x"00",
           126 => x"00",
           127 => x"00",
           128 => x"00",
           129 => x"04",
           130 => x"0c",
           131 => x"2d",
           132 => x"08",
           133 => x"04",
           134 => x"0c",
           135 => x"2d",
           136 => x"08",
           137 => x"04",
           138 => x"0c",
           139 => x"2d",
           140 => x"08",
           141 => x"04",
           142 => x"0c",
           143 => x"2d",
           144 => x"08",
           145 => x"04",
           146 => x"0c",
           147 => x"2d",
           148 => x"08",
           149 => x"04",
           150 => x"0c",
           151 => x"2d",
           152 => x"08",
           153 => x"04",
           154 => x"0c",
           155 => x"2d",
           156 => x"08",
           157 => x"04",
           158 => x"0c",
           159 => x"2d",
           160 => x"08",
           161 => x"04",
           162 => x"0c",
           163 => x"2d",
           164 => x"08",
           165 => x"04",
           166 => x"0c",
           167 => x"2d",
           168 => x"08",
           169 => x"04",
           170 => x"0c",
           171 => x"2d",
           172 => x"08",
           173 => x"04",
           174 => x"0c",
           175 => x"2d",
           176 => x"08",
           177 => x"04",
           178 => x"0c",
           179 => x"2d",
           180 => x"08",
           181 => x"04",
           182 => x"0c",
           183 => x"2d",
           184 => x"08",
           185 => x"04",
           186 => x"0c",
           187 => x"2d",
           188 => x"08",
           189 => x"04",
           190 => x"0c",
           191 => x"2d",
           192 => x"08",
           193 => x"04",
           194 => x"0c",
           195 => x"2d",
           196 => x"08",
           197 => x"04",
           198 => x"0c",
           199 => x"2d",
           200 => x"08",
           201 => x"04",
           202 => x"0c",
           203 => x"2d",
           204 => x"08",
           205 => x"04",
           206 => x"0c",
           207 => x"2d",
           208 => x"08",
           209 => x"04",
           210 => x"0c",
           211 => x"2d",
           212 => x"08",
           213 => x"04",
           214 => x"0c",
           215 => x"2d",
           216 => x"08",
           217 => x"04",
           218 => x"0c",
           219 => x"2d",
           220 => x"08",
           221 => x"04",
           222 => x"0c",
           223 => x"2d",
           224 => x"08",
           225 => x"04",
           226 => x"0c",
           227 => x"2d",
           228 => x"08",
           229 => x"04",
           230 => x"0c",
           231 => x"2d",
           232 => x"08",
           233 => x"04",
           234 => x"0c",
           235 => x"2d",
           236 => x"08",
           237 => x"04",
           238 => x"0c",
           239 => x"2d",
           240 => x"08",
           241 => x"04",
           242 => x"0c",
           243 => x"2d",
           244 => x"08",
           245 => x"04",
           246 => x"0c",
           247 => x"2d",
           248 => x"08",
           249 => x"04",
           250 => x"0c",
           251 => x"2d",
           252 => x"08",
           253 => x"04",
           254 => x"0c",
           255 => x"2d",
           256 => x"08",
           257 => x"04",
           258 => x"0c",
           259 => x"2d",
           260 => x"08",
           261 => x"04",
           262 => x"0c",
           263 => x"2d",
           264 => x"08",
           265 => x"04",
           266 => x"0c",
           267 => x"2d",
           268 => x"08",
           269 => x"04",
           270 => x"0c",
           271 => x"2d",
           272 => x"08",
           273 => x"04",
           274 => x"0c",
           275 => x"2d",
           276 => x"08",
           277 => x"04",
           278 => x"0c",
           279 => x"2d",
           280 => x"08",
           281 => x"04",
           282 => x"0c",
           283 => x"2d",
           284 => x"08",
           285 => x"04",
           286 => x"0c",
           287 => x"2d",
           288 => x"08",
           289 => x"04",
           290 => x"0c",
           291 => x"2d",
           292 => x"08",
           293 => x"04",
           294 => x"0c",
           295 => x"2d",
           296 => x"08",
           297 => x"04",
           298 => x"0c",
           299 => x"2d",
           300 => x"08",
           301 => x"04",
           302 => x"0c",
           303 => x"2d",
           304 => x"08",
           305 => x"04",
           306 => x"0c",
           307 => x"2d",
           308 => x"08",
           309 => x"04",
           310 => x"0c",
           311 => x"2d",
           312 => x"08",
           313 => x"04",
           314 => x"0c",
           315 => x"2d",
           316 => x"08",
           317 => x"04",
           318 => x"0c",
           319 => x"2d",
           320 => x"08",
           321 => x"04",
           322 => x"0c",
           323 => x"2d",
           324 => x"08",
           325 => x"04",
           326 => x"70",
           327 => x"27",
           328 => x"71",
           329 => x"53",
           330 => x"90",
           331 => x"90",
           332 => x"91",
           333 => x"3c",
           334 => x"d4",
           335 => x"d3",
           336 => x"3d",
           337 => x"91",
           338 => x"8c",
           339 => x"91",
           340 => x"88",
           341 => x"80",
           342 => x"d3",
           343 => x"91",
           344 => x"54",
           345 => x"91",
           346 => x"04",
           347 => x"08",
           348 => x"d4",
           349 => x"0d",
           350 => x"d3",
           351 => x"05",
           352 => x"d3",
           353 => x"05",
           354 => x"3f",
           355 => x"08",
           356 => x"c8",
           357 => x"3d",
           358 => x"d4",
           359 => x"d3",
           360 => x"91",
           361 => x"fd",
           362 => x"0b",
           363 => x"08",
           364 => x"80",
           365 => x"d4",
           366 => x"0c",
           367 => x"08",
           368 => x"91",
           369 => x"88",
           370 => x"b9",
           371 => x"d4",
           372 => x"08",
           373 => x"38",
           374 => x"d3",
           375 => x"05",
           376 => x"38",
           377 => x"08",
           378 => x"10",
           379 => x"08",
           380 => x"91",
           381 => x"fc",
           382 => x"91",
           383 => x"fc",
           384 => x"b8",
           385 => x"d4",
           386 => x"08",
           387 => x"e1",
           388 => x"d4",
           389 => x"08",
           390 => x"08",
           391 => x"26",
           392 => x"d3",
           393 => x"05",
           394 => x"d4",
           395 => x"08",
           396 => x"d4",
           397 => x"0c",
           398 => x"08",
           399 => x"91",
           400 => x"fc",
           401 => x"91",
           402 => x"f8",
           403 => x"d3",
           404 => x"05",
           405 => x"91",
           406 => x"fc",
           407 => x"d3",
           408 => x"05",
           409 => x"91",
           410 => x"8c",
           411 => x"95",
           412 => x"d4",
           413 => x"08",
           414 => x"38",
           415 => x"08",
           416 => x"70",
           417 => x"08",
           418 => x"51",
           419 => x"d3",
           420 => x"05",
           421 => x"d3",
           422 => x"05",
           423 => x"d3",
           424 => x"05",
           425 => x"c8",
           426 => x"0d",
           427 => x"0c",
           428 => x"0d",
           429 => x"02",
           430 => x"05",
           431 => x"53",
           432 => x"27",
           433 => x"83",
           434 => x"80",
           435 => x"ff",
           436 => x"ff",
           437 => x"73",
           438 => x"05",
           439 => x"12",
           440 => x"2e",
           441 => x"ef",
           442 => x"d3",
           443 => x"3d",
           444 => x"74",
           445 => x"07",
           446 => x"2b",
           447 => x"51",
           448 => x"a5",
           449 => x"70",
           450 => x"0c",
           451 => x"84",
           452 => x"72",
           453 => x"05",
           454 => x"71",
           455 => x"53",
           456 => x"52",
           457 => x"dd",
           458 => x"27",
           459 => x"71",
           460 => x"53",
           461 => x"52",
           462 => x"f2",
           463 => x"ff",
           464 => x"3d",
           465 => x"70",
           466 => x"06",
           467 => x"70",
           468 => x"73",
           469 => x"56",
           470 => x"08",
           471 => x"38",
           472 => x"52",
           473 => x"81",
           474 => x"54",
           475 => x"9d",
           476 => x"55",
           477 => x"09",
           478 => x"38",
           479 => x"14",
           480 => x"81",
           481 => x"56",
           482 => x"e5",
           483 => x"55",
           484 => x"06",
           485 => x"06",
           486 => x"91",
           487 => x"52",
           488 => x"0d",
           489 => x"70",
           490 => x"ff",
           491 => x"f8",
           492 => x"80",
           493 => x"51",
           494 => x"84",
           495 => x"71",
           496 => x"54",
           497 => x"2e",
           498 => x"75",
           499 => x"94",
           500 => x"91",
           501 => x"87",
           502 => x"fe",
           503 => x"70",
           504 => x"88",
           505 => x"9b",
           506 => x"c8",
           507 => x"06",
           508 => x"14",
           509 => x"73",
           510 => x"71",
           511 => x"0c",
           512 => x"04",
           513 => x"76",
           514 => x"53",
           515 => x"80",
           516 => x"38",
           517 => x"70",
           518 => x"81",
           519 => x"81",
           520 => x"52",
           521 => x"2e",
           522 => x"52",
           523 => x"12",
           524 => x"33",
           525 => x"a0",
           526 => x"81",
           527 => x"70",
           528 => x"06",
           529 => x"e6",
           530 => x"51",
           531 => x"09",
           532 => x"38",
           533 => x"81",
           534 => x"71",
           535 => x"51",
           536 => x"c8",
           537 => x"0d",
           538 => x"0d",
           539 => x"08",
           540 => x"38",
           541 => x"05",
           542 => x"99",
           543 => x"d3",
           544 => x"38",
           545 => x"39",
           546 => x"91",
           547 => x"86",
           548 => x"f5",
           549 => x"82",
           550 => x"05",
           551 => x"5b",
           552 => x"81",
           553 => x"1c",
           554 => x"5a",
           555 => x"9e",
           556 => x"38",
           557 => x"5a",
           558 => x"97",
           559 => x"38",
           560 => x"5a",
           561 => x"bb",
           562 => x"38",
           563 => x"5a",
           564 => x"bb",
           565 => x"38",
           566 => x"5a",
           567 => x"87",
           568 => x"80",
           569 => x"22",
           570 => x"79",
           571 => x"80",
           572 => x"1c",
           573 => x"1c",
           574 => x"1c",
           575 => x"1c",
           576 => x"1c",
           577 => x"1c",
           578 => x"1c",
           579 => x"22",
           580 => x"a8",
           581 => x"3f",
           582 => x"9c",
           583 => x"0c",
           584 => x"c0",
           585 => x"82",
           586 => x"c0",
           587 => x"83",
           588 => x"c0",
           589 => x"84",
           590 => x"c0",
           591 => x"85",
           592 => x"c0",
           593 => x"86",
           594 => x"c0",
           595 => x"88",
           596 => x"c0",
           597 => x"8a",
           598 => x"c0",
           599 => x"80",
           600 => x"5b",
           601 => x"c8",
           602 => x"0d",
           603 => x"0d",
           604 => x"c0",
           605 => x"81",
           606 => x"c0",
           607 => x"5b",
           608 => x"87",
           609 => x"08",
           610 => x"1b",
           611 => x"98",
           612 => x"7a",
           613 => x"87",
           614 => x"08",
           615 => x"1b",
           616 => x"98",
           617 => x"7a",
           618 => x"87",
           619 => x"08",
           620 => x"1b",
           621 => x"98",
           622 => x"7a",
           623 => x"87",
           624 => x"08",
           625 => x"1b",
           626 => x"0c",
           627 => x"59",
           628 => x"58",
           629 => x"57",
           630 => x"56",
           631 => x"55",
           632 => x"54",
           633 => x"53",
           634 => x"91",
           635 => x"92",
           636 => x"3d",
           637 => x"3d",
           638 => x"05",
           639 => x"70",
           640 => x"51",
           641 => x"0b",
           642 => x"34",
           643 => x"04",
           644 => x"75",
           645 => x"cb",
           646 => x"54",
           647 => x"84",
           648 => x"2e",
           649 => x"c0",
           650 => x"70",
           651 => x"2a",
           652 => x"51",
           653 => x"80",
           654 => x"71",
           655 => x"81",
           656 => x"70",
           657 => x"96",
           658 => x"70",
           659 => x"51",
           660 => x"8d",
           661 => x"2a",
           662 => x"51",
           663 => x"bc",
           664 => x"91",
           665 => x"51",
           666 => x"80",
           667 => x"2e",
           668 => x"c0",
           669 => x"73",
           670 => x"91",
           671 => x"85",
           672 => x"fd",
           673 => x"97",
           674 => x"0b",
           675 => x"33",
           676 => x"c0",
           677 => x"72",
           678 => x"38",
           679 => x"94",
           680 => x"70",
           681 => x"81",
           682 => x"52",
           683 => x"8c",
           684 => x"2a",
           685 => x"51",
           686 => x"38",
           687 => x"81",
           688 => x"06",
           689 => x"80",
           690 => x"71",
           691 => x"81",
           692 => x"70",
           693 => x"0b",
           694 => x"c0",
           695 => x"c0",
           696 => x"70",
           697 => x"38",
           698 => x"90",
           699 => x"0c",
           700 => x"04",
           701 => x"77",
           702 => x"33",
           703 => x"76",
           704 => x"38",
           705 => x"05",
           706 => x"0b",
           707 => x"33",
           708 => x"c0",
           709 => x"72",
           710 => x"38",
           711 => x"94",
           712 => x"70",
           713 => x"81",
           714 => x"52",
           715 => x"8c",
           716 => x"2a",
           717 => x"51",
           718 => x"38",
           719 => x"81",
           720 => x"06",
           721 => x"80",
           722 => x"71",
           723 => x"81",
           724 => x"70",
           725 => x"0b",
           726 => x"c0",
           727 => x"c0",
           728 => x"70",
           729 => x"38",
           730 => x"90",
           731 => x"0c",
           732 => x"33",
           733 => x"ff",
           734 => x"91",
           735 => x"87",
           736 => x"ff",
           737 => x"0b",
           738 => x"33",
           739 => x"94",
           740 => x"80",
           741 => x"87",
           742 => x"51",
           743 => x"82",
           744 => x"06",
           745 => x"70",
           746 => x"38",
           747 => x"cb",
           748 => x"87",
           749 => x"52",
           750 => x"86",
           751 => x"94",
           752 => x"08",
           753 => x"06",
           754 => x"0c",
           755 => x"0d",
           756 => x"0d",
           757 => x"cb",
           758 => x"87",
           759 => x"52",
           760 => x"86",
           761 => x"94",
           762 => x"08",
           763 => x"70",
           764 => x"51",
           765 => x"70",
           766 => x"38",
           767 => x"cb",
           768 => x"87",
           769 => x"52",
           770 => x"86",
           771 => x"94",
           772 => x"08",
           773 => x"70",
           774 => x"53",
           775 => x"d3",
           776 => x"3d",
           777 => x"3d",
           778 => x"9e",
           779 => x"70",
           780 => x"06",
           781 => x"70",
           782 => x"9f",
           783 => x"c4",
           784 => x"9e",
           785 => x"0c",
           786 => x"c0",
           787 => x"71",
           788 => x"11",
           789 => x"8c",
           790 => x"52",
           791 => x"c0",
           792 => x"71",
           793 => x"11",
           794 => x"94",
           795 => x"52",
           796 => x"c0",
           797 => x"71",
           798 => x"11",
           799 => x"a4",
           800 => x"52",
           801 => x"c0",
           802 => x"71",
           803 => x"11",
           804 => x"ac",
           805 => x"52",
           806 => x"52",
           807 => x"23",
           808 => x"c0",
           809 => x"71",
           810 => x"0b",
           811 => x"ad",
           812 => x"0b",
           813 => x"88",
           814 => x"80",
           815 => x"53",
           816 => x"83",
           817 => x"72",
           818 => x"0b",
           819 => x"88",
           820 => x"80",
           821 => x"52",
           822 => x"2e",
           823 => x"52",
           824 => x"f2",
           825 => x"87",
           826 => x"08",
           827 => x"80",
           828 => x"52",
           829 => x"83",
           830 => x"71",
           831 => x"34",
           832 => x"c0",
           833 => x"70",
           834 => x"51",
           835 => x"80",
           836 => x"81",
           837 => x"cb",
           838 => x"0b",
           839 => x"88",
           840 => x"80",
           841 => x"52",
           842 => x"83",
           843 => x"71",
           844 => x"34",
           845 => x"c0",
           846 => x"70",
           847 => x"51",
           848 => x"80",
           849 => x"81",
           850 => x"cb",
           851 => x"0b",
           852 => x"88",
           853 => x"80",
           854 => x"52",
           855 => x"83",
           856 => x"71",
           857 => x"34",
           858 => x"c0",
           859 => x"70",
           860 => x"51",
           861 => x"80",
           862 => x"81",
           863 => x"cb",
           864 => x"cb",
           865 => x"c0",
           866 => x"08",
           867 => x"06",
           868 => x"51",
           869 => x"70",
           870 => x"05",
           871 => x"54",
           872 => x"70",
           873 => x"52",
           874 => x"2e",
           875 => x"52",
           876 => x"80",
           877 => x"9e",
           878 => x"88",
           879 => x"52",
           880 => x"83",
           881 => x"71",
           882 => x"34",
           883 => x"88",
           884 => x"06",
           885 => x"91",
           886 => x"85",
           887 => x"fc",
           888 => x"b6",
           889 => x"be",
           890 => x"f0",
           891 => x"80",
           892 => x"91",
           893 => x"84",
           894 => x"b6",
           895 => x"a6",
           896 => x"f1",
           897 => x"55",
           898 => x"91",
           899 => x"08",
           900 => x"c4",
           901 => x"b7",
           902 => x"84",
           903 => x"f2",
           904 => x"55",
           905 => x"90",
           906 => x"08",
           907 => x"08",
           908 => x"a8",
           909 => x"3f",
           910 => x"70",
           911 => x"73",
           912 => x"15",
           913 => x"80",
           914 => x"91",
           915 => x"08",
           916 => x"08",
           917 => x"b7",
           918 => x"c4",
           919 => x"f5",
           920 => x"80",
           921 => x"91",
           922 => x"83",
           923 => x"cb",
           924 => x"73",
           925 => x"38",
           926 => x"51",
           927 => x"91",
           928 => x"54",
           929 => x"88",
           930 => x"88",
           931 => x"3f",
           932 => x"70",
           933 => x"73",
           934 => x"38",
           935 => x"52",
           936 => x"51",
           937 => x"91",
           938 => x"54",
           939 => x"88",
           940 => x"b4",
           941 => x"3f",
           942 => x"70",
           943 => x"73",
           944 => x"38",
           945 => x"52",
           946 => x"51",
           947 => x"91",
           948 => x"82",
           949 => x"cb",
           950 => x"70",
           951 => x"08",
           952 => x"f8",
           953 => x"88",
           954 => x"08",
           955 => x"a0",
           956 => x"3f",
           957 => x"52",
           958 => x"51",
           959 => x"8c",
           960 => x"91",
           961 => x"88",
           962 => x"15",
           963 => x"ba",
           964 => x"8c",
           965 => x"0d",
           966 => x"0d",
           967 => x"33",
           968 => x"26",
           969 => x"10",
           970 => x"91",
           971 => x"52",
           972 => x"91",
           973 => x"f7",
           974 => x"39",
           975 => x"51",
           976 => x"a3",
           977 => x"d0",
           978 => x"3f",
           979 => x"ba",
           980 => x"a0",
           981 => x"91",
           982 => x"f7",
           983 => x"39",
           984 => x"51",
           985 => x"83",
           986 => x"71",
           987 => x"04",
           988 => x"c0",
           989 => x"04",
           990 => x"87",
           991 => x"70",
           992 => x"80",
           993 => x"74",
           994 => x"cc",
           995 => x"0c",
           996 => x"04",
           997 => x"87",
           998 => x"70",
           999 => x"80",
          1000 => x"72",
          1001 => x"70",
          1002 => x"08",
          1003 => x"cc",
          1004 => x"0c",
          1005 => x"0d",
          1006 => x"80",
          1007 => x"96",
          1008 => x"fe",
          1009 => x"93",
          1010 => x"72",
          1011 => x"81",
          1012 => x"8d",
          1013 => x"91",
          1014 => x"80",
          1015 => x"91",
          1016 => x"52",
          1017 => x"91",
          1018 => x"81",
          1019 => x"e0",
          1020 => x"91",
          1021 => x"80",
          1022 => x"72",
          1023 => x"d8",
          1024 => x"2d",
          1025 => x"04",
          1026 => x"02",
          1027 => x"91",
          1028 => x"76",
          1029 => x"0c",
          1030 => x"a7",
          1031 => x"d3",
          1032 => x"3d",
          1033 => x"3d",
          1034 => x"33",
          1035 => x"80",
          1036 => x"72",
          1037 => x"54",
          1038 => x"87",
          1039 => x"52",
          1040 => x"84",
          1041 => x"fd",
          1042 => x"91",
          1043 => x"77",
          1044 => x"0c",
          1045 => x"55",
          1046 => x"2e",
          1047 => x"70",
          1048 => x"33",
          1049 => x"3f",
          1050 => x"71",
          1051 => x"91",
          1052 => x"85",
          1053 => x"ec",
          1054 => x"68",
          1055 => x"70",
          1056 => x"33",
          1057 => x"2e",
          1058 => x"75",
          1059 => x"38",
          1060 => x"af",
          1061 => x"80",
          1062 => x"81",
          1063 => x"58",
          1064 => x"b0",
          1065 => x"06",
          1066 => x"79",
          1067 => x"5b",
          1068 => x"92",
          1069 => x"2e",
          1070 => x"8a",
          1071 => x"70",
          1072 => x"33",
          1073 => x"aa",
          1074 => x"06",
          1075 => x"84",
          1076 => x"7b",
          1077 => x"5d",
          1078 => x"5d",
          1079 => x"d0",
          1080 => x"89",
          1081 => x"79",
          1082 => x"d0",
          1083 => x"81",
          1084 => x"d0",
          1085 => x"5a",
          1086 => x"eb",
          1087 => x"ec",
          1088 => x"70",
          1089 => x"25",
          1090 => x"32",
          1091 => x"72",
          1092 => x"73",
          1093 => x"52",
          1094 => x"73",
          1095 => x"38",
          1096 => x"79",
          1097 => x"5b",
          1098 => x"75",
          1099 => x"ec",
          1100 => x"80",
          1101 => x"89",
          1102 => x"70",
          1103 => x"56",
          1104 => x"15",
          1105 => x"26",
          1106 => x"72",
          1107 => x"b0",
          1108 => x"72",
          1109 => x"84",
          1110 => x"57",
          1111 => x"75",
          1112 => x"72",
          1113 => x"38",
          1114 => x"16",
          1115 => x"54",
          1116 => x"38",
          1117 => x"70",
          1118 => x"53",
          1119 => x"73",
          1120 => x"53",
          1121 => x"99",
          1122 => x"2a",
          1123 => x"a0",
          1124 => x"3f",
          1125 => x"73",
          1126 => x"53",
          1127 => x"ef",
          1128 => x"fd",
          1129 => x"81",
          1130 => x"72",
          1131 => x"ce",
          1132 => x"fc",
          1133 => x"81",
          1134 => x"79",
          1135 => x"38",
          1136 => x"7b",
          1137 => x"12",
          1138 => x"53",
          1139 => x"fd",
          1140 => x"5b",
          1141 => x"5b",
          1142 => x"5b",
          1143 => x"5b",
          1144 => x"51",
          1145 => x"fd",
          1146 => x"82",
          1147 => x"06",
          1148 => x"80",
          1149 => x"7b",
          1150 => x"08",
          1151 => x"9c",
          1152 => x"c4",
          1153 => x"06",
          1154 => x"84",
          1155 => x"59",
          1156 => x"39",
          1157 => x"71",
          1158 => x"53",
          1159 => x"32",
          1160 => x"72",
          1161 => x"70",
          1162 => x"06",
          1163 => x"53",
          1164 => x"88",
          1165 => x"7d",
          1166 => x"57",
          1167 => x"52",
          1168 => x"a8",
          1169 => x"c8",
          1170 => x"06",
          1171 => x"52",
          1172 => x"3f",
          1173 => x"08",
          1174 => x"27",
          1175 => x"a7",
          1176 => x"ff",
          1177 => x"54",
          1178 => x"2e",
          1179 => x"14",
          1180 => x"06",
          1181 => x"3d",
          1182 => x"05",
          1183 => x"54",
          1184 => x"81",
          1185 => x"70",
          1186 => x"2a",
          1187 => x"27",
          1188 => x"54",
          1189 => x"a6",
          1190 => x"2a",
          1191 => x"51",
          1192 => x"2e",
          1193 => x"3d",
          1194 => x"05",
          1195 => x"34",
          1196 => x"77",
          1197 => x"54",
          1198 => x"72",
          1199 => x"55",
          1200 => x"70",
          1201 => x"53",
          1202 => x"73",
          1203 => x"53",
          1204 => x"99",
          1205 => x"2a",
          1206 => x"74",
          1207 => x"3f",
          1208 => x"73",
          1209 => x"53",
          1210 => x"ef",
          1211 => x"97",
          1212 => x"11",
          1213 => x"54",
          1214 => x"3f",
          1215 => x"73",
          1216 => x"53",
          1217 => x"fa",
          1218 => x"51",
          1219 => x"73",
          1220 => x"53",
          1221 => x"f2",
          1222 => x"39",
          1223 => x"04",
          1224 => x"86",
          1225 => x"84",
          1226 => x"55",
          1227 => x"fa",
          1228 => x"3d",
          1229 => x"3d",
          1230 => x"d3",
          1231 => x"3d",
          1232 => x"75",
          1233 => x"3f",
          1234 => x"08",
          1235 => x"34",
          1236 => x"d3",
          1237 => x"3d",
          1238 => x"3d",
          1239 => x"d8",
          1240 => x"d3",
          1241 => x"3d",
          1242 => x"77",
          1243 => x"87",
          1244 => x"d3",
          1245 => x"3d",
          1246 => x"3d",
          1247 => x"57",
          1248 => x"91",
          1249 => x"73",
          1250 => x"38",
          1251 => x"53",
          1252 => x"80",
          1253 => x"dc",
          1254 => x"2d",
          1255 => x"08",
          1256 => x"54",
          1257 => x"e6",
          1258 => x"2e",
          1259 => x"73",
          1260 => x"30",
          1261 => x"78",
          1262 => x"72",
          1263 => x"52",
          1264 => x"72",
          1265 => x"38",
          1266 => x"81",
          1267 => x"55",
          1268 => x"c1",
          1269 => x"25",
          1270 => x"ff",
          1271 => x"72",
          1272 => x"38",
          1273 => x"73",
          1274 => x"15",
          1275 => x"06",
          1276 => x"cf",
          1277 => x"39",
          1278 => x"80",
          1279 => x"51",
          1280 => x"81",
          1281 => x"d3",
          1282 => x"3d",
          1283 => x"3d",
          1284 => x"dc",
          1285 => x"d3",
          1286 => x"53",
          1287 => x"fe",
          1288 => x"91",
          1289 => x"84",
          1290 => x"f8",
          1291 => x"7c",
          1292 => x"70",
          1293 => x"08",
          1294 => x"54",
          1295 => x"2e",
          1296 => x"92",
          1297 => x"81",
          1298 => x"74",
          1299 => x"55",
          1300 => x"2e",
          1301 => x"ad",
          1302 => x"06",
          1303 => x"75",
          1304 => x"0c",
          1305 => x"33",
          1306 => x"73",
          1307 => x"81",
          1308 => x"38",
          1309 => x"05",
          1310 => x"08",
          1311 => x"53",
          1312 => x"2e",
          1313 => x"80",
          1314 => x"81",
          1315 => x"90",
          1316 => x"76",
          1317 => x"70",
          1318 => x"57",
          1319 => x"82",
          1320 => x"05",
          1321 => x"08",
          1322 => x"54",
          1323 => x"81",
          1324 => x"27",
          1325 => x"d0",
          1326 => x"56",
          1327 => x"73",
          1328 => x"80",
          1329 => x"14",
          1330 => x"72",
          1331 => x"e8",
          1332 => x"80",
          1333 => x"39",
          1334 => x"dc",
          1335 => x"80",
          1336 => x"27",
          1337 => x"80",
          1338 => x"89",
          1339 => x"70",
          1340 => x"55",
          1341 => x"70",
          1342 => x"55",
          1343 => x"27",
          1344 => x"14",
          1345 => x"06",
          1346 => x"74",
          1347 => x"73",
          1348 => x"38",
          1349 => x"14",
          1350 => x"05",
          1351 => x"08",
          1352 => x"54",
          1353 => x"26",
          1354 => x"77",
          1355 => x"38",
          1356 => x"75",
          1357 => x"56",
          1358 => x"c8",
          1359 => x"0d",
          1360 => x"0d",
          1361 => x"55",
          1362 => x"0c",
          1363 => x"33",
          1364 => x"73",
          1365 => x"81",
          1366 => x"74",
          1367 => x"75",
          1368 => x"70",
          1369 => x"73",
          1370 => x"38",
          1371 => x"09",
          1372 => x"38",
          1373 => x"11",
          1374 => x"08",
          1375 => x"54",
          1376 => x"2e",
          1377 => x"80",
          1378 => x"08",
          1379 => x"0c",
          1380 => x"33",
          1381 => x"80",
          1382 => x"38",
          1383 => x"2e",
          1384 => x"a1",
          1385 => x"81",
          1386 => x"75",
          1387 => x"56",
          1388 => x"c1",
          1389 => x"08",
          1390 => x"0c",
          1391 => x"33",
          1392 => x"b1",
          1393 => x"a0",
          1394 => x"82",
          1395 => x"53",
          1396 => x"57",
          1397 => x"9d",
          1398 => x"39",
          1399 => x"80",
          1400 => x"26",
          1401 => x"8b",
          1402 => x"80",
          1403 => x"56",
          1404 => x"8a",
          1405 => x"a0",
          1406 => x"c5",
          1407 => x"74",
          1408 => x"e0",
          1409 => x"ff",
          1410 => x"d0",
          1411 => x"ff",
          1412 => x"90",
          1413 => x"38",
          1414 => x"81",
          1415 => x"53",
          1416 => x"c5",
          1417 => x"27",
          1418 => x"76",
          1419 => x"08",
          1420 => x"0c",
          1421 => x"33",
          1422 => x"73",
          1423 => x"bd",
          1424 => x"2e",
          1425 => x"30",
          1426 => x"0c",
          1427 => x"91",
          1428 => x"8a",
          1429 => x"ff",
          1430 => x"8f",
          1431 => x"81",
          1432 => x"26",
          1433 => x"cc",
          1434 => x"52",
          1435 => x"c8",
          1436 => x"0d",
          1437 => x"0d",
          1438 => x"33",
          1439 => x"9b",
          1440 => x"53",
          1441 => x"81",
          1442 => x"38",
          1443 => x"87",
          1444 => x"05",
          1445 => x"73",
          1446 => x"38",
          1447 => x"71",
          1448 => x"90",
          1449 => x"92",
          1450 => x"81",
          1451 => x"0b",
          1452 => x"8c",
          1453 => x"87",
          1454 => x"54",
          1455 => x"82",
          1456 => x"70",
          1457 => x"38",
          1458 => x"70",
          1459 => x"90",
          1460 => x"92",
          1461 => x"08",
          1462 => x"06",
          1463 => x"92",
          1464 => x"98",
          1465 => x"70",
          1466 => x"38",
          1467 => x"84",
          1468 => x"cc",
          1469 => x"51",
          1470 => x"c8",
          1471 => x"0d",
          1472 => x"0d",
          1473 => x"02",
          1474 => x"c3",
          1475 => x"41",
          1476 => x"73",
          1477 => x"bf",
          1478 => x"c8",
          1479 => x"7b",
          1480 => x"81",
          1481 => x"70",
          1482 => x"c0",
          1483 => x"84",
          1484 => x"92",
          1485 => x"c0",
          1486 => x"72",
          1487 => x"5b",
          1488 => x"0c",
          1489 => x"80",
          1490 => x"0c",
          1491 => x"0c",
          1492 => x"85",
          1493 => x"06",
          1494 => x"71",
          1495 => x"38",
          1496 => x"71",
          1497 => x"05",
          1498 => x"17",
          1499 => x"06",
          1500 => x"2e",
          1501 => x"08",
          1502 => x"38",
          1503 => x"71",
          1504 => x"38",
          1505 => x"2e",
          1506 => x"75",
          1507 => x"92",
          1508 => x"72",
          1509 => x"06",
          1510 => x"f7",
          1511 => x"5b",
          1512 => x"80",
          1513 => x"70",
          1514 => x"5f",
          1515 => x"80",
          1516 => x"73",
          1517 => x"06",
          1518 => x"38",
          1519 => x"ff",
          1520 => x"fc",
          1521 => x"52",
          1522 => x"83",
          1523 => x"71",
          1524 => x"d3",
          1525 => x"3d",
          1526 => x"3d",
          1527 => x"64",
          1528 => x"bf",
          1529 => x"40",
          1530 => x"73",
          1531 => x"e7",
          1532 => x"c8",
          1533 => x"7a",
          1534 => x"81",
          1535 => x"5c",
          1536 => x"8c",
          1537 => x"87",
          1538 => x"11",
          1539 => x"84",
          1540 => x"5b",
          1541 => x"85",
          1542 => x"c0",
          1543 => x"7b",
          1544 => x"82",
          1545 => x"53",
          1546 => x"84",
          1547 => x"06",
          1548 => x"71",
          1549 => x"38",
          1550 => x"05",
          1551 => x"0c",
          1552 => x"73",
          1553 => x"81",
          1554 => x"71",
          1555 => x"38",
          1556 => x"71",
          1557 => x"08",
          1558 => x"2e",
          1559 => x"84",
          1560 => x"38",
          1561 => x"87",
          1562 => x"1d",
          1563 => x"70",
          1564 => x"52",
          1565 => x"ff",
          1566 => x"39",
          1567 => x"81",
          1568 => x"80",
          1569 => x"52",
          1570 => x"90",
          1571 => x"80",
          1572 => x"71",
          1573 => x"7c",
          1574 => x"38",
          1575 => x"80",
          1576 => x"80",
          1577 => x"81",
          1578 => x"73",
          1579 => x"0c",
          1580 => x"04",
          1581 => x"7d",
          1582 => x"af",
          1583 => x"88",
          1584 => x"33",
          1585 => x"56",
          1586 => x"3f",
          1587 => x"08",
          1588 => x"83",
          1589 => x"38",
          1590 => x"74",
          1591 => x"72",
          1592 => x"38",
          1593 => x"8a",
          1594 => x"72",
          1595 => x"38",
          1596 => x"90",
          1597 => x"92",
          1598 => x"08",
          1599 => x"39",
          1600 => x"76",
          1601 => x"8b",
          1602 => x"76",
          1603 => x"83",
          1604 => x"73",
          1605 => x"0c",
          1606 => x"04",
          1607 => x"73",
          1608 => x"12",
          1609 => x"2b",
          1610 => x"d3",
          1611 => x"52",
          1612 => x"0d",
          1613 => x"0d",
          1614 => x"33",
          1615 => x"71",
          1616 => x"88",
          1617 => x"14",
          1618 => x"74",
          1619 => x"2b",
          1620 => x"c8",
          1621 => x"56",
          1622 => x"3d",
          1623 => x"3d",
          1624 => x"84",
          1625 => x"22",
          1626 => x"72",
          1627 => x"54",
          1628 => x"2a",
          1629 => x"34",
          1630 => x"04",
          1631 => x"73",
          1632 => x"70",
          1633 => x"05",
          1634 => x"88",
          1635 => x"72",
          1636 => x"54",
          1637 => x"2a",
          1638 => x"70",
          1639 => x"34",
          1640 => x"51",
          1641 => x"83",
          1642 => x"fe",
          1643 => x"75",
          1644 => x"51",
          1645 => x"93",
          1646 => x"81",
          1647 => x"73",
          1648 => x"55",
          1649 => x"51",
          1650 => x"84",
          1651 => x"fe",
          1652 => x"77",
          1653 => x"53",
          1654 => x"81",
          1655 => x"ff",
          1656 => x"f4",
          1657 => x"0d",
          1658 => x"0d",
          1659 => x"56",
          1660 => x"70",
          1661 => x"33",
          1662 => x"05",
          1663 => x"71",
          1664 => x"56",
          1665 => x"72",
          1666 => x"38",
          1667 => x"e2",
          1668 => x"d3",
          1669 => x"3d",
          1670 => x"3d",
          1671 => x"71",
          1672 => x"52",
          1673 => x"99",
          1674 => x"2e",
          1675 => x"12",
          1676 => x"52",
          1677 => x"89",
          1678 => x"2e",
          1679 => x"ee",
          1680 => x"91",
          1681 => x"84",
          1682 => x"80",
          1683 => x"c8",
          1684 => x"0b",
          1685 => x"0c",
          1686 => x"0d",
          1687 => x"0b",
          1688 => x"56",
          1689 => x"2e",
          1690 => x"81",
          1691 => x"08",
          1692 => x"70",
          1693 => x"33",
          1694 => x"de",
          1695 => x"c8",
          1696 => x"09",
          1697 => x"38",
          1698 => x"08",
          1699 => x"b0",
          1700 => x"17",
          1701 => x"74",
          1702 => x"27",
          1703 => x"16",
          1704 => x"82",
          1705 => x"06",
          1706 => x"54",
          1707 => x"9c",
          1708 => x"53",
          1709 => x"16",
          1710 => x"9e",
          1711 => x"81",
          1712 => x"d3",
          1713 => x"3d",
          1714 => x"3d",
          1715 => x"56",
          1716 => x"b0",
          1717 => x"2e",
          1718 => x"51",
          1719 => x"91",
          1720 => x"56",
          1721 => x"08",
          1722 => x"54",
          1723 => x"17",
          1724 => x"33",
          1725 => x"3f",
          1726 => x"08",
          1727 => x"38",
          1728 => x"56",
          1729 => x"0c",
          1730 => x"c8",
          1731 => x"0d",
          1732 => x"0d",
          1733 => x"57",
          1734 => x"91",
          1735 => x"58",
          1736 => x"08",
          1737 => x"76",
          1738 => x"83",
          1739 => x"06",
          1740 => x"84",
          1741 => x"78",
          1742 => x"81",
          1743 => x"38",
          1744 => x"91",
          1745 => x"52",
          1746 => x"52",
          1747 => x"3f",
          1748 => x"52",
          1749 => x"51",
          1750 => x"84",
          1751 => x"d2",
          1752 => x"fc",
          1753 => x"8a",
          1754 => x"52",
          1755 => x"51",
          1756 => x"90",
          1757 => x"84",
          1758 => x"fb",
          1759 => x"17",
          1760 => x"a0",
          1761 => x"f4",
          1762 => x"08",
          1763 => x"b0",
          1764 => x"55",
          1765 => x"81",
          1766 => x"f8",
          1767 => x"84",
          1768 => x"53",
          1769 => x"17",
          1770 => x"88",
          1771 => x"c8",
          1772 => x"83",
          1773 => x"77",
          1774 => x"0c",
          1775 => x"04",
          1776 => x"77",
          1777 => x"12",
          1778 => x"55",
          1779 => x"56",
          1780 => x"8d",
          1781 => x"22",
          1782 => x"ac",
          1783 => x"57",
          1784 => x"d3",
          1785 => x"3d",
          1786 => x"3d",
          1787 => x"70",
          1788 => x"55",
          1789 => x"88",
          1790 => x"08",
          1791 => x"38",
          1792 => x"d9",
          1793 => x"33",
          1794 => x"82",
          1795 => x"38",
          1796 => x"89",
          1797 => x"2e",
          1798 => x"bf",
          1799 => x"2e",
          1800 => x"81",
          1801 => x"81",
          1802 => x"89",
          1803 => x"08",
          1804 => x"52",
          1805 => x"3f",
          1806 => x"08",
          1807 => x"76",
          1808 => x"14",
          1809 => x"81",
          1810 => x"2a",
          1811 => x"05",
          1812 => x"59",
          1813 => x"f2",
          1814 => x"c8",
          1815 => x"38",
          1816 => x"06",
          1817 => x"33",
          1818 => x"7a",
          1819 => x"06",
          1820 => x"5a",
          1821 => x"53",
          1822 => x"38",
          1823 => x"06",
          1824 => x"39",
          1825 => x"a4",
          1826 => x"52",
          1827 => x"ba",
          1828 => x"c8",
          1829 => x"38",
          1830 => x"ff",
          1831 => x"b4",
          1832 => x"f8",
          1833 => x"c8",
          1834 => x"ff",
          1835 => x"39",
          1836 => x"a4",
          1837 => x"52",
          1838 => x"8e",
          1839 => x"c8",
          1840 => x"74",
          1841 => x"fc",
          1842 => x"b4",
          1843 => x"e5",
          1844 => x"c8",
          1845 => x"06",
          1846 => x"81",
          1847 => x"d3",
          1848 => x"3d",
          1849 => x"3d",
          1850 => x"7f",
          1851 => x"82",
          1852 => x"27",
          1853 => x"73",
          1854 => x"27",
          1855 => x"74",
          1856 => x"77",
          1857 => x"38",
          1858 => x"89",
          1859 => x"2e",
          1860 => x"91",
          1861 => x"2e",
          1862 => x"82",
          1863 => x"81",
          1864 => x"89",
          1865 => x"08",
          1866 => x"52",
          1867 => x"3f",
          1868 => x"08",
          1869 => x"c8",
          1870 => x"38",
          1871 => x"06",
          1872 => x"81",
          1873 => x"06",
          1874 => x"58",
          1875 => x"80",
          1876 => x"75",
          1877 => x"f0",
          1878 => x"8f",
          1879 => x"58",
          1880 => x"34",
          1881 => x"16",
          1882 => x"2a",
          1883 => x"05",
          1884 => x"fa",
          1885 => x"d3",
          1886 => x"91",
          1887 => x"81",
          1888 => x"83",
          1889 => x"b4",
          1890 => x"06",
          1891 => x"57",
          1892 => x"72",
          1893 => x"88",
          1894 => x"57",
          1895 => x"81",
          1896 => x"54",
          1897 => x"81",
          1898 => x"34",
          1899 => x"73",
          1900 => x"16",
          1901 => x"74",
          1902 => x"3f",
          1903 => x"08",
          1904 => x"c8",
          1905 => x"38",
          1906 => x"ff",
          1907 => x"14",
          1908 => x"75",
          1909 => x"51",
          1910 => x"81",
          1911 => x"34",
          1912 => x"73",
          1913 => x"16",
          1914 => x"74",
          1915 => x"3f",
          1916 => x"08",
          1917 => x"c8",
          1918 => x"75",
          1919 => x"74",
          1920 => x"fc",
          1921 => x"b4",
          1922 => x"51",
          1923 => x"a5",
          1924 => x"c8",
          1925 => x"06",
          1926 => x"72",
          1927 => x"3f",
          1928 => x"16",
          1929 => x"d3",
          1930 => x"3d",
          1931 => x"3d",
          1932 => x"7d",
          1933 => x"58",
          1934 => x"74",
          1935 => x"98",
          1936 => x"26",
          1937 => x"56",
          1938 => x"75",
          1939 => x"38",
          1940 => x"52",
          1941 => x"8e",
          1942 => x"c8",
          1943 => x"d3",
          1944 => x"f4",
          1945 => x"82",
          1946 => x"39",
          1947 => x"e8",
          1948 => x"c8",
          1949 => x"e0",
          1950 => x"76",
          1951 => x"3f",
          1952 => x"08",
          1953 => x"c8",
          1954 => x"80",
          1955 => x"d3",
          1956 => x"2e",
          1957 => x"d3",
          1958 => x"2e",
          1959 => x"53",
          1960 => x"51",
          1961 => x"91",
          1962 => x"c5",
          1963 => x"08",
          1964 => x"90",
          1965 => x"27",
          1966 => x"15",
          1967 => x"90",
          1968 => x"15",
          1969 => x"54",
          1970 => x"34",
          1971 => x"15",
          1972 => x"ff",
          1973 => x"56",
          1974 => x"c8",
          1975 => x"0d",
          1976 => x"0d",
          1977 => x"08",
          1978 => x"7a",
          1979 => x"19",
          1980 => x"80",
          1981 => x"98",
          1982 => x"26",
          1983 => x"58",
          1984 => x"52",
          1985 => x"e2",
          1986 => x"74",
          1987 => x"08",
          1988 => x"38",
          1989 => x"08",
          1990 => x"c8",
          1991 => x"82",
          1992 => x"d3",
          1993 => x"98",
          1994 => x"d3",
          1995 => x"82",
          1996 => x"58",
          1997 => x"19",
          1998 => x"82",
          1999 => x"57",
          2000 => x"09",
          2001 => x"db",
          2002 => x"57",
          2003 => x"77",
          2004 => x"82",
          2005 => x"7b",
          2006 => x"3f",
          2007 => x"08",
          2008 => x"91",
          2009 => x"81",
          2010 => x"06",
          2011 => x"d3",
          2012 => x"75",
          2013 => x"30",
          2014 => x"80",
          2015 => x"07",
          2016 => x"52",
          2017 => x"81",
          2018 => x"80",
          2019 => x"8c",
          2020 => x"81",
          2021 => x"38",
          2022 => x"08",
          2023 => x"75",
          2024 => x"76",
          2025 => x"77",
          2026 => x"57",
          2027 => x"77",
          2028 => x"82",
          2029 => x"26",
          2030 => x"76",
          2031 => x"f8",
          2032 => x"d3",
          2033 => x"91",
          2034 => x"80",
          2035 => x"80",
          2036 => x"c8",
          2037 => x"09",
          2038 => x"38",
          2039 => x"08",
          2040 => x"32",
          2041 => x"72",
          2042 => x"70",
          2043 => x"52",
          2044 => x"80",
          2045 => x"78",
          2046 => x"06",
          2047 => x"80",
          2048 => x"39",
          2049 => x"52",
          2050 => x"da",
          2051 => x"c8",
          2052 => x"c8",
          2053 => x"91",
          2054 => x"07",
          2055 => x"30",
          2056 => x"9f",
          2057 => x"52",
          2058 => x"56",
          2059 => x"8f",
          2060 => x"7a",
          2061 => x"f9",
          2062 => x"d3",
          2063 => x"75",
          2064 => x"8c",
          2065 => x"19",
          2066 => x"54",
          2067 => x"74",
          2068 => x"90",
          2069 => x"05",
          2070 => x"84",
          2071 => x"07",
          2072 => x"1a",
          2073 => x"ff",
          2074 => x"2e",
          2075 => x"39",
          2076 => x"39",
          2077 => x"39",
          2078 => x"55",
          2079 => x"c8",
          2080 => x"0d",
          2081 => x"0d",
          2082 => x"57",
          2083 => x"81",
          2084 => x"c8",
          2085 => x"38",
          2086 => x"51",
          2087 => x"91",
          2088 => x"91",
          2089 => x"b0",
          2090 => x"84",
          2091 => x"52",
          2092 => x"52",
          2093 => x"3f",
          2094 => x"58",
          2095 => x"39",
          2096 => x"8a",
          2097 => x"75",
          2098 => x"38",
          2099 => x"1a",
          2100 => x"81",
          2101 => x"ee",
          2102 => x"d3",
          2103 => x"2e",
          2104 => x"0b",
          2105 => x"56",
          2106 => x"2e",
          2107 => x"58",
          2108 => x"91",
          2109 => x"8b",
          2110 => x"f8",
          2111 => x"7c",
          2112 => x"56",
          2113 => x"80",
          2114 => x"38",
          2115 => x"53",
          2116 => x"86",
          2117 => x"81",
          2118 => x"90",
          2119 => x"17",
          2120 => x"aa",
          2121 => x"53",
          2122 => x"85",
          2123 => x"08",
          2124 => x"38",
          2125 => x"53",
          2126 => x"17",
          2127 => x"72",
          2128 => x"83",
          2129 => x"08",
          2130 => x"80",
          2131 => x"16",
          2132 => x"2b",
          2133 => x"75",
          2134 => x"73",
          2135 => x"f5",
          2136 => x"d3",
          2137 => x"91",
          2138 => x"ff",
          2139 => x"81",
          2140 => x"c8",
          2141 => x"38",
          2142 => x"91",
          2143 => x"26",
          2144 => x"58",
          2145 => x"74",
          2146 => x"74",
          2147 => x"38",
          2148 => x"51",
          2149 => x"91",
          2150 => x"98",
          2151 => x"94",
          2152 => x"58",
          2153 => x"80",
          2154 => x"85",
          2155 => x"97",
          2156 => x"2a",
          2157 => x"05",
          2158 => x"74",
          2159 => x"16",
          2160 => x"18",
          2161 => x"77",
          2162 => x"0c",
          2163 => x"04",
          2164 => x"79",
          2165 => x"90",
          2166 => x"05",
          2167 => x"55",
          2168 => x"76",
          2169 => x"80",
          2170 => x"0c",
          2171 => x"15",
          2172 => x"81",
          2173 => x"83",
          2174 => x"73",
          2175 => x"98",
          2176 => x"05",
          2177 => x"94",
          2178 => x"38",
          2179 => x"88",
          2180 => x"53",
          2181 => x"81",
          2182 => x"98",
          2183 => x"53",
          2184 => x"8a",
          2185 => x"11",
          2186 => x"06",
          2187 => x"81",
          2188 => x"15",
          2189 => x"51",
          2190 => x"91",
          2191 => x"54",
          2192 => x"0b",
          2193 => x"08",
          2194 => x"38",
          2195 => x"d3",
          2196 => x"2e",
          2197 => x"98",
          2198 => x"d3",
          2199 => x"80",
          2200 => x"8a",
          2201 => x"16",
          2202 => x"80",
          2203 => x"15",
          2204 => x"51",
          2205 => x"91",
          2206 => x"54",
          2207 => x"d3",
          2208 => x"2e",
          2209 => x"82",
          2210 => x"c8",
          2211 => x"bf",
          2212 => x"91",
          2213 => x"ff",
          2214 => x"91",
          2215 => x"52",
          2216 => x"e1",
          2217 => x"91",
          2218 => x"a3",
          2219 => x"16",
          2220 => x"76",
          2221 => x"3f",
          2222 => x"08",
          2223 => x"75",
          2224 => x"75",
          2225 => x"17",
          2226 => x"16",
          2227 => x"72",
          2228 => x"0c",
          2229 => x"04",
          2230 => x"7a",
          2231 => x"5a",
          2232 => x"52",
          2233 => x"93",
          2234 => x"c8",
          2235 => x"d3",
          2236 => x"e1",
          2237 => x"c8",
          2238 => x"16",
          2239 => x"51",
          2240 => x"91",
          2241 => x"54",
          2242 => x"08",
          2243 => x"91",
          2244 => x"9c",
          2245 => x"33",
          2246 => x"72",
          2247 => x"09",
          2248 => x"38",
          2249 => x"30",
          2250 => x"76",
          2251 => x"72",
          2252 => x"38",
          2253 => x"76",
          2254 => x"38",
          2255 => x"57",
          2256 => x"51",
          2257 => x"91",
          2258 => x"54",
          2259 => x"08",
          2260 => x"a6",
          2261 => x"2e",
          2262 => x"83",
          2263 => x"73",
          2264 => x"0c",
          2265 => x"04",
          2266 => x"76",
          2267 => x"54",
          2268 => x"91",
          2269 => x"83",
          2270 => x"76",
          2271 => x"53",
          2272 => x"2e",
          2273 => x"90",
          2274 => x"51",
          2275 => x"91",
          2276 => x"90",
          2277 => x"53",
          2278 => x"c8",
          2279 => x"0d",
          2280 => x"0d",
          2281 => x"83",
          2282 => x"54",
          2283 => x"55",
          2284 => x"3f",
          2285 => x"51",
          2286 => x"2e",
          2287 => x"8b",
          2288 => x"2a",
          2289 => x"51",
          2290 => x"86",
          2291 => x"f7",
          2292 => x"7d",
          2293 => x"76",
          2294 => x"98",
          2295 => x"2e",
          2296 => x"98",
          2297 => x"78",
          2298 => x"3f",
          2299 => x"08",
          2300 => x"c8",
          2301 => x"38",
          2302 => x"70",
          2303 => x"74",
          2304 => x"58",
          2305 => x"9c",
          2306 => x"11",
          2307 => x"06",
          2308 => x"06",
          2309 => x"53",
          2310 => x"34",
          2311 => x"32",
          2312 => x"ae",
          2313 => x"70",
          2314 => x"2a",
          2315 => x"51",
          2316 => x"2e",
          2317 => x"8f",
          2318 => x"80",
          2319 => x"54",
          2320 => x"2e",
          2321 => x"83",
          2322 => x"73",
          2323 => x"38",
          2324 => x"51",
          2325 => x"91",
          2326 => x"58",
          2327 => x"08",
          2328 => x"16",
          2329 => x"38",
          2330 => x"86",
          2331 => x"98",
          2332 => x"91",
          2333 => x"8b",
          2334 => x"f8",
          2335 => x"70",
          2336 => x"80",
          2337 => x"f8",
          2338 => x"d3",
          2339 => x"91",
          2340 => x"80",
          2341 => x"39",
          2342 => x"e6",
          2343 => x"08",
          2344 => x"ec",
          2345 => x"d3",
          2346 => x"91",
          2347 => x"80",
          2348 => x"16",
          2349 => x"51",
          2350 => x"2e",
          2351 => x"16",
          2352 => x"33",
          2353 => x"55",
          2354 => x"34",
          2355 => x"70",
          2356 => x"81",
          2357 => x"59",
          2358 => x"8b",
          2359 => x"52",
          2360 => x"85",
          2361 => x"c8",
          2362 => x"96",
          2363 => x"75",
          2364 => x"3f",
          2365 => x"08",
          2366 => x"c8",
          2367 => x"ff",
          2368 => x"54",
          2369 => x"c8",
          2370 => x"0d",
          2371 => x"0d",
          2372 => x"57",
          2373 => x"73",
          2374 => x"3f",
          2375 => x"08",
          2376 => x"c8",
          2377 => x"98",
          2378 => x"75",
          2379 => x"3f",
          2380 => x"08",
          2381 => x"c8",
          2382 => x"a0",
          2383 => x"c8",
          2384 => x"14",
          2385 => x"87",
          2386 => x"a0",
          2387 => x"14",
          2388 => x"d7",
          2389 => x"83",
          2390 => x"91",
          2391 => x"87",
          2392 => x"fc",
          2393 => x"70",
          2394 => x"08",
          2395 => x"56",
          2396 => x"3f",
          2397 => x"08",
          2398 => x"c8",
          2399 => x"9c",
          2400 => x"e5",
          2401 => x"0b",
          2402 => x"73",
          2403 => x"0c",
          2404 => x"04",
          2405 => x"78",
          2406 => x"80",
          2407 => x"34",
          2408 => x"80",
          2409 => x"38",
          2410 => x"55",
          2411 => x"14",
          2412 => x"16",
          2413 => x"72",
          2414 => x"38",
          2415 => x"09",
          2416 => x"38",
          2417 => x"73",
          2418 => x"81",
          2419 => x"75",
          2420 => x"52",
          2421 => x"13",
          2422 => x"55",
          2423 => x"05",
          2424 => x"13",
          2425 => x"55",
          2426 => x"c0",
          2427 => x"88",
          2428 => x"0b",
          2429 => x"9c",
          2430 => x"8b",
          2431 => x"17",
          2432 => x"08",
          2433 => x"e6",
          2434 => x"d3",
          2435 => x"0c",
          2436 => x"96",
          2437 => x"84",
          2438 => x"c8",
          2439 => x"23",
          2440 => x"98",
          2441 => x"f4",
          2442 => x"c8",
          2443 => x"23",
          2444 => x"04",
          2445 => x"7e",
          2446 => x"a0",
          2447 => x"5c",
          2448 => x"52",
          2449 => x"87",
          2450 => x"58",
          2451 => x"33",
          2452 => x"ae",
          2453 => x"06",
          2454 => x"78",
          2455 => x"81",
          2456 => x"32",
          2457 => x"9f",
          2458 => x"26",
          2459 => x"53",
          2460 => x"73",
          2461 => x"18",
          2462 => x"34",
          2463 => x"db",
          2464 => x"32",
          2465 => x"80",
          2466 => x"30",
          2467 => x"9f",
          2468 => x"56",
          2469 => x"80",
          2470 => x"86",
          2471 => x"26",
          2472 => x"76",
          2473 => x"a4",
          2474 => x"27",
          2475 => x"54",
          2476 => x"34",
          2477 => x"ce",
          2478 => x"70",
          2479 => x"59",
          2480 => x"76",
          2481 => x"38",
          2482 => x"70",
          2483 => x"dc",
          2484 => x"72",
          2485 => x"80",
          2486 => x"51",
          2487 => x"74",
          2488 => x"38",
          2489 => x"17",
          2490 => x"1a",
          2491 => x"55",
          2492 => x"2e",
          2493 => x"83",
          2494 => x"80",
          2495 => x"33",
          2496 => x"73",
          2497 => x"09",
          2498 => x"38",
          2499 => x"75",
          2500 => x"d2",
          2501 => x"39",
          2502 => x"70",
          2503 => x"25",
          2504 => x"07",
          2505 => x"73",
          2506 => x"38",
          2507 => x"70",
          2508 => x"32",
          2509 => x"80",
          2510 => x"2a",
          2511 => x"56",
          2512 => x"81",
          2513 => x"58",
          2514 => x"ed",
          2515 => x"2b",
          2516 => x"25",
          2517 => x"80",
          2518 => x"bb",
          2519 => x"57",
          2520 => x"e5",
          2521 => x"d3",
          2522 => x"2e",
          2523 => x"17",
          2524 => x"19",
          2525 => x"56",
          2526 => x"3f",
          2527 => x"08",
          2528 => x"38",
          2529 => x"73",
          2530 => x"38",
          2531 => x"f6",
          2532 => x"54",
          2533 => x"81",
          2534 => x"55",
          2535 => x"34",
          2536 => x"fe",
          2537 => x"52",
          2538 => x"51",
          2539 => x"91",
          2540 => x"80",
          2541 => x"9f",
          2542 => x"99",
          2543 => x"e0",
          2544 => x"ff",
          2545 => x"7a",
          2546 => x"74",
          2547 => x"58",
          2548 => x"76",
          2549 => x"86",
          2550 => x"2e",
          2551 => x"33",
          2552 => x"e5",
          2553 => x"06",
          2554 => x"7b",
          2555 => x"a0",
          2556 => x"38",
          2557 => x"54",
          2558 => x"54",
          2559 => x"54",
          2560 => x"34",
          2561 => x"91",
          2562 => x"8d",
          2563 => x"fa",
          2564 => x"70",
          2565 => x"80",
          2566 => x"51",
          2567 => x"af",
          2568 => x"81",
          2569 => x"70",
          2570 => x"54",
          2571 => x"2e",
          2572 => x"54",
          2573 => x"53",
          2574 => x"8c",
          2575 => x"08",
          2576 => x"b3",
          2577 => x"5a",
          2578 => x"33",
          2579 => x"72",
          2580 => x"81",
          2581 => x"81",
          2582 => x"70",
          2583 => x"54",
          2584 => x"2e",
          2585 => x"83",
          2586 => x"74",
          2587 => x"72",
          2588 => x"0b",
          2589 => x"79",
          2590 => x"53",
          2591 => x"9b",
          2592 => x"0b",
          2593 => x"80",
          2594 => x"f0",
          2595 => x"d3",
          2596 => x"81",
          2597 => x"55",
          2598 => x"89",
          2599 => x"52",
          2600 => x"90",
          2601 => x"c8",
          2602 => x"d3",
          2603 => x"8f",
          2604 => x"f7",
          2605 => x"d3",
          2606 => x"17",
          2607 => x"91",
          2608 => x"80",
          2609 => x"38",
          2610 => x"08",
          2611 => x"81",
          2612 => x"38",
          2613 => x"70",
          2614 => x"53",
          2615 => x"9a",
          2616 => x"2a",
          2617 => x"51",
          2618 => x"2e",
          2619 => x"ff",
          2620 => x"17",
          2621 => x"80",
          2622 => x"82",
          2623 => x"06",
          2624 => x"bb",
          2625 => x"b7",
          2626 => x"2a",
          2627 => x"51",
          2628 => x"38",
          2629 => x"70",
          2630 => x"81",
          2631 => x"54",
          2632 => x"fe",
          2633 => x"16",
          2634 => x"06",
          2635 => x"52",
          2636 => x"b4",
          2637 => x"c8",
          2638 => x"0c",
          2639 => x"74",
          2640 => x"0c",
          2641 => x"04",
          2642 => x"7c",
          2643 => x"08",
          2644 => x"59",
          2645 => x"80",
          2646 => x"38",
          2647 => x"05",
          2648 => x"ba",
          2649 => x"72",
          2650 => x"9f",
          2651 => x"51",
          2652 => x"e8",
          2653 => x"2e",
          2654 => x"81",
          2655 => x"33",
          2656 => x"52",
          2657 => x"92",
          2658 => x"72",
          2659 => x"d0",
          2660 => x"51",
          2661 => x"80",
          2662 => x"0b",
          2663 => x"5c",
          2664 => x"10",
          2665 => x"7a",
          2666 => x"51",
          2667 => x"05",
          2668 => x"70",
          2669 => x"33",
          2670 => x"53",
          2671 => x"99",
          2672 => x"e0",
          2673 => x"ff",
          2674 => x"ff",
          2675 => x"70",
          2676 => x"38",
          2677 => x"81",
          2678 => x"51",
          2679 => x"74",
          2680 => x"70",
          2681 => x"25",
          2682 => x"06",
          2683 => x"51",
          2684 => x"38",
          2685 => x"78",
          2686 => x"70",
          2687 => x"2a",
          2688 => x"07",
          2689 => x"51",
          2690 => x"8c",
          2691 => x"58",
          2692 => x"ff",
          2693 => x"39",
          2694 => x"86",
          2695 => x"7a",
          2696 => x"51",
          2697 => x"d3",
          2698 => x"70",
          2699 => x"0c",
          2700 => x"04",
          2701 => x"77",
          2702 => x"83",
          2703 => x"0b",
          2704 => x"78",
          2705 => x"e1",
          2706 => x"55",
          2707 => x"08",
          2708 => x"84",
          2709 => x"dd",
          2710 => x"d3",
          2711 => x"ff",
          2712 => x"83",
          2713 => x"d4",
          2714 => x"81",
          2715 => x"38",
          2716 => x"17",
          2717 => x"73",
          2718 => x"09",
          2719 => x"38",
          2720 => x"81",
          2721 => x"30",
          2722 => x"77",
          2723 => x"54",
          2724 => x"b4",
          2725 => x"73",
          2726 => x"09",
          2727 => x"38",
          2728 => x"bb",
          2729 => x"ea",
          2730 => x"bd",
          2731 => x"c8",
          2732 => x"d3",
          2733 => x"2e",
          2734 => x"53",
          2735 => x"52",
          2736 => x"51",
          2737 => x"91",
          2738 => x"55",
          2739 => x"08",
          2740 => x"38",
          2741 => x"91",
          2742 => x"87",
          2743 => x"f3",
          2744 => x"02",
          2745 => x"c7",
          2746 => x"54",
          2747 => x"7f",
          2748 => x"3f",
          2749 => x"08",
          2750 => x"80",
          2751 => x"c8",
          2752 => x"9e",
          2753 => x"c8",
          2754 => x"91",
          2755 => x"70",
          2756 => x"8c",
          2757 => x"2e",
          2758 => x"74",
          2759 => x"81",
          2760 => x"33",
          2761 => x"80",
          2762 => x"81",
          2763 => x"d6",
          2764 => x"d3",
          2765 => x"ff",
          2766 => x"06",
          2767 => x"99",
          2768 => x"2e",
          2769 => x"82",
          2770 => x"06",
          2771 => x"56",
          2772 => x"38",
          2773 => x"ca",
          2774 => x"34",
          2775 => x"34",
          2776 => x"15",
          2777 => x"8d",
          2778 => x"c8",
          2779 => x"06",
          2780 => x"54",
          2781 => x"72",
          2782 => x"76",
          2783 => x"38",
          2784 => x"70",
          2785 => x"53",
          2786 => x"86",
          2787 => x"70",
          2788 => x"5a",
          2789 => x"91",
          2790 => x"81",
          2791 => x"76",
          2792 => x"81",
          2793 => x"38",
          2794 => x"90",
          2795 => x"3d",
          2796 => x"05",
          2797 => x"f6",
          2798 => x"59",
          2799 => x"72",
          2800 => x"38",
          2801 => x"51",
          2802 => x"91",
          2803 => x"57",
          2804 => x"81",
          2805 => x"74",
          2806 => x"80",
          2807 => x"74",
          2808 => x"f0",
          2809 => x"53",
          2810 => x"80",
          2811 => x"79",
          2812 => x"fc",
          2813 => x"d3",
          2814 => x"ff",
          2815 => x"77",
          2816 => x"81",
          2817 => x"74",
          2818 => x"81",
          2819 => x"2e",
          2820 => x"8d",
          2821 => x"26",
          2822 => x"bf",
          2823 => x"fc",
          2824 => x"c8",
          2825 => x"ff",
          2826 => x"56",
          2827 => x"2e",
          2828 => x"84",
          2829 => x"ca",
          2830 => x"e0",
          2831 => x"c8",
          2832 => x"ff",
          2833 => x"8d",
          2834 => x"15",
          2835 => x"3f",
          2836 => x"08",
          2837 => x"16",
          2838 => x"15",
          2839 => x"34",
          2840 => x"33",
          2841 => x"8d",
          2842 => x"26",
          2843 => x"82",
          2844 => x"71",
          2845 => x"17",
          2846 => x"53",
          2847 => x"23",
          2848 => x"ff",
          2849 => x"80",
          2850 => x"ff",
          2851 => x"53",
          2852 => x"86",
          2853 => x"84",
          2854 => x"c5",
          2855 => x"fc",
          2856 => x"c8",
          2857 => x"23",
          2858 => x"08",
          2859 => x"06",
          2860 => x"8d",
          2861 => x"ea",
          2862 => x"15",
          2863 => x"3f",
          2864 => x"08",
          2865 => x"06",
          2866 => x"38",
          2867 => x"51",
          2868 => x"91",
          2869 => x"53",
          2870 => x"51",
          2871 => x"91",
          2872 => x"83",
          2873 => x"59",
          2874 => x"80",
          2875 => x"38",
          2876 => x"74",
          2877 => x"2a",
          2878 => x"8d",
          2879 => x"26",
          2880 => x"8a",
          2881 => x"72",
          2882 => x"ff",
          2883 => x"91",
          2884 => x"53",
          2885 => x"d3",
          2886 => x"2e",
          2887 => x"80",
          2888 => x"c8",
          2889 => x"ff",
          2890 => x"83",
          2891 => x"72",
          2892 => x"26",
          2893 => x"57",
          2894 => x"26",
          2895 => x"57",
          2896 => x"80",
          2897 => x"38",
          2898 => x"16",
          2899 => x"16",
          2900 => x"a4",
          2901 => x"1a",
          2902 => x"76",
          2903 => x"81",
          2904 => x"80",
          2905 => x"d7",
          2906 => x"d3",
          2907 => x"ff",
          2908 => x"8d",
          2909 => x"aa",
          2910 => x"22",
          2911 => x"72",
          2912 => x"80",
          2913 => x"d7",
          2914 => x"d3",
          2915 => x"16",
          2916 => x"08",
          2917 => x"b6",
          2918 => x"22",
          2919 => x"72",
          2920 => x"fe",
          2921 => x"08",
          2922 => x"0c",
          2923 => x"09",
          2924 => x"38",
          2925 => x"10",
          2926 => x"98",
          2927 => x"98",
          2928 => x"70",
          2929 => x"17",
          2930 => x"05",
          2931 => x"ff",
          2932 => x"53",
          2933 => x"9c",
          2934 => x"81",
          2935 => x"0b",
          2936 => x"ff",
          2937 => x"0c",
          2938 => x"84",
          2939 => x"83",
          2940 => x"06",
          2941 => x"80",
          2942 => x"d6",
          2943 => x"d3",
          2944 => x"ff",
          2945 => x"72",
          2946 => x"81",
          2947 => x"38",
          2948 => x"74",
          2949 => x"3f",
          2950 => x"08",
          2951 => x"91",
          2952 => x"84",
          2953 => x"b2",
          2954 => x"f0",
          2955 => x"c8",
          2956 => x"ff",
          2957 => x"82",
          2958 => x"09",
          2959 => x"c8",
          2960 => x"51",
          2961 => x"91",
          2962 => x"84",
          2963 => x"d2",
          2964 => x"06",
          2965 => x"98",
          2966 => x"d9",
          2967 => x"c8",
          2968 => x"85",
          2969 => x"09",
          2970 => x"38",
          2971 => x"51",
          2972 => x"91",
          2973 => x"90",
          2974 => x"a0",
          2975 => x"b5",
          2976 => x"c8",
          2977 => x"0c",
          2978 => x"91",
          2979 => x"81",
          2980 => x"91",
          2981 => x"72",
          2982 => x"80",
          2983 => x"0c",
          2984 => x"91",
          2985 => x"8f",
          2986 => x"fb",
          2987 => x"54",
          2988 => x"80",
          2989 => x"73",
          2990 => x"af",
          2991 => x"70",
          2992 => x"71",
          2993 => x"38",
          2994 => x"86",
          2995 => x"52",
          2996 => x"09",
          2997 => x"38",
          2998 => x"51",
          2999 => x"91",
          3000 => x"81",
          3001 => x"83",
          3002 => x"80",
          3003 => x"2e",
          3004 => x"84",
          3005 => x"53",
          3006 => x"0c",
          3007 => x"d3",
          3008 => x"3d",
          3009 => x"3d",
          3010 => x"05",
          3011 => x"89",
          3012 => x"52",
          3013 => x"3f",
          3014 => x"08",
          3015 => x"80",
          3016 => x"c8",
          3017 => x"c4",
          3018 => x"c8",
          3019 => x"91",
          3020 => x"70",
          3021 => x"73",
          3022 => x"38",
          3023 => x"78",
          3024 => x"38",
          3025 => x"74",
          3026 => x"10",
          3027 => x"05",
          3028 => x"54",
          3029 => x"80",
          3030 => x"80",
          3031 => x"70",
          3032 => x"51",
          3033 => x"91",
          3034 => x"54",
          3035 => x"c8",
          3036 => x"0d",
          3037 => x"0d",
          3038 => x"05",
          3039 => x"33",
          3040 => x"55",
          3041 => x"84",
          3042 => x"bf",
          3043 => x"98",
          3044 => x"53",
          3045 => x"05",
          3046 => x"c3",
          3047 => x"c8",
          3048 => x"d3",
          3049 => x"c5",
          3050 => x"68",
          3051 => x"d4",
          3052 => x"db",
          3053 => x"c8",
          3054 => x"d3",
          3055 => x"38",
          3056 => x"05",
          3057 => x"2b",
          3058 => x"80",
          3059 => x"86",
          3060 => x"06",
          3061 => x"2e",
          3062 => x"75",
          3063 => x"38",
          3064 => x"09",
          3065 => x"38",
          3066 => x"05",
          3067 => x"3f",
          3068 => x"08",
          3069 => x"07",
          3070 => x"02",
          3071 => x"91",
          3072 => x"80",
          3073 => x"87",
          3074 => x"76",
          3075 => x"81",
          3076 => x"74",
          3077 => x"38",
          3078 => x"83",
          3079 => x"83",
          3080 => x"06",
          3081 => x"80",
          3082 => x"38",
          3083 => x"51",
          3084 => x"91",
          3085 => x"59",
          3086 => x"0a",
          3087 => x"05",
          3088 => x"3f",
          3089 => x"0b",
          3090 => x"75",
          3091 => x"7a",
          3092 => x"3f",
          3093 => x"9c",
          3094 => x"a0",
          3095 => x"81",
          3096 => x"34",
          3097 => x"80",
          3098 => x"b0",
          3099 => x"55",
          3100 => x"3d",
          3101 => x"51",
          3102 => x"3f",
          3103 => x"08",
          3104 => x"c8",
          3105 => x"38",
          3106 => x"51",
          3107 => x"91",
          3108 => x"7b",
          3109 => x"12",
          3110 => x"b6",
          3111 => x"cd",
          3112 => x"05",
          3113 => x"2a",
          3114 => x"51",
          3115 => x"80",
          3116 => x"84",
          3117 => x"76",
          3118 => x"81",
          3119 => x"74",
          3120 => x"38",
          3121 => x"33",
          3122 => x"74",
          3123 => x"38",
          3124 => x"82",
          3125 => x"83",
          3126 => x"06",
          3127 => x"80",
          3128 => x"76",
          3129 => x"57",
          3130 => x"08",
          3131 => x"63",
          3132 => x"55",
          3133 => x"38",
          3134 => x"51",
          3135 => x"91",
          3136 => x"88",
          3137 => x"9c",
          3138 => x"a9",
          3139 => x"c8",
          3140 => x"0c",
          3141 => x"86",
          3142 => x"19",
          3143 => x"19",
          3144 => x"19",
          3145 => x"19",
          3146 => x"19",
          3147 => x"53",
          3148 => x"18",
          3149 => x"3f",
          3150 => x"70",
          3151 => x"55",
          3152 => x"81",
          3153 => x"18",
          3154 => x"81",
          3155 => x"18",
          3156 => x"0c",
          3157 => x"22",
          3158 => x"88",
          3159 => x"1c",
          3160 => x"5c",
          3161 => x"39",
          3162 => x"51",
          3163 => x"91",
          3164 => x"57",
          3165 => x"08",
          3166 => x"38",
          3167 => x"ff",
          3168 => x"06",
          3169 => x"56",
          3170 => x"59",
          3171 => x"77",
          3172 => x"70",
          3173 => x"06",
          3174 => x"74",
          3175 => x"98",
          3176 => x"80",
          3177 => x"83",
          3178 => x"74",
          3179 => x"38",
          3180 => x"51",
          3181 => x"91",
          3182 => x"85",
          3183 => x"a8",
          3184 => x"2a",
          3185 => x"08",
          3186 => x"1a",
          3187 => x"54",
          3188 => x"18",
          3189 => x"11",
          3190 => x"ca",
          3191 => x"d3",
          3192 => x"2e",
          3193 => x"56",
          3194 => x"84",
          3195 => x"0c",
          3196 => x"91",
          3197 => x"97",
          3198 => x"f3",
          3199 => x"62",
          3200 => x"5f",
          3201 => x"7d",
          3202 => x"fc",
          3203 => x"51",
          3204 => x"91",
          3205 => x"55",
          3206 => x"08",
          3207 => x"17",
          3208 => x"80",
          3209 => x"74",
          3210 => x"39",
          3211 => x"81",
          3212 => x"56",
          3213 => x"83",
          3214 => x"39",
          3215 => x"18",
          3216 => x"83",
          3217 => x"0b",
          3218 => x"81",
          3219 => x"39",
          3220 => x"18",
          3221 => x"83",
          3222 => x"0b",
          3223 => x"81",
          3224 => x"39",
          3225 => x"18",
          3226 => x"82",
          3227 => x"0b",
          3228 => x"81",
          3229 => x"39",
          3230 => x"94",
          3231 => x"55",
          3232 => x"83",
          3233 => x"78",
          3234 => x"cb",
          3235 => x"08",
          3236 => x"06",
          3237 => x"82",
          3238 => x"8a",
          3239 => x"05",
          3240 => x"06",
          3241 => x"a8",
          3242 => x"38",
          3243 => x"55",
          3244 => x"17",
          3245 => x"51",
          3246 => x"91",
          3247 => x"55",
          3248 => x"fe",
          3249 => x"ff",
          3250 => x"38",
          3251 => x"0c",
          3252 => x"52",
          3253 => x"e8",
          3254 => x"c8",
          3255 => x"fe",
          3256 => x"d3",
          3257 => x"79",
          3258 => x"58",
          3259 => x"80",
          3260 => x"1b",
          3261 => x"22",
          3262 => x"74",
          3263 => x"38",
          3264 => x"5a",
          3265 => x"53",
          3266 => x"81",
          3267 => x"55",
          3268 => x"91",
          3269 => x"fe",
          3270 => x"17",
          3271 => x"2b",
          3272 => x"80",
          3273 => x"9c",
          3274 => x"31",
          3275 => x"27",
          3276 => x"80",
          3277 => x"52",
          3278 => x"29",
          3279 => x"eb",
          3280 => x"2b",
          3281 => x"39",
          3282 => x"78",
          3283 => x"38",
          3284 => x"70",
          3285 => x"56",
          3286 => x"a5",
          3287 => x"9c",
          3288 => x"a8",
          3289 => x"81",
          3290 => x"55",
          3291 => x"91",
          3292 => x"fd",
          3293 => x"17",
          3294 => x"06",
          3295 => x"18",
          3296 => x"77",
          3297 => x"52",
          3298 => x"33",
          3299 => x"f1",
          3300 => x"c8",
          3301 => x"38",
          3302 => x"0c",
          3303 => x"83",
          3304 => x"80",
          3305 => x"55",
          3306 => x"83",
          3307 => x"75",
          3308 => x"08",
          3309 => x"17",
          3310 => x"7b",
          3311 => x"3f",
          3312 => x"7d",
          3313 => x"0c",
          3314 => x"19",
          3315 => x"1a",
          3316 => x"78",
          3317 => x"80",
          3318 => x"d3",
          3319 => x"3d",
          3320 => x"3d",
          3321 => x"64",
          3322 => x"5a",
          3323 => x"0c",
          3324 => x"05",
          3325 => x"f5",
          3326 => x"d3",
          3327 => x"91",
          3328 => x"8a",
          3329 => x"33",
          3330 => x"2e",
          3331 => x"56",
          3332 => x"90",
          3333 => x"81",
          3334 => x"06",
          3335 => x"87",
          3336 => x"2e",
          3337 => x"bd",
          3338 => x"91",
          3339 => x"56",
          3340 => x"81",
          3341 => x"34",
          3342 => x"d8",
          3343 => x"91",
          3344 => x"56",
          3345 => x"82",
          3346 => x"34",
          3347 => x"c4",
          3348 => x"91",
          3349 => x"56",
          3350 => x"81",
          3351 => x"34",
          3352 => x"b0",
          3353 => x"08",
          3354 => x"94",
          3355 => x"86",
          3356 => x"08",
          3357 => x"80",
          3358 => x"38",
          3359 => x"70",
          3360 => x"56",
          3361 => x"a8",
          3362 => x"11",
          3363 => x"77",
          3364 => x"5c",
          3365 => x"c6",
          3366 => x"38",
          3367 => x"55",
          3368 => x"7a",
          3369 => x"d4",
          3370 => x"d3",
          3371 => x"8f",
          3372 => x"08",
          3373 => x"d4",
          3374 => x"d3",
          3375 => x"74",
          3376 => x"c3",
          3377 => x"2e",
          3378 => x"74",
          3379 => x"e3",
          3380 => x"18",
          3381 => x"08",
          3382 => x"88",
          3383 => x"17",
          3384 => x"2b",
          3385 => x"80",
          3386 => x"81",
          3387 => x"08",
          3388 => x"52",
          3389 => x"33",
          3390 => x"de",
          3391 => x"c8",
          3392 => x"38",
          3393 => x"80",
          3394 => x"74",
          3395 => x"98",
          3396 => x"7d",
          3397 => x"3f",
          3398 => x"08",
          3399 => x"a7",
          3400 => x"c8",
          3401 => x"89",
          3402 => x"79",
          3403 => x"d5",
          3404 => x"7e",
          3405 => x"51",
          3406 => x"76",
          3407 => x"74",
          3408 => x"79",
          3409 => x"7b",
          3410 => x"11",
          3411 => x"c5",
          3412 => x"d3",
          3413 => x"f9",
          3414 => x"08",
          3415 => x"74",
          3416 => x"38",
          3417 => x"74",
          3418 => x"1c",
          3419 => x"51",
          3420 => x"90",
          3421 => x"ff",
          3422 => x"90",
          3423 => x"89",
          3424 => x"db",
          3425 => x"08",
          3426 => x"38",
          3427 => x"8c",
          3428 => x"98",
          3429 => x"77",
          3430 => x"52",
          3431 => x"33",
          3432 => x"dd",
          3433 => x"c8",
          3434 => x"38",
          3435 => x"0c",
          3436 => x"83",
          3437 => x"80",
          3438 => x"55",
          3439 => x"83",
          3440 => x"75",
          3441 => x"94",
          3442 => x"ff",
          3443 => x"05",
          3444 => x"3f",
          3445 => x"ff",
          3446 => x"74",
          3447 => x"78",
          3448 => x"08",
          3449 => x"76",
          3450 => x"08",
          3451 => x"1b",
          3452 => x"08",
          3453 => x"59",
          3454 => x"83",
          3455 => x"74",
          3456 => x"78",
          3457 => x"90",
          3458 => x"c0",
          3459 => x"90",
          3460 => x"56",
          3461 => x"c8",
          3462 => x"0d",
          3463 => x"0d",
          3464 => x"fc",
          3465 => x"52",
          3466 => x"3f",
          3467 => x"08",
          3468 => x"c8",
          3469 => x"38",
          3470 => x"70",
          3471 => x"81",
          3472 => x"56",
          3473 => x"81",
          3474 => x"98",
          3475 => x"80",
          3476 => x"81",
          3477 => x"08",
          3478 => x"52",
          3479 => x"33",
          3480 => x"f6",
          3481 => x"91",
          3482 => x"80",
          3483 => x"18",
          3484 => x"06",
          3485 => x"19",
          3486 => x"08",
          3487 => x"c8",
          3488 => x"d3",
          3489 => x"91",
          3490 => x"80",
          3491 => x"18",
          3492 => x"33",
          3493 => x"56",
          3494 => x"34",
          3495 => x"53",
          3496 => x"08",
          3497 => x"3f",
          3498 => x"52",
          3499 => x"c5",
          3500 => x"88",
          3501 => x"96",
          3502 => x"c0",
          3503 => x"92",
          3504 => x"9a",
          3505 => x"81",
          3506 => x"34",
          3507 => x"c1",
          3508 => x"c8",
          3509 => x"33",
          3510 => x"56",
          3511 => x"19",
          3512 => x"74",
          3513 => x"0c",
          3514 => x"04",
          3515 => x"76",
          3516 => x"fe",
          3517 => x"d3",
          3518 => x"91",
          3519 => x"9c",
          3520 => x"fc",
          3521 => x"51",
          3522 => x"91",
          3523 => x"53",
          3524 => x"08",
          3525 => x"d3",
          3526 => x"0c",
          3527 => x"c8",
          3528 => x"0d",
          3529 => x"0d",
          3530 => x"e4",
          3531 => x"53",
          3532 => x"d3",
          3533 => x"8b",
          3534 => x"c8",
          3535 => x"f8",
          3536 => x"72",
          3537 => x"0c",
          3538 => x"04",
          3539 => x"80",
          3540 => x"d0",
          3541 => x"3d",
          3542 => x"3f",
          3543 => x"08",
          3544 => x"c8",
          3545 => x"38",
          3546 => x"52",
          3547 => x"05",
          3548 => x"3f",
          3549 => x"08",
          3550 => x"c8",
          3551 => x"02",
          3552 => x"33",
          3553 => x"55",
          3554 => x"25",
          3555 => x"7a",
          3556 => x"54",
          3557 => x"a2",
          3558 => x"84",
          3559 => x"06",
          3560 => x"73",
          3561 => x"38",
          3562 => x"70",
          3563 => x"b8",
          3564 => x"c8",
          3565 => x"0c",
          3566 => x"55",
          3567 => x"09",
          3568 => x"38",
          3569 => x"91",
          3570 => x"93",
          3571 => x"e1",
          3572 => x"3d",
          3573 => x"08",
          3574 => x"7a",
          3575 => x"a1",
          3576 => x"05",
          3577 => x"51",
          3578 => x"91",
          3579 => x"57",
          3580 => x"08",
          3581 => x"7e",
          3582 => x"94",
          3583 => x"55",
          3584 => x"74",
          3585 => x"f9",
          3586 => x"70",
          3587 => x"5e",
          3588 => x"7a",
          3589 => x"3f",
          3590 => x"08",
          3591 => x"c8",
          3592 => x"38",
          3593 => x"51",
          3594 => x"91",
          3595 => x"57",
          3596 => x"08",
          3597 => x"6c",
          3598 => x"d6",
          3599 => x"d3",
          3600 => x"76",
          3601 => x"d1",
          3602 => x"d3",
          3603 => x"91",
          3604 => x"81",
          3605 => x"54",
          3606 => x"51",
          3607 => x"91",
          3608 => x"57",
          3609 => x"08",
          3610 => x"52",
          3611 => x"f8",
          3612 => x"c8",
          3613 => x"95",
          3614 => x"73",
          3615 => x"3f",
          3616 => x"08",
          3617 => x"c8",
          3618 => x"cc",
          3619 => x"2e",
          3620 => x"83",
          3621 => x"76",
          3622 => x"a1",
          3623 => x"11",
          3624 => x"51",
          3625 => x"76",
          3626 => x"79",
          3627 => x"33",
          3628 => x"55",
          3629 => x"2e",
          3630 => x"16",
          3631 => x"11",
          3632 => x"56",
          3633 => x"81",
          3634 => x"74",
          3635 => x"91",
          3636 => x"75",
          3637 => x"38",
          3638 => x"19",
          3639 => x"11",
          3640 => x"1b",
          3641 => x"59",
          3642 => x"75",
          3643 => x"38",
          3644 => x"3d",
          3645 => x"59",
          3646 => x"67",
          3647 => x"91",
          3648 => x"85",
          3649 => x"2e",
          3650 => x"8c",
          3651 => x"a3",
          3652 => x"55",
          3653 => x"34",
          3654 => x"d3",
          3655 => x"10",
          3656 => x"e8",
          3657 => x"70",
          3658 => x"57",
          3659 => x"73",
          3660 => x"38",
          3661 => x"16",
          3662 => x"55",
          3663 => x"38",
          3664 => x"73",
          3665 => x"38",
          3666 => x"76",
          3667 => x"77",
          3668 => x"33",
          3669 => x"05",
          3670 => x"18",
          3671 => x"26",
          3672 => x"7a",
          3673 => x"5c",
          3674 => x"58",
          3675 => x"91",
          3676 => x"38",
          3677 => x"19",
          3678 => x"54",
          3679 => x"70",
          3680 => x"34",
          3681 => x"ec",
          3682 => x"34",
          3683 => x"c8",
          3684 => x"0d",
          3685 => x"0d",
          3686 => x"3d",
          3687 => x"71",
          3688 => x"ea",
          3689 => x"d3",
          3690 => x"91",
          3691 => x"8a",
          3692 => x"33",
          3693 => x"2e",
          3694 => x"55",
          3695 => x"8c",
          3696 => x"27",
          3697 => x"17",
          3698 => x"2a",
          3699 => x"51",
          3700 => x"85",
          3701 => x"08",
          3702 => x"08",
          3703 => x"94",
          3704 => x"77",
          3705 => x"b3",
          3706 => x"11",
          3707 => x"2b",
          3708 => x"75",
          3709 => x"38",
          3710 => x"18",
          3711 => x"b9",
          3712 => x"c8",
          3713 => x"7a",
          3714 => x"57",
          3715 => x"a9",
          3716 => x"c8",
          3717 => x"95",
          3718 => x"76",
          3719 => x"0c",
          3720 => x"08",
          3721 => x"08",
          3722 => x"c9",
          3723 => x"08",
          3724 => x"38",
          3725 => x"51",
          3726 => x"91",
          3727 => x"56",
          3728 => x"08",
          3729 => x"81",
          3730 => x"82",
          3731 => x"34",
          3732 => x"e3",
          3733 => x"c8",
          3734 => x"09",
          3735 => x"38",
          3736 => x"18",
          3737 => x"82",
          3738 => x"d3",
          3739 => x"18",
          3740 => x"18",
          3741 => x"2e",
          3742 => x"78",
          3743 => x"ea",
          3744 => x"31",
          3745 => x"1a",
          3746 => x"90",
          3747 => x"81",
          3748 => x"06",
          3749 => x"58",
          3750 => x"9a",
          3751 => x"76",
          3752 => x"3f",
          3753 => x"08",
          3754 => x"c8",
          3755 => x"91",
          3756 => x"58",
          3757 => x"52",
          3758 => x"ae",
          3759 => x"c8",
          3760 => x"ff",
          3761 => x"38",
          3762 => x"8a",
          3763 => x"98",
          3764 => x"26",
          3765 => x"0b",
          3766 => x"82",
          3767 => x"39",
          3768 => x"0c",
          3769 => x"ff",
          3770 => x"17",
          3771 => x"18",
          3772 => x"ff",
          3773 => x"80",
          3774 => x"75",
          3775 => x"c1",
          3776 => x"d3",
          3777 => x"38",
          3778 => x"18",
          3779 => x"81",
          3780 => x"89",
          3781 => x"c8",
          3782 => x"8c",
          3783 => x"18",
          3784 => x"38",
          3785 => x"8c",
          3786 => x"17",
          3787 => x"07",
          3788 => x"18",
          3789 => x"08",
          3790 => x"55",
          3791 => x"80",
          3792 => x"17",
          3793 => x"80",
          3794 => x"17",
          3795 => x"2b",
          3796 => x"80",
          3797 => x"81",
          3798 => x"08",
          3799 => x"52",
          3800 => x"33",
          3801 => x"b8",
          3802 => x"d3",
          3803 => x"2e",
          3804 => x"0b",
          3805 => x"81",
          3806 => x"90",
          3807 => x"ff",
          3808 => x"90",
          3809 => x"54",
          3810 => x"17",
          3811 => x"11",
          3812 => x"ff",
          3813 => x"91",
          3814 => x"80",
          3815 => x"81",
          3816 => x"34",
          3817 => x"39",
          3818 => x"18",
          3819 => x"87",
          3820 => x"18",
          3821 => x"74",
          3822 => x"0c",
          3823 => x"04",
          3824 => x"79",
          3825 => x"75",
          3826 => x"8f",
          3827 => x"89",
          3828 => x"52",
          3829 => x"05",
          3830 => x"3f",
          3831 => x"08",
          3832 => x"c8",
          3833 => x"38",
          3834 => x"7a",
          3835 => x"d8",
          3836 => x"d3",
          3837 => x"91",
          3838 => x"80",
          3839 => x"16",
          3840 => x"2b",
          3841 => x"74",
          3842 => x"86",
          3843 => x"84",
          3844 => x"06",
          3845 => x"73",
          3846 => x"38",
          3847 => x"52",
          3848 => x"c4",
          3849 => x"c8",
          3850 => x"0c",
          3851 => x"55",
          3852 => x"77",
          3853 => x"22",
          3854 => x"74",
          3855 => x"c9",
          3856 => x"d3",
          3857 => x"74",
          3858 => x"81",
          3859 => x"85",
          3860 => x"2e",
          3861 => x"76",
          3862 => x"73",
          3863 => x"0c",
          3864 => x"04",
          3865 => x"76",
          3866 => x"05",
          3867 => x"54",
          3868 => x"91",
          3869 => x"53",
          3870 => x"08",
          3871 => x"d3",
          3872 => x"0c",
          3873 => x"c8",
          3874 => x"0d",
          3875 => x"0d",
          3876 => x"3d",
          3877 => x"71",
          3878 => x"e4",
          3879 => x"d3",
          3880 => x"91",
          3881 => x"80",
          3882 => x"92",
          3883 => x"c8",
          3884 => x"51",
          3885 => x"91",
          3886 => x"53",
          3887 => x"52",
          3888 => x"8b",
          3889 => x"c8",
          3890 => x"d3",
          3891 => x"2e",
          3892 => x"83",
          3893 => x"72",
          3894 => x"52",
          3895 => x"b4",
          3896 => x"73",
          3897 => x"3f",
          3898 => x"08",
          3899 => x"c8",
          3900 => x"09",
          3901 => x"38",
          3902 => x"91",
          3903 => x"87",
          3904 => x"ef",
          3905 => x"56",
          3906 => x"3d",
          3907 => x"3d",
          3908 => x"cb",
          3909 => x"c8",
          3910 => x"d3",
          3911 => x"38",
          3912 => x"51",
          3913 => x"91",
          3914 => x"55",
          3915 => x"08",
          3916 => x"80",
          3917 => x"70",
          3918 => x"57",
          3919 => x"85",
          3920 => x"90",
          3921 => x"2e",
          3922 => x"52",
          3923 => x"05",
          3924 => x"3f",
          3925 => x"c8",
          3926 => x"0d",
          3927 => x"0d",
          3928 => x"5a",
          3929 => x"3d",
          3930 => x"91",
          3931 => x"ef",
          3932 => x"c8",
          3933 => x"d3",
          3934 => x"84",
          3935 => x"0c",
          3936 => x"11",
          3937 => x"55",
          3938 => x"08",
          3939 => x"38",
          3940 => x"7a",
          3941 => x"39",
          3942 => x"cf",
          3943 => x"81",
          3944 => x"7b",
          3945 => x"56",
          3946 => x"2e",
          3947 => x"80",
          3948 => x"75",
          3949 => x"52",
          3950 => x"05",
          3951 => x"aa",
          3952 => x"c8",
          3953 => x"d0",
          3954 => x"c8",
          3955 => x"cd",
          3956 => x"c8",
          3957 => x"91",
          3958 => x"07",
          3959 => x"05",
          3960 => x"53",
          3961 => x"98",
          3962 => x"26",
          3963 => x"fb",
          3964 => x"11",
          3965 => x"08",
          3966 => x"80",
          3967 => x"38",
          3968 => x"18",
          3969 => x"ff",
          3970 => x"91",
          3971 => x"59",
          3972 => x"08",
          3973 => x"7a",
          3974 => x"54",
          3975 => x"09",
          3976 => x"38",
          3977 => x"05",
          3978 => x"f0",
          3979 => x"c8",
          3980 => x"ff",
          3981 => x"70",
          3982 => x"82",
          3983 => x"51",
          3984 => x"7a",
          3985 => x"51",
          3986 => x"3f",
          3987 => x"08",
          3988 => x"70",
          3989 => x"25",
          3990 => x"58",
          3991 => x"74",
          3992 => x"ff",
          3993 => x"75",
          3994 => x"76",
          3995 => x"77",
          3996 => x"54",
          3997 => x"33",
          3998 => x"55",
          3999 => x"34",
          4000 => x"c8",
          4001 => x"0d",
          4002 => x"0d",
          4003 => x"fc",
          4004 => x"52",
          4005 => x"3f",
          4006 => x"08",
          4007 => x"c8",
          4008 => x"91",
          4009 => x"76",
          4010 => x"38",
          4011 => x"dc",
          4012 => x"33",
          4013 => x"70",
          4014 => x"56",
          4015 => x"74",
          4016 => x"c8",
          4017 => x"08",
          4018 => x"27",
          4019 => x"94",
          4020 => x"38",
          4021 => x"18",
          4022 => x"51",
          4023 => x"3f",
          4024 => x"08",
          4025 => x"88",
          4026 => x"ca",
          4027 => x"08",
          4028 => x"ff",
          4029 => x"91",
          4030 => x"91",
          4031 => x"ff",
          4032 => x"70",
          4033 => x"25",
          4034 => x"56",
          4035 => x"08",
          4036 => x"81",
          4037 => x"82",
          4038 => x"38",
          4039 => x"98",
          4040 => x"92",
          4041 => x"08",
          4042 => x"77",
          4043 => x"fe",
          4044 => x"c8",
          4045 => x"18",
          4046 => x"0c",
          4047 => x"80",
          4048 => x"74",
          4049 => x"76",
          4050 => x"98",
          4051 => x"80",
          4052 => x"81",
          4053 => x"08",
          4054 => x"52",
          4055 => x"33",
          4056 => x"b0",
          4057 => x"d3",
          4058 => x"2e",
          4059 => x"57",
          4060 => x"18",
          4061 => x"06",
          4062 => x"19",
          4063 => x"2e",
          4064 => x"91",
          4065 => x"56",
          4066 => x"56",
          4067 => x"c8",
          4068 => x"0d",
          4069 => x"0d",
          4070 => x"51",
          4071 => x"3f",
          4072 => x"3d",
          4073 => x"52",
          4074 => x"d6",
          4075 => x"d3",
          4076 => x"91",
          4077 => x"82",
          4078 => x"bb",
          4079 => x"96",
          4080 => x"44",
          4081 => x"3d",
          4082 => x"d0",
          4083 => x"d3",
          4084 => x"bb",
          4085 => x"ff",
          4086 => x"75",
          4087 => x"02",
          4088 => x"33",
          4089 => x"70",
          4090 => x"55",
          4091 => x"2e",
          4092 => x"56",
          4093 => x"38",
          4094 => x"51",
          4095 => x"3f",
          4096 => x"05",
          4097 => x"2b",
          4098 => x"80",
          4099 => x"86",
          4100 => x"02",
          4101 => x"33",
          4102 => x"73",
          4103 => x"38",
          4104 => x"81",
          4105 => x"52",
          4106 => x"bc",
          4107 => x"c8",
          4108 => x"05",
          4109 => x"33",
          4110 => x"70",
          4111 => x"56",
          4112 => x"80",
          4113 => x"38",
          4114 => x"51",
          4115 => x"3f",
          4116 => x"56",
          4117 => x"77",
          4118 => x"38",
          4119 => x"51",
          4120 => x"3f",
          4121 => x"5b",
          4122 => x"51",
          4123 => x"3f",
          4124 => x"3d",
          4125 => x"c1",
          4126 => x"d3",
          4127 => x"91",
          4128 => x"81",
          4129 => x"d3",
          4130 => x"73",
          4131 => x"3f",
          4132 => x"08",
          4133 => x"c8",
          4134 => x"87",
          4135 => x"32",
          4136 => x"72",
          4137 => x"78",
          4138 => x"54",
          4139 => x"38",
          4140 => x"51",
          4141 => x"3f",
          4142 => x"05",
          4143 => x"3f",
          4144 => x"08",
          4145 => x"08",
          4146 => x"d3",
          4147 => x"80",
          4148 => x"70",
          4149 => x"2a",
          4150 => x"57",
          4151 => x"74",
          4152 => x"38",
          4153 => x"51",
          4154 => x"3f",
          4155 => x"52",
          4156 => x"05",
          4157 => x"b6",
          4158 => x"c8",
          4159 => x"8c",
          4160 => x"ff",
          4161 => x"91",
          4162 => x"56",
          4163 => x"51",
          4164 => x"3f",
          4165 => x"c8",
          4166 => x"0d",
          4167 => x"0d",
          4168 => x"3d",
          4169 => x"99",
          4170 => x"b3",
          4171 => x"c8",
          4172 => x"d3",
          4173 => x"b5",
          4174 => x"68",
          4175 => x"d4",
          4176 => x"cb",
          4177 => x"c8",
          4178 => x"d3",
          4179 => x"38",
          4180 => x"84",
          4181 => x"06",
          4182 => x"02",
          4183 => x"33",
          4184 => x"70",
          4185 => x"55",
          4186 => x"2e",
          4187 => x"55",
          4188 => x"09",
          4189 => x"f5",
          4190 => x"80",
          4191 => x"c4",
          4192 => x"ba",
          4193 => x"d3",
          4194 => x"80",
          4195 => x"c8",
          4196 => x"09",
          4197 => x"38",
          4198 => x"81",
          4199 => x"06",
          4200 => x"55",
          4201 => x"09",
          4202 => x"38",
          4203 => x"88",
          4204 => x"74",
          4205 => x"75",
          4206 => x"ff",
          4207 => x"91",
          4208 => x"55",
          4209 => x"08",
          4210 => x"8b",
          4211 => x"b4",
          4212 => x"af",
          4213 => x"54",
          4214 => x"15",
          4215 => x"90",
          4216 => x"34",
          4217 => x"ca",
          4218 => x"af",
          4219 => x"53",
          4220 => x"77",
          4221 => x"3f",
          4222 => x"18",
          4223 => x"18",
          4224 => x"a7",
          4225 => x"ae",
          4226 => x"15",
          4227 => x"80",
          4228 => x"77",
          4229 => x"3f",
          4230 => x"0b",
          4231 => x"98",
          4232 => x"51",
          4233 => x"91",
          4234 => x"55",
          4235 => x"08",
          4236 => x"52",
          4237 => x"51",
          4238 => x"3f",
          4239 => x"52",
          4240 => x"dd",
          4241 => x"90",
          4242 => x"34",
          4243 => x"0b",
          4244 => x"77",
          4245 => x"b9",
          4246 => x"c8",
          4247 => x"39",
          4248 => x"52",
          4249 => x"05",
          4250 => x"c2",
          4251 => x"d3",
          4252 => x"3d",
          4253 => x"3d",
          4254 => x"84",
          4255 => x"c8",
          4256 => x"a7",
          4257 => x"05",
          4258 => x"51",
          4259 => x"91",
          4260 => x"55",
          4261 => x"08",
          4262 => x"77",
          4263 => x"08",
          4264 => x"d4",
          4265 => x"e7",
          4266 => x"c8",
          4267 => x"d3",
          4268 => x"bd",
          4269 => x"97",
          4270 => x"a0",
          4271 => x"80",
          4272 => x"86",
          4273 => x"a9",
          4274 => x"a3",
          4275 => x"a7",
          4276 => x"05",
          4277 => x"d3",
          4278 => x"a7",
          4279 => x"52",
          4280 => x"52",
          4281 => x"c3",
          4282 => x"08",
          4283 => x"ca",
          4284 => x"d3",
          4285 => x"91",
          4286 => x"94",
          4287 => x"2e",
          4288 => x"8a",
          4289 => x"64",
          4290 => x"2e",
          4291 => x"55",
          4292 => x"09",
          4293 => x"b8",
          4294 => x"ff",
          4295 => x"c3",
          4296 => x"d3",
          4297 => x"91",
          4298 => x"81",
          4299 => x"56",
          4300 => x"3d",
          4301 => x"52",
          4302 => x"ff",
          4303 => x"02",
          4304 => x"8b",
          4305 => x"16",
          4306 => x"2a",
          4307 => x"51",
          4308 => x"89",
          4309 => x"07",
          4310 => x"17",
          4311 => x"81",
          4312 => x"34",
          4313 => x"70",
          4314 => x"81",
          4315 => x"57",
          4316 => x"80",
          4317 => x"63",
          4318 => x"38",
          4319 => x"51",
          4320 => x"3f",
          4321 => x"08",
          4322 => x"ff",
          4323 => x"82",
          4324 => x"c8",
          4325 => x"b8",
          4326 => x"c8",
          4327 => x"51",
          4328 => x"3f",
          4329 => x"08",
          4330 => x"57",
          4331 => x"c8",
          4332 => x"81",
          4333 => x"73",
          4334 => x"81",
          4335 => x"62",
          4336 => x"77",
          4337 => x"d9",
          4338 => x"81",
          4339 => x"34",
          4340 => x"a7",
          4341 => x"51",
          4342 => x"91",
          4343 => x"55",
          4344 => x"08",
          4345 => x"51",
          4346 => x"3f",
          4347 => x"08",
          4348 => x"d3",
          4349 => x"3d",
          4350 => x"3d",
          4351 => x"db",
          4352 => x"84",
          4353 => x"05",
          4354 => x"82",
          4355 => x"d0",
          4356 => x"3d",
          4357 => x"3f",
          4358 => x"08",
          4359 => x"c8",
          4360 => x"38",
          4361 => x"52",
          4362 => x"05",
          4363 => x"3f",
          4364 => x"08",
          4365 => x"c8",
          4366 => x"02",
          4367 => x"33",
          4368 => x"54",
          4369 => x"83",
          4370 => x"74",
          4371 => x"a7",
          4372 => x"09",
          4373 => x"71",
          4374 => x"06",
          4375 => x"55",
          4376 => x"15",
          4377 => x"81",
          4378 => x"34",
          4379 => x"ad",
          4380 => x"d3",
          4381 => x"74",
          4382 => x"0c",
          4383 => x"04",
          4384 => x"65",
          4385 => x"94",
          4386 => x"52",
          4387 => x"cc",
          4388 => x"d3",
          4389 => x"91",
          4390 => x"80",
          4391 => x"59",
          4392 => x"3d",
          4393 => x"c6",
          4394 => x"d3",
          4395 => x"91",
          4396 => x"bc",
          4397 => x"cb",
          4398 => x"a0",
          4399 => x"80",
          4400 => x"86",
          4401 => x"38",
          4402 => x"84",
          4403 => x"90",
          4404 => x"54",
          4405 => x"96",
          4406 => x"a9",
          4407 => x"54",
          4408 => x"15",
          4409 => x"ff",
          4410 => x"91",
          4411 => x"55",
          4412 => x"c8",
          4413 => x"0d",
          4414 => x"0d",
          4415 => x"59",
          4416 => x"3d",
          4417 => x"99",
          4418 => x"d3",
          4419 => x"c8",
          4420 => x"c8",
          4421 => x"91",
          4422 => x"07",
          4423 => x"30",
          4424 => x"9f",
          4425 => x"52",
          4426 => x"56",
          4427 => x"80",
          4428 => x"5d",
          4429 => x"52",
          4430 => x"52",
          4431 => x"bb",
          4432 => x"c8",
          4433 => x"d3",
          4434 => x"ce",
          4435 => x"73",
          4436 => x"fb",
          4437 => x"c8",
          4438 => x"d3",
          4439 => x"38",
          4440 => x"08",
          4441 => x"08",
          4442 => x"58",
          4443 => x"18",
          4444 => x"58",
          4445 => x"74",
          4446 => x"58",
          4447 => x"ec",
          4448 => x"54",
          4449 => x"77",
          4450 => x"38",
          4451 => x"11",
          4452 => x"55",
          4453 => x"2e",
          4454 => x"84",
          4455 => x"06",
          4456 => x"79",
          4457 => x"75",
          4458 => x"07",
          4459 => x"30",
          4460 => x"9f",
          4461 => x"52",
          4462 => x"74",
          4463 => x"38",
          4464 => x"08",
          4465 => x"aa",
          4466 => x"d3",
          4467 => x"91",
          4468 => x"a7",
          4469 => x"33",
          4470 => x"c3",
          4471 => x"2e",
          4472 => x"e4",
          4473 => x"2e",
          4474 => x"58",
          4475 => x"05",
          4476 => x"c1",
          4477 => x"c8",
          4478 => x"75",
          4479 => x"0c",
          4480 => x"04",
          4481 => x"82",
          4482 => x"ff",
          4483 => x"9b",
          4484 => x"cb",
          4485 => x"c8",
          4486 => x"d3",
          4487 => x"c8",
          4488 => x"a0",
          4489 => x"ff",
          4490 => x"ff",
          4491 => x"80",
          4492 => x"33",
          4493 => x"57",
          4494 => x"81",
          4495 => x"33",
          4496 => x"4c",
          4497 => x"06",
          4498 => x"a7",
          4499 => x"d3",
          4500 => x"2e",
          4501 => x"70",
          4502 => x"51",
          4503 => x"f2",
          4504 => x"c8",
          4505 => x"8d",
          4506 => x"2b",
          4507 => x"81",
          4508 => x"83",
          4509 => x"ff",
          4510 => x"73",
          4511 => x"38",
          4512 => x"83",
          4513 => x"57",
          4514 => x"76",
          4515 => x"91",
          4516 => x"33",
          4517 => x"2e",
          4518 => x"52",
          4519 => x"51",
          4520 => x"3f",
          4521 => x"08",
          4522 => x"ff",
          4523 => x"38",
          4524 => x"88",
          4525 => x"8a",
          4526 => x"38",
          4527 => x"a8",
          4528 => x"76",
          4529 => x"9a",
          4530 => x"ff",
          4531 => x"88",
          4532 => x"73",
          4533 => x"17",
          4534 => x"77",
          4535 => x"05",
          4536 => x"34",
          4537 => x"70",
          4538 => x"57",
          4539 => x"fe",
          4540 => x"3d",
          4541 => x"55",
          4542 => x"2e",
          4543 => x"76",
          4544 => x"38",
          4545 => x"70",
          4546 => x"33",
          4547 => x"54",
          4548 => x"09",
          4549 => x"38",
          4550 => x"76",
          4551 => x"38",
          4552 => x"33",
          4553 => x"a0",
          4554 => x"77",
          4555 => x"80",
          4556 => x"70",
          4557 => x"b3",
          4558 => x"d3",
          4559 => x"91",
          4560 => x"81",
          4561 => x"52",
          4562 => x"b9",
          4563 => x"d3",
          4564 => x"91",
          4565 => x"b0",
          4566 => x"2e",
          4567 => x"53",
          4568 => x"bc",
          4569 => x"51",
          4570 => x"3f",
          4571 => x"54",
          4572 => x"77",
          4573 => x"83",
          4574 => x"51",
          4575 => x"3f",
          4576 => x"08",
          4577 => x"39",
          4578 => x"08",
          4579 => x"81",
          4580 => x"38",
          4581 => x"74",
          4582 => x"38",
          4583 => x"3d",
          4584 => x"ff",
          4585 => x"91",
          4586 => x"54",
          4587 => x"08",
          4588 => x"53",
          4589 => x"08",
          4590 => x"ff",
          4591 => x"65",
          4592 => x"8b",
          4593 => x"53",
          4594 => x"bc",
          4595 => x"51",
          4596 => x"3f",
          4597 => x"0b",
          4598 => x"77",
          4599 => x"b1",
          4600 => x"c8",
          4601 => x"55",
          4602 => x"c8",
          4603 => x"0d",
          4604 => x"0d",
          4605 => x"88",
          4606 => x"05",
          4607 => x"fc",
          4608 => x"54",
          4609 => x"cd",
          4610 => x"d3",
          4611 => x"91",
          4612 => x"8a",
          4613 => x"33",
          4614 => x"2e",
          4615 => x"54",
          4616 => x"7a",
          4617 => x"38",
          4618 => x"90",
          4619 => x"33",
          4620 => x"70",
          4621 => x"55",
          4622 => x"38",
          4623 => x"99",
          4624 => x"81",
          4625 => x"57",
          4626 => x"7f",
          4627 => x"70",
          4628 => x"55",
          4629 => x"51",
          4630 => x"dd",
          4631 => x"7b",
          4632 => x"70",
          4633 => x"2a",
          4634 => x"08",
          4635 => x"11",
          4636 => x"40",
          4637 => x"5f",
          4638 => x"88",
          4639 => x"08",
          4640 => x"38",
          4641 => x"79",
          4642 => x"5a",
          4643 => x"51",
          4644 => x"3f",
          4645 => x"08",
          4646 => x"56",
          4647 => x"14",
          4648 => x"83",
          4649 => x"75",
          4650 => x"95",
          4651 => x"2e",
          4652 => x"75",
          4653 => x"1a",
          4654 => x"2e",
          4655 => x"39",
          4656 => x"5a",
          4657 => x"09",
          4658 => x"38",
          4659 => x"81",
          4660 => x"80",
          4661 => x"7c",
          4662 => x"7d",
          4663 => x"38",
          4664 => x"75",
          4665 => x"81",
          4666 => x"ff",
          4667 => x"74",
          4668 => x"ff",
          4669 => x"91",
          4670 => x"57",
          4671 => x"08",
          4672 => x"81",
          4673 => x"58",
          4674 => x"d4",
          4675 => x"ff",
          4676 => x"80",
          4677 => x"7f",
          4678 => x"54",
          4679 => x"b7",
          4680 => x"19",
          4681 => x"19",
          4682 => x"33",
          4683 => x"54",
          4684 => x"34",
          4685 => x"08",
          4686 => x"55",
          4687 => x"74",
          4688 => x"90",
          4689 => x"31",
          4690 => x"7f",
          4691 => x"81",
          4692 => x"73",
          4693 => x"76",
          4694 => x"d3",
          4695 => x"3d",
          4696 => x"3d",
          4697 => x"84",
          4698 => x"05",
          4699 => x"53",
          4700 => x"bf",
          4701 => x"d3",
          4702 => x"8b",
          4703 => x"91",
          4704 => x"24",
          4705 => x"91",
          4706 => x"10",
          4707 => x"e4",
          4708 => x"08",
          4709 => x"38",
          4710 => x"80",
          4711 => x"81",
          4712 => x"81",
          4713 => x"ff",
          4714 => x"91",
          4715 => x"81",
          4716 => x"81",
          4717 => x"83",
          4718 => x"9b",
          4719 => x"2a",
          4720 => x"51",
          4721 => x"74",
          4722 => x"98",
          4723 => x"53",
          4724 => x"51",
          4725 => x"3f",
          4726 => x"08",
          4727 => x"80",
          4728 => x"66",
          4729 => x"26",
          4730 => x"ff",
          4731 => x"55",
          4732 => x"83",
          4733 => x"84",
          4734 => x"80",
          4735 => x"7d",
          4736 => x"38",
          4737 => x"0a",
          4738 => x"ff",
          4739 => x"55",
          4740 => x"86",
          4741 => x"8b",
          4742 => x"52",
          4743 => x"f6",
          4744 => x"d3",
          4745 => x"7f",
          4746 => x"40",
          4747 => x"89",
          4748 => x"c8",
          4749 => x"d3",
          4750 => x"60",
          4751 => x"07",
          4752 => x"d3",
          4753 => x"70",
          4754 => x"08",
          4755 => x"72",
          4756 => x"51",
          4757 => x"91",
          4758 => x"fb",
          4759 => x"f8",
          4760 => x"52",
          4761 => x"9c",
          4762 => x"57",
          4763 => x"08",
          4764 => x"7c",
          4765 => x"81",
          4766 => x"80",
          4767 => x"2e",
          4768 => x"83",
          4769 => x"8e",
          4770 => x"26",
          4771 => x"65",
          4772 => x"8e",
          4773 => x"66",
          4774 => x"38",
          4775 => x"81",
          4776 => x"b3",
          4777 => x"2a",
          4778 => x"51",
          4779 => x"2e",
          4780 => x"87",
          4781 => x"82",
          4782 => x"7c",
          4783 => x"74",
          4784 => x"42",
          4785 => x"81",
          4786 => x"57",
          4787 => x"80",
          4788 => x"38",
          4789 => x"83",
          4790 => x"06",
          4791 => x"77",
          4792 => x"91",
          4793 => x"57",
          4794 => x"bd",
          4795 => x"22",
          4796 => x"59",
          4797 => x"9d",
          4798 => x"26",
          4799 => x"1b",
          4800 => x"10",
          4801 => x"51",
          4802 => x"74",
          4803 => x"38",
          4804 => x"ea",
          4805 => x"65",
          4806 => x"9d",
          4807 => x"c8",
          4808 => x"c8",
          4809 => x"1f",
          4810 => x"05",
          4811 => x"f4",
          4812 => x"d3",
          4813 => x"a0",
          4814 => x"fc",
          4815 => x"56",
          4816 => x"f0",
          4817 => x"81",
          4818 => x"57",
          4819 => x"77",
          4820 => x"8c",
          4821 => x"57",
          4822 => x"bd",
          4823 => x"22",
          4824 => x"59",
          4825 => x"9d",
          4826 => x"26",
          4827 => x"1b",
          4828 => x"10",
          4829 => x"51",
          4830 => x"74",
          4831 => x"38",
          4832 => x"ea",
          4833 => x"65",
          4834 => x"ad",
          4835 => x"c8",
          4836 => x"05",
          4837 => x"c8",
          4838 => x"26",
          4839 => x"0b",
          4840 => x"08",
          4841 => x"70",
          4842 => x"05",
          4843 => x"7d",
          4844 => x"ff",
          4845 => x"f3",
          4846 => x"d3",
          4847 => x"81",
          4848 => x"81",
          4849 => x"fe",
          4850 => x"91",
          4851 => x"83",
          4852 => x"43",
          4853 => x"11",
          4854 => x"11",
          4855 => x"30",
          4856 => x"73",
          4857 => x"59",
          4858 => x"83",
          4859 => x"06",
          4860 => x"1b",
          4861 => x"5b",
          4862 => x"1c",
          4863 => x"29",
          4864 => x"31",
          4865 => x"66",
          4866 => x"38",
          4867 => x"7c",
          4868 => x"70",
          4869 => x"56",
          4870 => x"3f",
          4871 => x"08",
          4872 => x"2e",
          4873 => x"9b",
          4874 => x"c8",
          4875 => x"f5",
          4876 => x"77",
          4877 => x"81",
          4878 => x"fd",
          4879 => x"57",
          4880 => x"61",
          4881 => x"81",
          4882 => x"38",
          4883 => x"76",
          4884 => x"77",
          4885 => x"19",
          4886 => x"c0",
          4887 => x"74",
          4888 => x"39",
          4889 => x"81",
          4890 => x"80",
          4891 => x"83",
          4892 => x"39",
          4893 => x"78",
          4894 => x"80",
          4895 => x"d4",
          4896 => x"86",
          4897 => x"9f",
          4898 => x"38",
          4899 => x"78",
          4900 => x"80",
          4901 => x"bc",
          4902 => x"86",
          4903 => x"55",
          4904 => x"09",
          4905 => x"38",
          4906 => x"9f",
          4907 => x"06",
          4908 => x"74",
          4909 => x"7d",
          4910 => x"7e",
          4911 => x"8f",
          4912 => x"91",
          4913 => x"7e",
          4914 => x"df",
          4915 => x"8b",
          4916 => x"99",
          4917 => x"7f",
          4918 => x"7a",
          4919 => x"06",
          4920 => x"51",
          4921 => x"3f",
          4922 => x"05",
          4923 => x"32",
          4924 => x"96",
          4925 => x"06",
          4926 => x"91",
          4927 => x"98",
          4928 => x"83",
          4929 => x"90",
          4930 => x"d6",
          4931 => x"93",
          4932 => x"98",
          4933 => x"39",
          4934 => x"1f",
          4935 => x"dc",
          4936 => x"95",
          4937 => x"52",
          4938 => x"ff",
          4939 => x"81",
          4940 => x"1f",
          4941 => x"a6",
          4942 => x"9c",
          4943 => x"98",
          4944 => x"83",
          4945 => x"06",
          4946 => x"82",
          4947 => x"52",
          4948 => x"51",
          4949 => x"3f",
          4950 => x"1f",
          4951 => x"9c",
          4952 => x"ac",
          4953 => x"98",
          4954 => x"52",
          4955 => x"ff",
          4956 => x"86",
          4957 => x"51",
          4958 => x"3f",
          4959 => x"80",
          4960 => x"a9",
          4961 => x"05",
          4962 => x"91",
          4963 => x"80",
          4964 => x"ff",
          4965 => x"b2",
          4966 => x"b2",
          4967 => x"1f",
          4968 => x"d8",
          4969 => x"ff",
          4970 => x"96",
          4971 => x"97",
          4972 => x"80",
          4973 => x"34",
          4974 => x"05",
          4975 => x"91",
          4976 => x"ab",
          4977 => x"97",
          4978 => x"d4",
          4979 => x"fe",
          4980 => x"97",
          4981 => x"54",
          4982 => x"52",
          4983 => x"93",
          4984 => x"57",
          4985 => x"08",
          4986 => x"61",
          4987 => x"81",
          4988 => x"38",
          4989 => x"86",
          4990 => x"52",
          4991 => x"93",
          4992 => x"53",
          4993 => x"51",
          4994 => x"3f",
          4995 => x"a4",
          4996 => x"51",
          4997 => x"3f",
          4998 => x"e4",
          4999 => x"e4",
          5000 => x"96",
          5001 => x"16",
          5002 => x"1f",
          5003 => x"cc",
          5004 => x"83",
          5005 => x"ff",
          5006 => x"82",
          5007 => x"83",
          5008 => x"ff",
          5009 => x"81",
          5010 => x"05",
          5011 => x"79",
          5012 => x"86",
          5013 => x"63",
          5014 => x"7e",
          5015 => x"ff",
          5016 => x"64",
          5017 => x"7e",
          5018 => x"e3",
          5019 => x"80",
          5020 => x"2e",
          5021 => x"9e",
          5022 => x"7e",
          5023 => x"fc",
          5024 => x"84",
          5025 => x"95",
          5026 => x"0a",
          5027 => x"51",
          5028 => x"3f",
          5029 => x"ff",
          5030 => x"61",
          5031 => x"38",
          5032 => x"52",
          5033 => x"95",
          5034 => x"55",
          5035 => x"61",
          5036 => x"74",
          5037 => x"75",
          5038 => x"79",
          5039 => x"9a",
          5040 => x"c8",
          5041 => x"38",
          5042 => x"52",
          5043 => x"95",
          5044 => x"16",
          5045 => x"56",
          5046 => x"38",
          5047 => x"7a",
          5048 => x"8d",
          5049 => x"61",
          5050 => x"38",
          5051 => x"57",
          5052 => x"83",
          5053 => x"76",
          5054 => x"7e",
          5055 => x"ff",
          5056 => x"91",
          5057 => x"81",
          5058 => x"16",
          5059 => x"56",
          5060 => x"38",
          5061 => x"83",
          5062 => x"86",
          5063 => x"ff",
          5064 => x"38",
          5065 => x"82",
          5066 => x"81",
          5067 => x"2a",
          5068 => x"77",
          5069 => x"7d",
          5070 => x"7e",
          5071 => x"8f",
          5072 => x"d5",
          5073 => x"1f",
          5074 => x"92",
          5075 => x"1f",
          5076 => x"34",
          5077 => x"17",
          5078 => x"82",
          5079 => x"83",
          5080 => x"84",
          5081 => x"66",
          5082 => x"fd",
          5083 => x"51",
          5084 => x"3f",
          5085 => x"17",
          5086 => x"c8",
          5087 => x"bf",
          5088 => x"86",
          5089 => x"d3",
          5090 => x"17",
          5091 => x"83",
          5092 => x"ff",
          5093 => x"65",
          5094 => x"1f",
          5095 => x"dc",
          5096 => x"77",
          5097 => x"79",
          5098 => x"ae",
          5099 => x"91",
          5100 => x"a3",
          5101 => x"80",
          5102 => x"ff",
          5103 => x"81",
          5104 => x"c8",
          5105 => x"8d",
          5106 => x"8b",
          5107 => x"87",
          5108 => x"83",
          5109 => x"76",
          5110 => x"0c",
          5111 => x"04",
          5112 => x"73",
          5113 => x"26",
          5114 => x"71",
          5115 => x"b1",
          5116 => x"71",
          5117 => x"c1",
          5118 => x"80",
          5119 => x"d4",
          5120 => x"84",
          5121 => x"9e",
          5122 => x"39",
          5123 => x"51",
          5124 => x"3f",
          5125 => x"91",
          5126 => x"ff",
          5127 => x"81",
          5128 => x"c2",
          5129 => x"ff",
          5130 => x"a8",
          5131 => x"cc",
          5132 => x"f2",
          5133 => x"39",
          5134 => x"51",
          5135 => x"3f",
          5136 => x"91",
          5137 => x"fe",
          5138 => x"81",
          5139 => x"c3",
          5140 => x"ff",
          5141 => x"fc",
          5142 => x"a0",
          5143 => x"c6",
          5144 => x"39",
          5145 => x"51",
          5146 => x"3f",
          5147 => x"91",
          5148 => x"fe",
          5149 => x"80",
          5150 => x"c3",
          5151 => x"ff",
          5152 => x"d0",
          5153 => x"94",
          5154 => x"9a",
          5155 => x"39",
          5156 => x"51",
          5157 => x"3f",
          5158 => x"c4",
          5159 => x"ff",
          5160 => x"39",
          5161 => x"51",
          5162 => x"3f",
          5163 => x"c4",
          5164 => x"fe",
          5165 => x"39",
          5166 => x"51",
          5167 => x"3f",
          5168 => x"c5",
          5169 => x"fe",
          5170 => x"39",
          5171 => x"51",
          5172 => x"3f",
          5173 => x"04",
          5174 => x"77",
          5175 => x"74",
          5176 => x"93",
          5177 => x"75",
          5178 => x"51",
          5179 => x"3f",
          5180 => x"08",
          5181 => x"87",
          5182 => x"51",
          5183 => x"3f",
          5184 => x"08",
          5185 => x"fe",
          5186 => x"91",
          5187 => x"55",
          5188 => x"53",
          5189 => x"c5",
          5190 => x"84",
          5191 => x"3d",
          5192 => x"ec",
          5193 => x"97",
          5194 => x"99",
          5195 => x"88",
          5196 => x"05",
          5197 => x"30",
          5198 => x"80",
          5199 => x"75",
          5200 => x"59",
          5201 => x"58",
          5202 => x"81",
          5203 => x"53",
          5204 => x"96",
          5205 => x"05",
          5206 => x"99",
          5207 => x"c8",
          5208 => x"d3",
          5209 => x"38",
          5210 => x"08",
          5211 => x"88",
          5212 => x"c8",
          5213 => x"96",
          5214 => x"11",
          5215 => x"80",
          5216 => x"fb",
          5217 => x"c0",
          5218 => x"d3",
          5219 => x"91",
          5220 => x"8e",
          5221 => x"2e",
          5222 => x"19",
          5223 => x"59",
          5224 => x"96",
          5225 => x"05",
          5226 => x"3f",
          5227 => x"79",
          5228 => x"7b",
          5229 => x"2a",
          5230 => x"57",
          5231 => x"80",
          5232 => x"91",
          5233 => x"87",
          5234 => x"08",
          5235 => x"fe",
          5236 => x"55",
          5237 => x"c8",
          5238 => x"3d",
          5239 => x"3d",
          5240 => x"05",
          5241 => x"7d",
          5242 => x"53",
          5243 => x"51",
          5244 => x"91",
          5245 => x"a4",
          5246 => x"2e",
          5247 => x"81",
          5248 => x"98",
          5249 => x"60",
          5250 => x"c8",
          5251 => x"7e",
          5252 => x"91",
          5253 => x"59",
          5254 => x"04",
          5255 => x"c8",
          5256 => x"0d",
          5257 => x"0d",
          5258 => x"33",
          5259 => x"53",
          5260 => x"52",
          5261 => x"e8",
          5262 => x"e8",
          5263 => x"55",
          5264 => x"3f",
          5265 => x"54",
          5266 => x"53",
          5267 => x"52",
          5268 => x"51",
          5269 => x"3f",
          5270 => x"85",
          5271 => x"ff",
          5272 => x"0d",
          5273 => x"0d",
          5274 => x"80",
          5275 => x"f9",
          5276 => x"51",
          5277 => x"3f",
          5278 => x"51",
          5279 => x"3f",
          5280 => x"ee",
          5281 => x"81",
          5282 => x"06",
          5283 => x"80",
          5284 => x"81",
          5285 => x"de",
          5286 => x"cc",
          5287 => x"d4",
          5288 => x"fe",
          5289 => x"72",
          5290 => x"81",
          5291 => x"71",
          5292 => x"38",
          5293 => x"ee",
          5294 => x"c6",
          5295 => x"f0",
          5296 => x"51",
          5297 => x"3f",
          5298 => x"70",
          5299 => x"52",
          5300 => x"95",
          5301 => x"fe",
          5302 => x"91",
          5303 => x"fe",
          5304 => x"80",
          5305 => x"8e",
          5306 => x"2a",
          5307 => x"51",
          5308 => x"2e",
          5309 => x"51",
          5310 => x"3f",
          5311 => x"51",
          5312 => x"3f",
          5313 => x"ed",
          5314 => x"85",
          5315 => x"06",
          5316 => x"80",
          5317 => x"81",
          5318 => x"da",
          5319 => x"98",
          5320 => x"d0",
          5321 => x"fe",
          5322 => x"72",
          5323 => x"81",
          5324 => x"71",
          5325 => x"38",
          5326 => x"ed",
          5327 => x"c7",
          5328 => x"ef",
          5329 => x"51",
          5330 => x"3f",
          5331 => x"70",
          5332 => x"52",
          5333 => x"95",
          5334 => x"fe",
          5335 => x"91",
          5336 => x"fe",
          5337 => x"80",
          5338 => x"8a",
          5339 => x"2a",
          5340 => x"51",
          5341 => x"2e",
          5342 => x"51",
          5343 => x"3f",
          5344 => x"51",
          5345 => x"3f",
          5346 => x"ec",
          5347 => x"f8",
          5348 => x"3d",
          5349 => x"3d",
          5350 => x"08",
          5351 => x"57",
          5352 => x"80",
          5353 => x"39",
          5354 => x"85",
          5355 => x"80",
          5356 => x"15",
          5357 => x"33",
          5358 => x"a0",
          5359 => x"81",
          5360 => x"70",
          5361 => x"06",
          5362 => x"e6",
          5363 => x"53",
          5364 => x"09",
          5365 => x"38",
          5366 => x"81",
          5367 => x"80",
          5368 => x"29",
          5369 => x"05",
          5370 => x"70",
          5371 => x"fe",
          5372 => x"91",
          5373 => x"8b",
          5374 => x"33",
          5375 => x"2e",
          5376 => x"81",
          5377 => x"ff",
          5378 => x"bb",
          5379 => x"38",
          5380 => x"91",
          5381 => x"88",
          5382 => x"ce",
          5383 => x"70",
          5384 => x"72",
          5385 => x"5e",
          5386 => x"81",
          5387 => x"ff",
          5388 => x"91",
          5389 => x"81",
          5390 => x"78",
          5391 => x"81",
          5392 => x"91",
          5393 => x"96",
          5394 => x"59",
          5395 => x"3f",
          5396 => x"52",
          5397 => x"51",
          5398 => x"3f",
          5399 => x"08",
          5400 => x"2e",
          5401 => x"c8",
          5402 => x"fd",
          5403 => x"39",
          5404 => x"5c",
          5405 => x"51",
          5406 => x"3f",
          5407 => x"43",
          5408 => x"70",
          5409 => x"52",
          5410 => x"e4",
          5411 => x"52",
          5412 => x"fd",
          5413 => x"3d",
          5414 => x"51",
          5415 => x"91",
          5416 => x"90",
          5417 => x"2c",
          5418 => x"81",
          5419 => x"af",
          5420 => x"10",
          5421 => x"05",
          5422 => x"04",
          5423 => x"f4",
          5424 => x"f8",
          5425 => x"fe",
          5426 => x"d3",
          5427 => x"38",
          5428 => x"51",
          5429 => x"3f",
          5430 => x"b4",
          5431 => x"11",
          5432 => x"05",
          5433 => x"c3",
          5434 => x"c8",
          5435 => x"88",
          5436 => x"25",
          5437 => x"40",
          5438 => x"33",
          5439 => x"c3",
          5440 => x"ff",
          5441 => x"91",
          5442 => x"81",
          5443 => x"78",
          5444 => x"c8",
          5445 => x"f6",
          5446 => x"5d",
          5447 => x"91",
          5448 => x"fe",
          5449 => x"fe",
          5450 => x"3d",
          5451 => x"53",
          5452 => x"51",
          5453 => x"3f",
          5454 => x"08",
          5455 => x"b4",
          5456 => x"80",
          5457 => x"c3",
          5458 => x"ff",
          5459 => x"91",
          5460 => x"52",
          5461 => x"51",
          5462 => x"3f",
          5463 => x"b4",
          5464 => x"11",
          5465 => x"05",
          5466 => x"bf",
          5467 => x"c8",
          5468 => x"87",
          5469 => x"26",
          5470 => x"b4",
          5471 => x"11",
          5472 => x"05",
          5473 => x"a3",
          5474 => x"c8",
          5475 => x"91",
          5476 => x"40",
          5477 => x"c9",
          5478 => x"3d",
          5479 => x"fe",
          5480 => x"02",
          5481 => x"53",
          5482 => x"84",
          5483 => x"e0",
          5484 => x"ff",
          5485 => x"91",
          5486 => x"80",
          5487 => x"91",
          5488 => x"51",
          5489 => x"fd",
          5490 => x"c8",
          5491 => x"f4",
          5492 => x"5c",
          5493 => x"b4",
          5494 => x"05",
          5495 => x"a4",
          5496 => x"c8",
          5497 => x"fe",
          5498 => x"5b",
          5499 => x"3f",
          5500 => x"d3",
          5501 => x"7a",
          5502 => x"3f",
          5503 => x"08",
          5504 => x"f0",
          5505 => x"c8",
          5506 => x"d4",
          5507 => x"39",
          5508 => x"f8",
          5509 => x"e3",
          5510 => x"d3",
          5511 => x"3d",
          5512 => x"52",
          5513 => x"c1",
          5514 => x"c8",
          5515 => x"fe",
          5516 => x"5a",
          5517 => x"3f",
          5518 => x"08",
          5519 => x"f8",
          5520 => x"fe",
          5521 => x"91",
          5522 => x"91",
          5523 => x"80",
          5524 => x"91",
          5525 => x"81",
          5526 => x"78",
          5527 => x"7a",
          5528 => x"3f",
          5529 => x"08",
          5530 => x"88",
          5531 => x"c8",
          5532 => x"ec",
          5533 => x"39",
          5534 => x"51",
          5535 => x"3f",
          5536 => x"f2",
          5537 => x"ec",
          5538 => x"b0",
          5539 => x"96",
          5540 => x"fe",
          5541 => x"fb",
          5542 => x"80",
          5543 => x"c0",
          5544 => x"84",
          5545 => x"87",
          5546 => x"0c",
          5547 => x"51",
          5548 => x"3f",
          5549 => x"91",
          5550 => x"fe",
          5551 => x"8c",
          5552 => x"87",
          5553 => x"0c",
          5554 => x"0b",
          5555 => x"94",
          5556 => x"39",
          5557 => x"f4",
          5558 => x"f8",
          5559 => x"fa",
          5560 => x"d3",
          5561 => x"2e",
          5562 => x"60",
          5563 => x"f0",
          5564 => x"ac",
          5565 => x"78",
          5566 => x"fe",
          5567 => x"fe",
          5568 => x"fe",
          5569 => x"91",
          5570 => x"80",
          5571 => x"38",
          5572 => x"ca",
          5573 => x"f8",
          5574 => x"59",
          5575 => x"d3",
          5576 => x"91",
          5577 => x"80",
          5578 => x"38",
          5579 => x"08",
          5580 => x"a8",
          5581 => x"e8",
          5582 => x"39",
          5583 => x"51",
          5584 => x"3f",
          5585 => x"3f",
          5586 => x"91",
          5587 => x"fe",
          5588 => x"80",
          5589 => x"39",
          5590 => x"3f",
          5591 => x"61",
          5592 => x"59",
          5593 => x"fa",
          5594 => x"7c",
          5595 => x"80",
          5596 => x"38",
          5597 => x"f8",
          5598 => x"e1",
          5599 => x"ca",
          5600 => x"d3",
          5601 => x"91",
          5602 => x"80",
          5603 => x"fc",
          5604 => x"70",
          5605 => x"f7",
          5606 => x"cb",
          5607 => x"d3",
          5608 => x"56",
          5609 => x"42",
          5610 => x"54",
          5611 => x"53",
          5612 => x"52",
          5613 => x"a6",
          5614 => x"c8",
          5615 => x"81",
          5616 => x"32",
          5617 => x"8a",
          5618 => x"2e",
          5619 => x"f9",
          5620 => x"cb",
          5621 => x"f6",
          5622 => x"98",
          5623 => x"0d",
          5624 => x"d3",
          5625 => x"90",
          5626 => x"87",
          5627 => x"0c",
          5628 => x"e4",
          5629 => x"94",
          5630 => x"80",
          5631 => x"c0",
          5632 => x"8c",
          5633 => x"87",
          5634 => x"0c",
          5635 => x"0b",
          5636 => x"0c",
          5637 => x"0b",
          5638 => x"0c",
          5639 => x"3f",
          5640 => x"3f",
          5641 => x"51",
          5642 => x"3f",
          5643 => x"51",
          5644 => x"3f",
          5645 => x"51",
          5646 => x"3f",
          5647 => x"e5",
          5648 => x"3f",
          5649 => x"00",
          5650 => x"00",
          5651 => x"00",
          5652 => x"00",
          5653 => x"00",
          5654 => x"00",
          5655 => x"00",
          5656 => x"00",
          5657 => x"00",
          5658 => x"00",
          5659 => x"00",
          5660 => x"00",
          5661 => x"00",
          5662 => x"00",
          5663 => x"00",
          5664 => x"00",
          5665 => x"00",
          5666 => x"00",
          5667 => x"00",
          5668 => x"00",
          5669 => x"00",
          5670 => x"00",
          5671 => x"00",
          5672 => x"00",
          5673 => x"00",
          5674 => x"00",
          5675 => x"00",
          5676 => x"00",
          5677 => x"00",
          5678 => x"00",
          5679 => x"00",
          5680 => x"00",
          5681 => x"00",
          5682 => x"00",
          5683 => x"00",
          5684 => x"00",
          5685 => x"00",
          5686 => x"00",
          5687 => x"00",
          5688 => x"00",
          5689 => x"00",
          5690 => x"00",
          5691 => x"00",
          5692 => x"00",
          5693 => x"00",
          5694 => x"00",
          5695 => x"00",
          5696 => x"00",
          5697 => x"00",
          5698 => x"00",
          5699 => x"00",
          5700 => x"00",
          5701 => x"00",
          5702 => x"00",
          5703 => x"00",
          5704 => x"00",
          5705 => x"00",
          5706 => x"00",
          5707 => x"00",
          5708 => x"00",
          5709 => x"00",
          5710 => x"00",
          5711 => x"00",
          5712 => x"00",
          5713 => x"00",
          5714 => x"00",
          5715 => x"00",
          5716 => x"00",
          5717 => x"00",
          5718 => x"00",
          5719 => x"00",
          5720 => x"00",
          5721 => x"00",
          5722 => x"00",
          5723 => x"00",
          5724 => x"00",
          5725 => x"00",
          5726 => x"00",
          5727 => x"00",
          5728 => x"00",
          5729 => x"00",
          5730 => x"00",
          5731 => x"00",
          5732 => x"00",
          5733 => x"00",
          5734 => x"00",
          5735 => x"00",
          5736 => x"00",
          5737 => x"00",
          5738 => x"00",
          5739 => x"00",
          5740 => x"00",
          5741 => x"00",
          5742 => x"00",
          5743 => x"00",
          5744 => x"00",
          5745 => x"00",
          5746 => x"00",
          5747 => x"00",
          5748 => x"00",
          5749 => x"00",
          5750 => x"00",
          5751 => x"00",
          5752 => x"00",
          5753 => x"00",
          5754 => x"00",
          5755 => x"00",
          5756 => x"00",
          5757 => x"00",
          5758 => x"00",
          5759 => x"00",
          5760 => x"00",
          5761 => x"00",
          5762 => x"00",
          5763 => x"00",
          5764 => x"00",
          5765 => x"00",
          5766 => x"00",
          5767 => x"00",
          5768 => x"00",
          5769 => x"00",
          5770 => x"00",
          5771 => x"00",
          5772 => x"00",
          5773 => x"00",
          5774 => x"00",
          5775 => x"00",
          5776 => x"00",
          5777 => x"00",
          5778 => x"00",
          5779 => x"00",
          5780 => x"00",
          5781 => x"00",
          5782 => x"00",
          5783 => x"00",
          5784 => x"00",
          5785 => x"00",
          5786 => x"00",
          5787 => x"00",
          5788 => x"00",
          5789 => x"00",
          5790 => x"00",
          5791 => x"00",
          5792 => x"00",
          5793 => x"00",
          5794 => x"00",
          5795 => x"00",
          5796 => x"00",
          5797 => x"00",
          5798 => x"00",
          5799 => x"00",
          5800 => x"00",
          5801 => x"00",
          5802 => x"00",
          5803 => x"00",
          5804 => x"00",
          5805 => x"00",
          5806 => x"00",
          5807 => x"00",
          5808 => x"00",
          5809 => x"00",
          5810 => x"00",
          5811 => x"00",
          5812 => x"00",
          5813 => x"00",
          5814 => x"00",
          5815 => x"00",
          5816 => x"00",
          5817 => x"00",
          5818 => x"00",
          5819 => x"00",
          5820 => x"00",
          5821 => x"00",
          5822 => x"00",
          5823 => x"00",
          5824 => x"00",
          5825 => x"00",
          5826 => x"00",
          5827 => x"00",
          5828 => x"00",
          5829 => x"00",
          5830 => x"00",
          5831 => x"00",
          5832 => x"00",
          5833 => x"00",
          5834 => x"25",
          5835 => x"64",
          5836 => x"20",
          5837 => x"25",
          5838 => x"64",
          5839 => x"25",
          5840 => x"53",
          5841 => x"43",
          5842 => x"69",
          5843 => x"61",
          5844 => x"6e",
          5845 => x"20",
          5846 => x"6f",
          5847 => x"6f",
          5848 => x"6f",
          5849 => x"67",
          5850 => x"3a",
          5851 => x"76",
          5852 => x"73",
          5853 => x"70",
          5854 => x"65",
          5855 => x"64",
          5856 => x"20",
          5857 => x"49",
          5858 => x"20",
          5859 => x"4d",
          5860 => x"74",
          5861 => x"3d",
          5862 => x"58",
          5863 => x"69",
          5864 => x"25",
          5865 => x"29",
          5866 => x"20",
          5867 => x"42",
          5868 => x"20",
          5869 => x"61",
          5870 => x"25",
          5871 => x"2c",
          5872 => x"7a",
          5873 => x"30",
          5874 => x"2e",
          5875 => x"20",
          5876 => x"52",
          5877 => x"28",
          5878 => x"72",
          5879 => x"30",
          5880 => x"20",
          5881 => x"65",
          5882 => x"38",
          5883 => x"0a",
          5884 => x"20",
          5885 => x"49",
          5886 => x"4c",
          5887 => x"20",
          5888 => x"50",
          5889 => x"00",
          5890 => x"20",
          5891 => x"53",
          5892 => x"00",
          5893 => x"20",
          5894 => x"53",
          5895 => x"61",
          5896 => x"28",
          5897 => x"69",
          5898 => x"3d",
          5899 => x"58",
          5900 => x"00",
          5901 => x"20",
          5902 => x"49",
          5903 => x"52",
          5904 => x"54",
          5905 => x"4e",
          5906 => x"4c",
          5907 => x"0a",
          5908 => x"20",
          5909 => x"54",
          5910 => x"52",
          5911 => x"54",
          5912 => x"72",
          5913 => x"30",
          5914 => x"2e",
          5915 => x"41",
          5916 => x"65",
          5917 => x"73",
          5918 => x"20",
          5919 => x"43",
          5920 => x"52",
          5921 => x"74",
          5922 => x"63",
          5923 => x"20",
          5924 => x"72",
          5925 => x"20",
          5926 => x"30",
          5927 => x"00",
          5928 => x"20",
          5929 => x"43",
          5930 => x"4d",
          5931 => x"72",
          5932 => x"74",
          5933 => x"20",
          5934 => x"72",
          5935 => x"20",
          5936 => x"30",
          5937 => x"00",
          5938 => x"20",
          5939 => x"53",
          5940 => x"6b",
          5941 => x"61",
          5942 => x"41",
          5943 => x"65",
          5944 => x"20",
          5945 => x"20",
          5946 => x"30",
          5947 => x"00",
          5948 => x"20",
          5949 => x"5a",
          5950 => x"49",
          5951 => x"20",
          5952 => x"20",
          5953 => x"20",
          5954 => x"20",
          5955 => x"20",
          5956 => x"30",
          5957 => x"00",
          5958 => x"20",
          5959 => x"53",
          5960 => x"65",
          5961 => x"6c",
          5962 => x"20",
          5963 => x"71",
          5964 => x"20",
          5965 => x"20",
          5966 => x"30",
          5967 => x"00",
          5968 => x"53",
          5969 => x"6c",
          5970 => x"4d",
          5971 => x"75",
          5972 => x"46",
          5973 => x"00",
          5974 => x"45",
          5975 => x"45",
          5976 => x"69",
          5977 => x"55",
          5978 => x"6f",
          5979 => x"53",
          5980 => x"22",
          5981 => x"3a",
          5982 => x"3e",
          5983 => x"7c",
          5984 => x"46",
          5985 => x"46",
          5986 => x"32",
          5987 => x"30",
          5988 => x"31",
          5989 => x"32",
          5990 => x"33",
          5991 => x"35",
          5992 => x"36",
          5993 => x"37",
          5994 => x"38",
          5995 => x"39",
          5996 => x"31",
          5997 => x"eb",
          5998 => x"53",
          5999 => x"35",
          6000 => x"4e",
          6001 => x"41",
          6002 => x"20",
          6003 => x"41",
          6004 => x"20",
          6005 => x"4e",
          6006 => x"41",
          6007 => x"20",
          6008 => x"41",
          6009 => x"20",
          6010 => x"00",
          6011 => x"00",
          6012 => x"00",
          6013 => x"00",
          6014 => x"80",
          6015 => x"8e",
          6016 => x"45",
          6017 => x"49",
          6018 => x"90",
          6019 => x"99",
          6020 => x"59",
          6021 => x"9c",
          6022 => x"41",
          6023 => x"a5",
          6024 => x"a8",
          6025 => x"ac",
          6026 => x"b0",
          6027 => x"b4",
          6028 => x"b8",
          6029 => x"bc",
          6030 => x"c0",
          6031 => x"c4",
          6032 => x"c8",
          6033 => x"cc",
          6034 => x"d0",
          6035 => x"d4",
          6036 => x"d8",
          6037 => x"dc",
          6038 => x"e0",
          6039 => x"e4",
          6040 => x"e8",
          6041 => x"ec",
          6042 => x"f0",
          6043 => x"f4",
          6044 => x"f8",
          6045 => x"fc",
          6046 => x"2b",
          6047 => x"3d",
          6048 => x"5c",
          6049 => x"3c",
          6050 => x"7f",
          6051 => x"00",
          6052 => x"00",
          6053 => x"01",
          6054 => x"00",
          6055 => x"00",
          6056 => x"00",
          6057 => x"00",
          6058 => x"00",
          6059 => x"46",
          6060 => x"32",
          6061 => x"46",
          6062 => x"36",
          6063 => x"65",
          6064 => x"54",
          6065 => x"44",
          6066 => x"20",
          6067 => x"43",
          6068 => x"52",
          6069 => x"00",
          6070 => x"44",
          6071 => x"20",
          6072 => x"46",
          6073 => x"43",
          6074 => x"52",
          6075 => x"00",
          6076 => x"46",
          6077 => x"53",
          6078 => x"45",
          6079 => x"4f",
          6080 => x"4f",
          6081 => x"4d",
          6082 => x"52",
          6083 => x"48",
          6084 => x"57",
          6085 => x"00",
          6086 => x"54",
          6087 => x"49",
          6088 => x"45",
          6089 => x"55",
          6090 => x"4e",
          6091 => x"4d",
          6092 => x"20",
          6093 => x"4d",
          6094 => x"53",
          6095 => x"64",
          6096 => x"70",
          6097 => x"64",
          6098 => x"74",
          6099 => x"64",
          6100 => x"74",
          6101 => x"64",
          6102 => x"74",
          6103 => x"62",
          6104 => x"70",
          6105 => x"62",
          6106 => x"74",
          6107 => x"62",
          6108 => x"64",
          6109 => x"62",
          6110 => x"74",
          6111 => x"62",
          6112 => x"6c",
          6113 => x"62",
          6114 => x"00",
          6115 => x"66",
          6116 => x"74",
          6117 => x"66",
          6118 => x"6e",
          6119 => x"66",
          6120 => x"73",
          6121 => x"66",
          6122 => x"6b",
          6123 => x"66",
          6124 => x"64",
          6125 => x"66",
          6126 => x"70",
          6127 => x"00",
          6128 => x"66",
          6129 => x"74",
          6130 => x"66",
          6131 => x"6e",
          6132 => x"66",
          6133 => x"6f",
          6134 => x"66",
          6135 => x"72",
          6136 => x"66",
          6137 => x"65",
          6138 => x"66",
          6139 => x"61",
          6140 => x"66",
          6141 => x"00",
          6142 => x"66",
          6143 => x"69",
          6144 => x"66",
          6145 => x"74",
          6146 => x"66",
          6147 => x"00",
          6148 => x"66",
          6149 => x"00",
          6150 => x"66",
          6151 => x"66",
          6152 => x"63",
          6153 => x"66",
          6154 => x"61",
          6155 => x"66",
          6156 => x"64",
          6157 => x"66",
          6158 => x"63",
          6159 => x"66",
          6160 => x"65",
          6161 => x"66",
          6162 => x"70",
          6163 => x"66",
          6164 => x"66",
          6165 => x"76",
          6166 => x"66",
          6167 => x"77",
          6168 => x"00",
          6169 => x"66",
          6170 => x"65",
          6171 => x"66",
          6172 => x"73",
          6173 => x"6d",
          6174 => x"00",
          6175 => x"6d",
          6176 => x"70",
          6177 => x"6d",
          6178 => x"6d",
          6179 => x"6d",
          6180 => x"68",
          6181 => x"68",
          6182 => x"68",
          6183 => x"68",
          6184 => x"68",
          6185 => x"68",
          6186 => x"64",
          6187 => x"00",
          6188 => x"63",
          6189 => x"6d",
          6190 => x"00",
          6191 => x"63",
          6192 => x"00",
          6193 => x"6a",
          6194 => x"72",
          6195 => x"61",
          6196 => x"72",
          6197 => x"74",
          6198 => x"68",
          6199 => x"00",
          6200 => x"69",
          6201 => x"00",
          6202 => x"74",
          6203 => x"00",
          6204 => x"74",
          6205 => x"00",
          6206 => x"44",
          6207 => x"20",
          6208 => x"6f",
          6209 => x"49",
          6210 => x"72",
          6211 => x"20",
          6212 => x"6f",
          6213 => x"00",
          6214 => x"44",
          6215 => x"20",
          6216 => x"20",
          6217 => x"64",
          6218 => x"00",
          6219 => x"4e",
          6220 => x"69",
          6221 => x"66",
          6222 => x"64",
          6223 => x"4e",
          6224 => x"61",
          6225 => x"66",
          6226 => x"64",
          6227 => x"49",
          6228 => x"6c",
          6229 => x"66",
          6230 => x"6e",
          6231 => x"2e",
          6232 => x"41",
          6233 => x"73",
          6234 => x"65",
          6235 => x"64",
          6236 => x"46",
          6237 => x"20",
          6238 => x"65",
          6239 => x"20",
          6240 => x"73",
          6241 => x"0a",
          6242 => x"46",
          6243 => x"20",
          6244 => x"64",
          6245 => x"69",
          6246 => x"6c",
          6247 => x"0a",
          6248 => x"53",
          6249 => x"73",
          6250 => x"69",
          6251 => x"70",
          6252 => x"65",
          6253 => x"64",
          6254 => x"44",
          6255 => x"65",
          6256 => x"6d",
          6257 => x"20",
          6258 => x"69",
          6259 => x"6c",
          6260 => x"0a",
          6261 => x"44",
          6262 => x"20",
          6263 => x"20",
          6264 => x"62",
          6265 => x"2e",
          6266 => x"4e",
          6267 => x"6f",
          6268 => x"74",
          6269 => x"65",
          6270 => x"6c",
          6271 => x"73",
          6272 => x"20",
          6273 => x"6e",
          6274 => x"6e",
          6275 => x"73",
          6276 => x"00",
          6277 => x"46",
          6278 => x"61",
          6279 => x"62",
          6280 => x"65",
          6281 => x"00",
          6282 => x"54",
          6283 => x"6f",
          6284 => x"20",
          6285 => x"72",
          6286 => x"6f",
          6287 => x"61",
          6288 => x"6c",
          6289 => x"2e",
          6290 => x"46",
          6291 => x"20",
          6292 => x"6c",
          6293 => x"65",
          6294 => x"00",
          6295 => x"49",
          6296 => x"66",
          6297 => x"69",
          6298 => x"20",
          6299 => x"6f",
          6300 => x"0a",
          6301 => x"54",
          6302 => x"6d",
          6303 => x"20",
          6304 => x"6e",
          6305 => x"6c",
          6306 => x"0a",
          6307 => x"50",
          6308 => x"6d",
          6309 => x"72",
          6310 => x"6e",
          6311 => x"72",
          6312 => x"2e",
          6313 => x"53",
          6314 => x"65",
          6315 => x"0a",
          6316 => x"55",
          6317 => x"6f",
          6318 => x"65",
          6319 => x"72",
          6320 => x"0a",
          6321 => x"20",
          6322 => x"65",
          6323 => x"73",
          6324 => x"20",
          6325 => x"20",
          6326 => x"65",
          6327 => x"65",
          6328 => x"00",
          6329 => x"72",
          6330 => x"00",
          6331 => x"5a",
          6332 => x"41",
          6333 => x"0a",
          6334 => x"25",
          6335 => x"00",
          6336 => x"31",
          6337 => x"37",
          6338 => x"31",
          6339 => x"76",
          6340 => x"00",
          6341 => x"20",
          6342 => x"2c",
          6343 => x"76",
          6344 => x"32",
          6345 => x"25",
          6346 => x"73",
          6347 => x"0a",
          6348 => x"5a",
          6349 => x"41",
          6350 => x"74",
          6351 => x"75",
          6352 => x"48",
          6353 => x"6c",
          6354 => x"00",
          6355 => x"54",
          6356 => x"72",
          6357 => x"74",
          6358 => x"75",
          6359 => x"00",
          6360 => x"50",
          6361 => x"69",
          6362 => x"72",
          6363 => x"74",
          6364 => x"49",
          6365 => x"4c",
          6366 => x"20",
          6367 => x"65",
          6368 => x"70",
          6369 => x"49",
          6370 => x"4c",
          6371 => x"20",
          6372 => x"65",
          6373 => x"70",
          6374 => x"55",
          6375 => x"30",
          6376 => x"20",
          6377 => x"65",
          6378 => x"70",
          6379 => x"55",
          6380 => x"30",
          6381 => x"20",
          6382 => x"65",
          6383 => x"70",
          6384 => x"55",
          6385 => x"31",
          6386 => x"20",
          6387 => x"65",
          6388 => x"70",
          6389 => x"55",
          6390 => x"31",
          6391 => x"20",
          6392 => x"65",
          6393 => x"70",
          6394 => x"53",
          6395 => x"69",
          6396 => x"75",
          6397 => x"69",
          6398 => x"2e",
          6399 => x"00",
          6400 => x"45",
          6401 => x"6c",
          6402 => x"20",
          6403 => x"65",
          6404 => x"2e",
          6405 => x"30",
          6406 => x"46",
          6407 => x"65",
          6408 => x"6f",
          6409 => x"69",
          6410 => x"6c",
          6411 => x"20",
          6412 => x"63",
          6413 => x"20",
          6414 => x"70",
          6415 => x"73",
          6416 => x"6e",
          6417 => x"6d",
          6418 => x"61",
          6419 => x"2e",
          6420 => x"2a",
          6421 => x"42",
          6422 => x"64",
          6423 => x"20",
          6424 => x"0a",
          6425 => x"49",
          6426 => x"69",
          6427 => x"73",
          6428 => x"0a",
          6429 => x"46",
          6430 => x"65",
          6431 => x"6f",
          6432 => x"69",
          6433 => x"6c",
          6434 => x"2e",
          6435 => x"72",
          6436 => x"64",
          6437 => x"25",
          6438 => x"44",
          6439 => x"62",
          6440 => x"67",
          6441 => x"74",
          6442 => x"75",
          6443 => x"0a",
          6444 => x"45",
          6445 => x"6c",
          6446 => x"20",
          6447 => x"65",
          6448 => x"70",
          6449 => x"00",
          6450 => x"44",
          6451 => x"62",
          6452 => x"20",
          6453 => x"74",
          6454 => x"66",
          6455 => x"45",
          6456 => x"6c",
          6457 => x"20",
          6458 => x"74",
          6459 => x"66",
          6460 => x"45",
          6461 => x"75",
          6462 => x"67",
          6463 => x"64",
          6464 => x"20",
          6465 => x"78",
          6466 => x"2e",
          6467 => x"43",
          6468 => x"69",
          6469 => x"63",
          6470 => x"20",
          6471 => x"30",
          6472 => x"2e",
          6473 => x"00",
          6474 => x"43",
          6475 => x"20",
          6476 => x"75",
          6477 => x"64",
          6478 => x"64",
          6479 => x"25",
          6480 => x"0a",
          6481 => x"52",
          6482 => x"61",
          6483 => x"6e",
          6484 => x"70",
          6485 => x"63",
          6486 => x"6f",
          6487 => x"2e",
          6488 => x"43",
          6489 => x"20",
          6490 => x"6f",
          6491 => x"6e",
          6492 => x"2e",
          6493 => x"5a",
          6494 => x"62",
          6495 => x"25",
          6496 => x"25",
          6497 => x"73",
          6498 => x"00",
          6499 => x"42",
          6500 => x"63",
          6501 => x"61",
          6502 => x"0a",
          6503 => x"52",
          6504 => x"69",
          6505 => x"2e",
          6506 => x"45",
          6507 => x"6c",
          6508 => x"20",
          6509 => x"65",
          6510 => x"70",
          6511 => x"2e",
          6512 => x"00",
          6513 => x"00",
          6514 => x"00",
          6515 => x"00",
          6516 => x"00",
          6517 => x"00",
          6518 => x"00",
          6519 => x"00",
          6520 => x"00",
          6521 => x"00",
          6522 => x"00",
          6523 => x"05",
          6524 => x"00",
          6525 => x"01",
          6526 => x"80",
          6527 => x"01",
          6528 => x"00",
          6529 => x"01",
          6530 => x"00",
          6531 => x"00",
          6532 => x"00",
          6533 => x"00",
          6534 => x"00",
          6535 => x"01",
          6536 => x"00",
          6537 => x"00",
          6538 => x"00",
          6539 => x"00",
          6540 => x"00",
          6541 => x"00",
          6542 => x"00",
          6543 => x"01",
          6544 => x"00",
          6545 => x"00",
          6546 => x"00",
          6547 => x"00",
          6548 => x"00",
          6549 => x"00",
          6550 => x"00",
          6551 => x"00",
          6552 => x"00",
          6553 => x"00",
          6554 => x"00",
          6555 => x"00",
          6556 => x"00",
          6557 => x"00",
          6558 => x"00",
          6559 => x"00",
          6560 => x"00",
          6561 => x"00",
          6562 => x"00",
          6563 => x"00",
          6564 => x"00",
          6565 => x"00",
          6566 => x"00",
          6567 => x"00",
          6568 => x"00",
          6569 => x"00",
          6570 => x"00",
          6571 => x"01",
          6572 => x"00",
          6573 => x"00",
          6574 => x"00",
          6575 => x"00",
          6576 => x"00",
          6577 => x"00",
          6578 => x"00",
          6579 => x"00",
          6580 => x"00",
          6581 => x"00",
          6582 => x"00",
          6583 => x"00",
          6584 => x"00",
          6585 => x"00",
          6586 => x"00",
          6587 => x"00",
          6588 => x"00",
          6589 => x"00",
          6590 => x"00",
          6591 => x"00",
          6592 => x"00",
          6593 => x"00",
          6594 => x"00",
          6595 => x"00",
          6596 => x"00",
          6597 => x"00",
          6598 => x"00",
          6599 => x"00",
          6600 => x"00",
          6601 => x"00",
          6602 => x"00",
          6603 => x"00",
          6604 => x"00",
          6605 => x"00",
          6606 => x"00",
          6607 => x"00",
          6608 => x"00",
          6609 => x"00",
          6610 => x"00",
          6611 => x"00",
          6612 => x"00",
          6613 => x"00",
          6614 => x"00",
          6615 => x"00",
          6616 => x"00",
          6617 => x"00",
          6618 => x"00",
          6619 => x"00",
          6620 => x"00",
          6621 => x"00",
          6622 => x"00",
          6623 => x"00",
          6624 => x"00",
          6625 => x"00",
          6626 => x"00",
          6627 => x"00",
          6628 => x"00",
          6629 => x"00",
          6630 => x"00",
          6631 => x"00",
          6632 => x"00",
          6633 => x"00",
          6634 => x"00",
          6635 => x"00",
          6636 => x"00",
          6637 => x"00",
          6638 => x"00",
          6639 => x"00",
          6640 => x"00",
          6641 => x"00",
          6642 => x"00",
          6643 => x"00",
          6644 => x"00",
          6645 => x"00",
          6646 => x"00",
          6647 => x"00",
          6648 => x"00",
          6649 => x"00",
          6650 => x"00",
          6651 => x"01",
          6652 => x"00",
          6653 => x"00",
          6654 => x"00",
          6655 => x"01",
          6656 => x"00",
          6657 => x"00",
          6658 => x"00",
          6659 => x"00",
          6660 => x"00",
          6661 => x"00",
          6662 => x"00",
          6663 => x"00",
          6664 => x"00",
          6665 => x"00",
          6666 => x"00",
          6667 => x"00",
          6668 => x"00",
          6669 => x"00",
          6670 => x"00",
          6671 => x"00",
          6672 => x"00",
          6673 => x"00",
          6674 => x"00",
          6675 => x"00",
          6676 => x"00",
          6677 => x"00",
          6678 => x"00",
          6679 => x"00",
          6680 => x"00",
          6681 => x"00",
          6682 => x"00",
          6683 => x"00",
          6684 => x"00",
          6685 => x"00",
          6686 => x"00",
          6687 => x"00",
          6688 => x"00",
          6689 => x"00",
          6690 => x"00",
          6691 => x"00",
          6692 => x"00",
          6693 => x"00",
          6694 => x"00",
          6695 => x"00",
          6696 => x"00",
          6697 => x"00",
          6698 => x"00",
          6699 => x"00",
          6700 => x"00",
          6701 => x"00",
          6702 => x"00",
          6703 => x"00",
          6704 => x"00",
          6705 => x"00",
          6706 => x"00",
          6707 => x"01",
          6708 => x"00",
          6709 => x"00",
          6710 => x"00",
          6711 => x"01",
          6712 => x"00",
          6713 => x"00",
          6714 => x"00",
          6715 => x"00",
          6716 => x"00",
          6717 => x"00",
          6718 => x"00",
          6719 => x"00",
          6720 => x"00",
          6721 => x"00",
          6722 => x"00",
          6723 => x"01",
          6724 => x"00",
          6725 => x"00",
          6726 => x"00",
          6727 => x"01",
          6728 => x"00",
          6729 => x"00",
          6730 => x"00",
          6731 => x"00",
          6732 => x"00",
          6733 => x"00",
          6734 => x"00",
          6735 => x"00",
          6736 => x"00",
          6737 => x"00",
          6738 => x"00",
          6739 => x"01",
          6740 => x"00",
          6741 => x"00",
          6742 => x"00",
          6743 => x"01",
          6744 => x"00",
          6745 => x"00",
          6746 => x"00",
          6747 => x"01",
          6748 => x"00",
          6749 => x"00",
          6750 => x"00",
          6751 => x"01",
          6752 => x"00",
          6753 => x"00",
          6754 => x"00",
          6755 => x"00",
          6756 => x"00",
          6757 => x"00",
          6758 => x"00",
          6759 => x"01",
          6760 => x"00",
          6761 => x"00",
          6762 => x"00",
          6763 => x"00",
          6764 => x"00",
          6765 => x"00",
          6766 => x"00",
          6767 => x"01",
          6768 => x"00",
          6769 => x"00",
        others => X"00"
    );

    signal RAM0_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM1_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM2_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM3_DATA                       : std_logic_vector(7 downto 0);   -- Buffer for byte in word to be written.
    signal RAM0_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM1_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM2_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.
    signal RAM3_WREN                       : std_logic;                      -- Write Enable for this particular byte in word.

begin

    RAM0_DATA <= memAWrite(7 downto 0);
    RAM0_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "00") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM1_DATA <= memAWrite(15 downto 8)  when (memAWriteByte = '0' and memAWriteHalfWord = '0') or memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM1_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "01") or (memAWriteHalfWord = '1' and memAAddr(1) = '0'))
                 else '0';
    RAM2_DATA <= memAWrite(23 downto 16) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(7 downto 0);
    RAM2_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "10") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';
    RAM3_DATA <= memAWrite(31 downto 24) when (memAWriteByte = '0' and memAWriteHalfWord = '0')
                 else
                 memAWrite(15 downto 8)  when memAWriteHalfWord = '1'
                 else
                 memAWrite(7 downto 0);
    RAM3_WREN <= '1' when memAWriteEnable = '1' and ((memAWriteByte = '0' and memAWriteHalfWord = '0') or (memAWriteByte = '1' and memAAddr(1 downto 0) = "11") or (memAWriteHalfWord = '1' and memAAddr(1) = '1'))
                 else '0';

    -- RAM Byte 0 - Port A - bits 7 to 0
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM0_WREN = '1' then
                RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM0_DATA;
            else
                memARead(7 downto 0) <= RAM0(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 1 - Port A - bits 15 to 8
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM1_WREN = '1' then
                RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM1_DATA;
            else
                memARead(15 downto 8) <= RAM1(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 2 - Port A - bits 23 to 16 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM2_WREN = '1' then
                RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM2_DATA;
            else
                memARead(23 downto 16) <= RAM2(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;

    -- RAM Byte 3 - Port A - bits 31 to 24 
    process(clk)
    begin
        if rising_edge(clk) then
            if RAM3_WREN = '1' then
                RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2)))) := RAM3_DATA;
            else
                memARead(31 downto 24) <= RAM3(to_integer(unsigned(memAAddr(addrbits-1 downto 2))));
            end if;
        end if;
    end process;
end arch;
